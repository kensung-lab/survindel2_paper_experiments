SRR1766442.42445526 chr6 40209513 N chr6 40209764 N DUP 22
SRR1766469.1573710 chr6 40209513 N chr6 40209764 N DUP 22
SRR1766469.2711675 chr6 40209267 N chr6 40209776 N DEL 21
SRR1766444.5330388 chr6 40209267 N chr6 40209812 N DEL 23
SRR1766472.1493340 chr6 40209267 N chr6 40209812 N DEL 23
SRR1766450.2073233 chr6 40209343 N chr6 40209416 N DEL 23
SRR1766475.10669225 chr6 40209327 N chr6 40209528 N DEL 28
SRR1766449.5984102 chr6 40209267 N chr6 40209704 N DEL 22
SRR1766464.7652180 chr6 40209267 N chr6 40209704 N DEL 22
SRR1766442.26017208 chr6 40209267 N chr6 40209740 N DEL 24
SRR1766472.4368075 chr6 40209267 N chr6 40209740 N DEL 24
SRR1766459.619374 chr6 40209389 N chr6 40209812 N DEL 21
SRR1766466.2830877 chr6 40209389 N chr6 40209812 N DEL 21
SRR1766473.7390458 chr6 40209309 N chr6 40209422 N DEL 20
SRR1766462.2079898 chr6 40209327 N chr6 40209792 N DEL 29
SRR1766455.914097 chr6 40209327 N chr6 40209792 N DEL 28
SRR1766478.7660085 chr6 40209309 N chr6 40209422 N DEL 20
SRR1766472.8450164 chr6 40209322 N chr6 40209805 N DEL 23
SRR1766460.7211391 chr6 40209322 N chr6 40209805 N DEL 24
SRR1766451.1403969 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766481.6328673 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766477.7553933 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766442.33120376 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766450.3168715 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766445.9878414 chr6 40209470 N chr6 40209805 N DEL 25
SRR1766457.3977199 chr6 40209292 N chr6 40209805 N DEL 36
SRR1766462.2718922 chr6 40209297 N chr6 40209792 N DEL 31
SRR1766469.6318633 chr6 40209535 N chr6 40209850 N DUP 21
SRR1766462.670452 chr6 40209327 N chr6 40209528 N DEL 24
SRR1766446.6025057 chr6 40209597 N chr6 40209828 N DEL 23
SRR1766447.8376972 chr6 40209597 N chr6 40209828 N DEL 21
SRR1766485.5998535 chr6 40209605 N chr6 40209864 N DEL 31
SRR1766482.12819399 chr6 40209605 N chr6 40209864 N DEL 28
SRR1766468.5053632 chr6 40209605 N chr6 40209864 N DEL 22
SRR1766457.8845115 chr6 40209789 N chr6 40209910 N DUP 28
SRR1766471.5915735 chr6 40209710 N chr6 40209933 N DUP 27
SRR1766447.4273536 chr6 40209710 N chr6 40209933 N DUP 28
SRR1766448.7464201 chr6 40209594 N chr6 40209789 N DEL 22
SRR1766444.1954797 chr6 40209576 N chr6 40209771 N DEL 26
SRR1766443.8549389 chr6 40209602 N chr6 40209789 N DEL 25
SRR1766450.6976269 chr6 40209710 N chr6 40209933 N DUP 35
SRR1766454.7416014 chr6 40209710 N chr6 40209933 N DUP 33
SRR1766442.38069493 chr6 40209710 N chr6 40209933 N DUP 32
SRR1766474.4657954 chr6 40209710 N chr6 40209933 N DUP 29
SRR1766476.4536931 chr6 40209710 N chr6 40209933 N DUP 28
SRR1766461.10258966 chr6 40209699 N chr6 40209910 N DUP 22
SRR1766462.11185331 chr6 40209446 N chr6 40209799 N DEL 24
SRR1766453.1324498 chr6 40209446 N chr6 40209799 N DEL 24
SRR1766443.5327830 chr6 40209446 N chr6 40209799 N DEL 23
SRR1766443.2709190 chr6 40209581 N chr6 40209792 N DEL 27
SRR1766467.10408201 chr6 40209439 N chr6 40209792 N DEL 23
SRR1766482.5377961 chr6 40209297 N chr6 40209792 N DEL 25
SRR1766442.26986129 chr6 40209710 N chr6 40209933 N DUP 31
SRR1766444.2847076 chr6 40209789 N chr6 40209910 N DUP 27
SRR1766442.27163626 chr6 40209563 N chr6 40209800 N DEL 22
SRR1766463.2468135 chr6 40209605 N chr6 40209864 N DEL 28
SRR1766462.4603369 chr2 10015918 N chr2 10016004 N DUP 34
SRR1766442.6929645 chr2 10015632 N chr2 10015918 N DEL 20
SRR1766461.5928700 chr2 10015545 N chr2 10015918 N DEL 32
SRR1766444.5811458 chr2 10016098 N chr2 10016354 N DEL 22
SRR1766449.1832322 chr5 92251215 N chr5 92251326 N DUP 21
SRR1766451.4329725 chr15 21777066 N chr15 21777415 N DEL 25
SRR1766482.9682475 chr2 208177113 N chr2 208177164 N DEL 27
SRR1766469.7791650 chr2 208177089 N chr2 208177164 N DEL 21
SRR1766442.2128103 chr19 40349976 N chr19 40350279 N DEL 20
SRR1766446.6764419 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766472.4613969 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766458.3116698 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766466.1567353 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766476.854244 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766453.110206 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766468.7577578 chr3 111167155 N chr3 111167254 N DEL 24
SRR1766453.7906072 chr8 121201742 N chr8 121201797 N DUP 27
SRR1766466.5978198 chr8 121201742 N chr8 121201797 N DUP 31
SRR1766461.9745147 chr8 121201743 N chr8 121201798 N DUP 36
SRR1766473.10430545 chr8 121201731 N chr8 121201814 N DUP 37
SRR1766482.12682478 chr8 121201731 N chr8 121201814 N DUP 37
SRR1766442.30384333 chr8 121201731 N chr8 121201814 N DUP 36
SRR1766472.4290844 chr8 121201742 N chr8 121201797 N DUP 36
SRR1766479.7782704 chr8 121201731 N chr8 121201814 N DUP 38
SRR1766476.1120260 chr8 121201731 N chr8 121201814 N DUP 36
SRR1766442.10320318 chr8 121201731 N chr8 121201814 N DUP 36
SRR1766479.12075917 chr8 121201731 N chr8 121201814 N DUP 36
SRR1766484.3570631 chr8 121201742 N chr8 121201797 N DUP 23
SRR1766445.6162180 chr8 121201760 N chr8 121201851 N DUP 21
SRR1766442.32155005 chr8 121201742 N chr8 121201797 N DUP 23
SRR1766451.288703 chr8 121201731 N chr8 121201814 N DUP 34
SRR1766454.3139006 chr8 121201731 N chr8 121201814 N DUP 34
SRR1766464.1264448 chr8 121201742 N chr8 121201797 N DUP 36
SRR1766463.1769967 chr7 157994701 N chr7 157994819 N DEL 29
SRR1766481.5622972 chr7 157994701 N chr7 157994819 N DEL 30
SRR1766463.10420251 chr7 157994701 N chr7 157994819 N DEL 30
SRR1766468.1303758 chr7 157994657 N chr7 157994738 N DUP 24
SRR1766442.35192898 chr7 157994652 N chr7 157994733 N DUP 25
SRR1766462.881771 chr7 157994652 N chr7 157994733 N DUP 32
SRR1766478.1854747 chr7 157994652 N chr7 157994733 N DUP 24
SRR1766464.5066659 chr7 157994771 N chr7 157994852 N DUP 20
SRR1766483.9778397 chr7 157994771 N chr7 157994852 N DUP 25
SRR1766458.626563 chr7 157994701 N chr7 157994819 N DEL 30
SRR1766459.4770473 chr1 42324194 N chr1 42324285 N DEL 27
SRR1766486.692995 chr2 122274144 N chr2 122274269 N DEL 21
SRR1766467.1461203 chrX 62523742 N chrX 62524252 N DEL 25
SRR1766470.3183711 chr6 168044327 N chr6 168044789 N DEL 23
SRR1766485.7620708 chr1 154714107 N chr1 154714760 N DEL 22
SRR1766484.6011862 chr1 154714107 N chr1 154714760 N DEL 22
SRR1766460.8417822 chr1 154714117 N chr1 154714693 N DEL 25
SRR1766442.19833827 chr1 154714274 N chr1 154714331 N DEL 23
SRR1766455.3191781 chr1 154714297 N chr1 154714354 N DEL 29
SRR1766442.21178965 chr1 154714141 N chr1 154714587 N DUP 26
SRR1766446.6990697 chr1 154714457 N chr1 154714607 N DEL 27
SRR1766481.10293459 chr1 154714139 N chr1 154714587 N DUP 24
SRR1766456.140230 chr1 154714457 N chr1 154714607 N DEL 35
SRR1766467.10907432 chr1 154714134 N chr1 154714687 N DUP 26
SRR1766460.126957 chr1 154714655 N chr1 154714786 N DEL 27
SRR1766479.2708796 chr18 76587105 N chr18 76587412 N DEL 33
SRR1766455.5916173 chr18 76587139 N chr18 76587293 N DEL 33
SRR1766481.4038627 chr18 76587178 N chr18 76587332 N DEL 20
SRR1766456.3999652 chr18 76587048 N chr18 76587338 N DEL 30
SRR1766461.3207899 chr5 32158173 N chr5 32158287 N DUP 24
SRR1766483.5987532 chr13 108258355 N chr13 108258404 N DUP 25
SRR1766486.7066633 chr13 108258351 N chr13 108258400 N DUP 25
SRR1766465.4632427 chr13 108258351 N chr13 108258400 N DUP 25
SRR1766442.22260542 chr13 108258351 N chr13 108258400 N DUP 25
SRR1766469.18885 chr13 108258351 N chr13 108258400 N DUP 25
SRR1766455.1415730 chr13 108258351 N chr13 108258400 N DUP 27
SRR1766458.3779198 chr13 108258351 N chr13 108258400 N DUP 38
SRR1766459.1118596 chr13 108258351 N chr13 108258400 N DUP 20
SRR1766457.626318 chr13 108258351 N chr13 108258400 N DUP 24
SRR1766474.11674704 chr1 3502172 N chr1 3502250 N DUP 25
SRR1766448.97907 chr19 52554530 N chr19 52555035 N DEL 30
SRR1766456.2387469 chr19 52555013 N chr19 52555182 N DEL 25
SRR1766458.46167 chr19 52554544 N chr19 52555049 N DEL 30
SRR1766453.750168 chr6 1054124 N chr6 1054177 N DUP 23
SRR1766442.8735881 chr22 48757304 N chr22 48757589 N DUP 31
SRR1766485.7566056 chr22 48757461 N chr22 48757593 N DUP 32
SRR1766445.9601123 chr22 48757462 N chr22 48757594 N DUP 32
SRR1766470.9224590 chr22 48757461 N chr22 48757593 N DUP 32
SRR1766463.9759456 chr22 48757461 N chr22 48757593 N DUP 27
SRR1766450.234388 chr22 48757304 N chr22 48757508 N DUP 21
SRR1766478.11778193 chr22 48757304 N chr22 48757446 N DUP 23
SRR1766446.9710512 chr8 93833664 N chr8 93833999 N DEL 20
SRR1766442.27394378 chr18 29511893 N chr18 29511946 N DEL 22
SRR1766443.10079627 chr18 29511893 N chr18 29511946 N DEL 21
SRR1766447.730327 chr18 29512116 N chr18 29512199 N DUP 22
SRR1766486.6897880 chr18 29512102 N chr18 29512175 N DUP 20
SRR1766451.10200674 chr18 29512116 N chr18 29512199 N DUP 29
SRR1766476.1767158 chr18 29512133 N chr18 29512346 N DUP 21
SRR1766481.2297823 chr18 29512133 N chr18 29512346 N DUP 21
SRR1766442.28760933 chr18 29512204 N chr18 29512344 N DUP 27
SRR1766486.4476584 chr18 29512230 N chr18 29512344 N DUP 25
SRR1766450.1116268 chr18 29511666 N chr18 29512230 N DEL 20
SRR1766479.9912839 chr18 29511666 N chr18 29512230 N DEL 20
SRR1766442.8245711 chr18 29511666 N chr18 29512230 N DEL 20
SRR1766469.3902827 chr18 29511666 N chr18 29512230 N DEL 20
SRR1766481.11859953 chr18 29512199 N chr18 29512282 N DEL 26
SRR1766442.44756759 chr18 29512163 N chr18 29512282 N DEL 28
SRR1766454.325548 chr18 29512230 N chr18 29512344 N DUP 27
SRR1766442.42093179 chr4 162764161 N chr4 162764228 N DUP 22
SRR1766445.10545933 chr4 162764161 N chr4 162764228 N DUP 28
SRR1766446.4231808 chr4 162764120 N chr4 162764228 N DUP 30
SRR1766484.9703071 chr4 162764120 N chr4 162764228 N DUP 30
SRR1766445.6231410 chr4 162764160 N chr4 162764209 N DUP 37
SRR1766466.3922666 chr4 162764120 N chr4 162764228 N DUP 24
SRR1766476.10399494 chr4 162764120 N chr4 162764228 N DUP 24
SRR1766465.7415466 chr4 162764120 N chr4 162764228 N DUP 29
SRR1766476.10864049 chr4 162764120 N chr4 162764228 N DUP 29
SRR1766468.575116 chr4 162764160 N chr4 162764209 N DUP 34
SRR1766456.5541965 chr4 162764160 N chr4 162764209 N DUP 36
SRR1766464.10343395 chr4 162764160 N chr4 162764209 N DUP 36
SRR1766483.5105017 chr4 162764143 N chr4 162764201 N DEL 23
SRR1766446.4776360 chr4 162764143 N chr4 162764201 N DEL 21
SRR1766477.9642725 chr4 162764143 N chr4 162764201 N DEL 21
SRR1766462.59031 chr4 162764143 N chr4 162764201 N DEL 21
SRR1766443.1572423 chr4 162764143 N chr4 162764201 N DEL 23
SRR1766455.7585734 chr4 162764143 N chr4 162764201 N DEL 23
SRR1766442.33744957 chr20 64105723 N chr20 64105875 N DEL 20
SRR1766483.9561670 chr20 64105722 N chr20 64105874 N DEL 20
SRR1766461.8523351 chr20 64105722 N chr20 64105874 N DEL 20
SRR1766468.5538195 chr20 64105681 N chr20 64105875 N DEL 20
SRR1766482.5469074 chr3 77323092 N chr3 77323173 N DUP 20
SRR1766480.4069988 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766471.6636310 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766468.7840055 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766480.6578666 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766471.8305279 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766462.7983021 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766446.10526335 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766486.8071106 chr12 7197426 N chr12 7197528 N DUP 20
SRR1766442.17743676 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766467.8277990 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766483.7669952 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766483.7090183 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766464.2949238 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766462.11102186 chr12 7197464 N chr12 7197544 N DUP 27
SRR1766486.11792641 chr12 7197427 N chr12 7197580 N DUP 23
SRR1766478.3221258 chr12 7197427 N chr12 7197580 N DUP 28
SRR1766459.6053149 chr12 7197464 N chr12 7197544 N DUP 27
SRR1766460.4289330 chr12 7197484 N chr12 7197563 N DUP 28
SRR1766457.550630 chr12 7197464 N chr12 7197570 N DUP 31
SRR1766479.5202926 chr12 7197464 N chr12 7197570 N DUP 31
SRR1766467.8998667 chr12 7197482 N chr12 7197564 N DUP 25
SRR1766486.6579404 chr6 166824831 N chr6 166824926 N DEL 22
SRR1766467.7704282 chrY 6081085 N chrY 6081406 N DEL 21
SRR1766475.586435 chr10 16646073 N chr10 16646156 N DEL 23
SRR1766446.1990774 chr13 87990186 N chr13 87990243 N DEL 32
SRR1766462.1762920 chr13 87990186 N chr13 87990243 N DEL 36
SRR1766464.3248739 chr13 87990186 N chr13 87990243 N DEL 35
SRR1766486.10295875 chr8 142116246 N chr8 142116435 N DEL 21
SRR1766465.6279546 chr8 1698407 N chr8 1698698 N DEL 20
SRR1766461.6908107 chr8 1698752 N chr8 1698808 N DUP 22
SRR1766455.2025403 chr8 1698664 N chr8 1698808 N DUP 20
SRR1766447.5521092 chr8 1698709 N chr8 1698765 N DUP 22
SRR1766453.1875414 chr8 1698450 N chr8 1698798 N DEL 30
SRR1766480.4328314 chr18 78755872 N chr18 78756029 N DEL 25
SRR1766443.7223220 chr4 117740001 N chr4 117740063 N DUP 20
SRR1766486.714908 chr4 117740001 N chr4 117740063 N DUP 20
SRR1766481.1396643 chr4 117740001 N chr4 117740063 N DUP 26
SRR1766453.5765675 chr4 117740001 N chr4 117740063 N DUP 27
SRR1766485.2393910 chr4 117740001 N chr4 117740063 N DUP 34
SRR1766471.2332312 chr4 117740001 N chr4 117740063 N DUP 36
SRR1766448.1984575 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766442.113303 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766462.4751505 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766470.7062168 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766467.6169663 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766455.7778042 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766442.23983098 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766464.5262491 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766442.11958196 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766445.9433921 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766469.2490008 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766465.11141919 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766477.4403156 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766459.1191571 chr4 117740001 N chr4 117740063 N DUP 39
SRR1766458.3851732 chr4 117740226 N chr4 117740320 N DEL 24
SRR1766462.8081067 chr4 117740226 N chr4 117740320 N DEL 24
SRR1766484.9652404 chr4 117740226 N chr4 117740320 N DEL 26
SRR1766458.1000470 chr4 117740226 N chr4 117740320 N DEL 26
SRR1766467.607608 chr4 117740226 N chr4 117740320 N DEL 26
SRR1766468.7713097 chr4 117740226 N chr4 117740320 N DEL 29
SRR1766474.1401520 chr4 117740226 N chr4 117740320 N DEL 30
SRR1766462.5862362 chr4 117740226 N chr4 117740320 N DEL 30
SRR1766464.4587641 chr4 117740226 N chr4 117740320 N DEL 31
SRR1766464.6645833 chr4 117740226 N chr4 117740320 N DEL 32
SRR1766450.4606567 chr16 89342033 N chr16 89342206 N DUP 20
SRR1766467.11546382 chr16 89342136 N chr16 89342227 N DEL 38
SRR1766448.733517 chr16 89342136 N chr16 89342227 N DEL 25
SRR1766448.8949338 chr16 89342136 N chr16 89342227 N DEL 23
SRR1766442.21173843 chr8 123315143 N chr8 123315495 N DEL 20
SRR1766456.4660246 chr8 123315143 N chr8 123315495 N DEL 20
SRR1766446.4033195 chr8 123315143 N chr8 123315495 N DEL 20
SRR1766453.9408663 chr8 123315184 N chr8 123315585 N DEL 24
SRR1766458.1257881 chrX 40616950 N chrX 40617023 N DUP 32
SRR1766475.768835 chrX 818492 N chrX 818546 N DEL 22
SRR1766476.5977634 chrX 818457 N chrX 818546 N DEL 20
SRR1766484.3957404 chrX 818457 N chrX 818546 N DEL 23
SRR1766455.2207311 chrX 818457 N chrX 818546 N DEL 20
SRR1766449.4400899 chrX 818457 N chrX 818546 N DEL 22
SRR1766484.12259432 chrX 818457 N chrX 818546 N DEL 24
SRR1766468.5777039 chr22 42087670 N chr22 42087976 N DEL 26
SRR1766473.8208453 chr22 42087669 N chr22 42088275 N DEL 20
SRR1766458.5155559 chr22 42088023 N chr22 42088324 N DEL 36
SRR1766466.11283389 chr9 20417146 N chr9 20417459 N DEL 20
SRR1766480.8641988 chr22 46194965 N chr22 46195295 N DEL 20
SRR1766442.46038382 chr22 46194970 N chr22 46195300 N DEL 20
SRR1766481.4088628 chr10 7526840 N chr10 7526973 N DUP 21
SRR1766478.7249718 chr10 7526840 N chr10 7526973 N DUP 20
SRR1766453.7469241 chr10 7526840 N chr10 7526973 N DUP 20
SRR1766483.3971877 chr10 92393448 N chr10 92393539 N DEL 25
SRR1766461.9158422 chr14 101245290 N chr14 101245651 N DEL 35
SRR1766446.311057 chr14 101245939 N chr14 101246622 N DUP 28
SRR1766460.4815622 chr14 101245373 N chr14 101246724 N DEL 27
SRR1766458.7111845 chr14 101245334 N chr14 101245425 N DEL 23
SRR1766468.7765869 chr14 101245356 N chr14 101245735 N DEL 24
SRR1766486.5330697 chr14 101246382 N chr14 101246707 N DEL 20
SRR1766481.1297127 chr14 101245451 N chr14 101246100 N DEL 20
SRR1766483.9148776 chr14 101245964 N chr14 101246379 N DEL 20
SRR1766482.5168333 chr14 101245478 N chr14 101245533 N DEL 25
SRR1766442.42666224 chr14 101245460 N chr14 101246379 N DEL 29
SRR1766444.5923801 chr14 101245496 N chr14 101245821 N DEL 24
SRR1766486.114319 chr14 101245460 N chr14 101246379 N DEL 31
SRR1766445.1439541 chr14 101245327 N chr14 101245470 N DUP 25
SRR1766463.7734475 chr14 101245282 N chr14 101245497 N DUP 21
SRR1766454.599539 chr14 101245560 N chr14 101245939 N DEL 20
SRR1766478.9781159 chr14 101245597 N chr14 101245904 N DEL 20
SRR1766478.6037459 chr14 101245362 N chr14 101245633 N DEL 25
SRR1766482.415829 chr14 101245636 N chr14 101245887 N DUP 20
SRR1766470.1895312 chr14 101245318 N chr14 101245695 N DUP 20
SRR1766477.2542897 chr14 101245633 N chr14 101245884 N DUP 20
SRR1766477.1493530 chr14 101245308 N chr14 101245633 N DEL 20
SRR1766479.6759241 chr14 101245293 N chr14 101245654 N DEL 20
SRR1766453.6240820 chr14 101245273 N chr14 101245704 N DUP 20
SRR1766442.33690140 chr14 101245374 N chr14 101245717 N DEL 26
SRR1766465.3000192 chr14 101245351 N chr14 101246738 N DEL 30
SRR1766484.10457121 chr14 101245374 N chr14 101245735 N DEL 30
SRR1766484.5382012 chr14 101245776 N chr14 101245831 N DEL 20
SRR1766447.9871520 chr14 101245370 N chr14 101245749 N DEL 26
SRR1766482.5168333 chr14 101245370 N chr14 101246487 N DEL 25
SRR1766478.1825873 chr14 101245488 N chr14 101245831 N DEL 20
SRR1766448.7476190 chr14 101245831 N chr14 101245884 N DUP 22
SRR1766481.5165580 chr14 101245317 N chr14 101245892 N DUP 22
SRR1766485.7749809 chr14 101245821 N chr14 101245892 N DUP 20
SRR1766478.11319565 chr14 101245293 N chr14 101245834 N DEL 20
SRR1766457.6100005 chr14 101245831 N chr14 101245884 N DUP 25
SRR1766484.2565051 chr14 101245831 N chr14 101245992 N DUP 24
SRR1766450.2080379 chr14 101245487 N chr14 101246100 N DEL 20
SRR1766442.5700407 chr14 101245362 N chr14 101245831 N DEL 22
SRR1766484.7193371 chr14 101246136 N chr14 101246605 N DEL 25
SRR1766466.7587906 chr14 101245478 N chr14 101245533 N DEL 20
SRR1766460.2051043 chr14 101245327 N chr14 101246046 N DUP 20
SRR1766446.2915964 chr14 101245831 N chr14 101246154 N DUP 30
SRR1766451.3372057 chr14 101245274 N chr14 101246173 N DUP 20
SRR1766471.3573507 chr14 101245896 N chr14 101246203 N DEL 20
SRR1766471.10486227 chr14 101245271 N chr14 101245756 N DUP 20
SRR1766479.5642890 chr14 101245299 N chr14 101246270 N DUP 20
SRR1766486.5168337 chr14 101245525 N chr14 101245902 N DUP 20
SRR1766452.9309309 chr14 101245273 N chr14 101246298 N DUP 20
SRR1766457.7217813 chr14 101246101 N chr14 101246334 N DUP 25
SRR1766450.8366300 chr14 101245478 N chr14 101246217 N DEL 25
SRR1766460.1657224 chr14 101245273 N chr14 101246352 N DUP 20
SRR1766475.1637672 chr14 101245831 N chr14 101246280 N DUP 20
SRR1766475.10583976 chr14 101245866 N chr14 101246101 N DEL 20
SRR1766449.1277676 chr14 101245998 N chr14 101246485 N DEL 25
SRR1766486.699950 chr14 101245299 N chr14 101246452 N DEL 20
SRR1766442.704320 chr14 101245350 N chr14 101246485 N DEL 30
SRR1766461.10770513 chr14 101245271 N chr14 101246242 N DUP 23
SRR1766485.980861 chr14 101245361 N chr14 101246604 N DEL 25
SRR1766465.4071350 chr14 101246559 N chr14 101246666 N DUP 20
SRR1766462.2601057 chr14 101245496 N chr14 101246091 N DEL 20
SRR1766455.8583754 chr14 101246135 N chr14 101246782 N DUP 20
SRR1766466.8118570 chr14 101245464 N chr14 101246689 N DEL 20
SRR1766475.10771606 chr14 101245921 N chr14 101246046 N DUP 20
SRR1766453.10345893 chr14 101246026 N chr14 101246819 N DEL 20
SRR1766474.7532084 chr2 60467296 N chr2 60467598 N DUP 20
SRR1766480.4112742 chr2 60467297 N chr2 60467611 N DUP 21
SRR1766458.1886098 chr2 60467291 N chr2 60467530 N DUP 20
SRR1766459.3303569 chr2 60467347 N chr2 60467879 N DEL 23
SRR1766445.10213320 chr2 60467331 N chr2 60467893 N DEL 29
SRR1766442.3002635 chr2 60467226 N chr2 60467966 N DUP 23
SRR1766455.9636460 chr2 60467346 N chr2 60468262 N DEL 20
SRR1766480.2776584 chr17 402226 N chr17 402302 N DUP 21
SRR1766460.158631 chr1 83013698 N chr1 83013789 N DEL 29
SRR1766483.9963672 chr1 83013698 N chr1 83013789 N DEL 22
SRR1766464.2046669 chr6 158157029 N chr6 158157108 N DUP 27
SRR1766454.5677670 chr12 122163820 N chr12 122164123 N DEL 25
SRR1766479.6732906 chr12 122164200 N chr12 122164798 N DEL 20
SRR1766475.7100167 chr9 9845155 N chr9 9845230 N DEL 24
SRR1766465.9503357 chr9 9845167 N chr9 9845242 N DEL 27
SRR1766479.13507727 chr7 34129758 N chr7 34129809 N DEL 22
SRR1766471.5341137 chr12 14179750 N chr12 14179989 N DUP 24
SRR1766470.1907208 chr12 14179750 N chr12 14179989 N DUP 24
SRR1766443.1479011 chr12 14179750 N chr12 14179989 N DUP 24
SRR1766463.9554293 chr15 97641268 N chr15 97641333 N DUP 28
SRR1766464.1175433 chr15 97641268 N chr15 97641333 N DUP 34
SRR1766461.10816161 chr15 97641268 N chr15 97641333 N DUP 28
SRR1766459.5931635 chr15 97641268 N chr15 97641333 N DUP 30
SRR1766442.22567980 chr15 97641268 N chr15 97641333 N DUP 29
SRR1766444.1225838 chr6 82306996 N chr6 82307055 N DEL 24
SRR1766442.22455973 chr6 82306996 N chr6 82307055 N DEL 21
SRR1766459.11232537 chr6 82306998 N chr6 82307077 N DEL 22
SRR1766448.10210807 chr6 82306998 N chr6 82307077 N DEL 22
SRR1766480.2123825 chr12 131327152 N chr12 131327394 N DEL 20
SRR1766478.2037580 chr12 131327103 N chr12 131327197 N DUP 22
SRR1766442.10665047 chr12 131327200 N chr12 131327347 N DEL 25
SRR1766465.8884821 chr12 132518428 N chr12 132518559 N DEL 36
SRR1766452.10646644 chrX 121079468 N chrX 121079768 N DEL 30
SRR1766483.259294 chr3 180873904 N chr3 180874227 N DEL 20
SRR1766471.6389135 chr7 14471315 N chr7 14471407 N DEL 20
SRR1766476.4369637 chr7 14471315 N chr7 14471407 N DEL 21
SRR1766459.2282115 chr7 14471315 N chr7 14471407 N DEL 26
SRR1766449.8432411 chr7 14471315 N chr7 14471469 N DEL 28
SRR1766454.1892234 chr7 14471315 N chr7 14471407 N DEL 25
SRR1766472.6711196 chr7 14471315 N chr7 14471407 N DEL 28
SRR1766442.12888009 chr7 14471315 N chr7 14471407 N DEL 24
SRR1766465.5927457 chr7 14471315 N chr7 14471407 N DEL 24
SRR1766450.3889651 chr7 14471315 N chr7 14471407 N DEL 24
SRR1766442.19631537 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766464.3823515 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766442.19519932 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766483.1302022 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766445.5578674 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766465.3333568 chr12 78626252 N chr12 78626307 N DUP 31
SRR1766445.6536061 chr17 18000173 N chr17 18000510 N DEL 27
SRR1766446.2399663 chr17 891839 N chr17 892061 N DEL 21
SRR1766476.4696548 chr17 891893 N chr17 892225 N DEL 20
SRR1766482.11089384 chr17 891874 N chr17 892206 N DEL 20
SRR1766459.2193542 chr17 891904 N chr17 892234 N DUP 20
SRR1766458.3689918 chr17 891911 N chr17 892169 N DEL 20
SRR1766486.2786602 chr17 891911 N chr17 892169 N DEL 20
SRR1766482.2243559 chr17 891913 N chr17 892208 N DEL 23
SRR1766449.1953732 chr17 891913 N chr17 892208 N DEL 20
SRR1766456.1177652 chr17 891913 N chr17 892208 N DEL 20
SRR1766467.4831609 chr17 891913 N chr17 892208 N DEL 20
SRR1766460.10169943 chr4 11191938 N chr4 11192036 N DUP 20
SRR1766447.460340 chr10 60240162 N chr10 60240282 N DUP 31
SRR1766457.6485003 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766461.10565373 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766451.8173222 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766443.2558803 chr10 60240271 N chr10 60240402 N DUP 20
SRR1766442.32666096 chr6 84395673 N chr6 84395763 N DUP 21
SRR1766467.11104608 chr6 84395673 N chr6 84395755 N DUP 21
SRR1766458.6309674 chr9 134977517 N chr9 134977632 N DEL 26
SRR1766442.14526898 chr8 58301684 N chr8 58301733 N DUP 20
SRR1766442.25935094 chr8 58301684 N chr8 58301733 N DUP 28
SRR1766448.3398217 chr8 58301684 N chr8 58301733 N DUP 28
SRR1766466.9953406 chr12 51858512 N chr12 51858817 N DEL 35
SRR1766481.589331 chr10 54332395 N chr10 54332497 N DUP 28
SRR1766442.46601613 chr10 54332451 N chr10 54332517 N DUP 28
SRR1766443.5132830 chr10 54332451 N chr10 54332517 N DUP 28
SRR1766452.1402192 chr10 54332451 N chr10 54332517 N DUP 28
SRR1766477.11894468 chr10 54332415 N chr10 54332481 N DUP 38
SRR1766479.1053038 chr10 54332415 N chr10 54332481 N DUP 38
SRR1766454.6419540 chr10 54332415 N chr10 54332517 N DUP 24
SRR1766484.4795239 chr10 54332415 N chr10 54332517 N DUP 26
SRR1766466.5574371 chr10 54332395 N chr10 54332502 N DUP 20
SRR1766457.2433659 chr10 54332415 N chr10 54332517 N DUP 30
SRR1766452.2995561 chr10 54332415 N chr10 54332481 N DUP 24
SRR1766456.4088960 chr10 54332415 N chr10 54332517 N DUP 23
SRR1766483.1231495 chr10 54332415 N chr10 54332517 N DUP 24
SRR1766450.9512239 chr10 54332415 N chr10 54332517 N DUP 25
SRR1766459.1646041 chr6 170114229 N chr6 170114318 N DUP 24
SRR1766450.5150588 chr6 170114229 N chr6 170114318 N DUP 24
SRR1766473.1731086 chr6 170114229 N chr6 170114318 N DUP 23
SRR1766465.10950306 chr15 101764198 N chr15 101764634 N DEL 20
SRR1766462.8782756 chr2 240812862 N chr2 240813161 N DUP 22
SRR1766469.6886259 chr2 240813030 N chr2 240813181 N DUP 27
SRR1766442.23769213 chr2 240813030 N chr2 240813105 N DUP 22
SRR1766464.2540435 chr2 240813053 N chr2 240813185 N DUP 22
SRR1766460.7765759 chr2 240813030 N chr2 240813105 N DUP 21
SRR1766465.11194010 chr2 240813025 N chr2 240813100 N DUP 20
SRR1766480.4629870 chr6 121497528 N chr6 121497841 N DEL 32
SRR1766464.8669415 chr1 222138942 N chr1 222139039 N DUP 22
SRR1766442.23570587 chr1 222138942 N chr1 222139039 N DUP 27
SRR1766475.1358042 chr1 222138977 N chr1 222139042 N DEL 23
SRR1766449.5092166 chr1 222138977 N chr1 222139042 N DEL 21
SRR1766481.5569726 chr1 248671537 N chr1 248671895 N DEL 24
SRR1766480.3023694 chr1 248671541 N chr1 248672154 N DEL 20
SRR1766470.10764973 chr1 248671698 N chr1 248671750 N DEL 20
SRR1766477.7562770 chr1 248671698 N chr1 248671750 N DEL 20
SRR1766444.3160027 chr1 248671700 N chr1 248671854 N DEL 25
SRR1766463.1988046 chr1 248671700 N chr1 248671854 N DEL 20
SRR1766453.3847903 chr3 79771313 N chr3 79771366 N DEL 23
SRR1766452.10372461 chr3 79771313 N chr3 79771366 N DEL 28
SRR1766476.6189739 chr3 79771313 N chr3 79771366 N DEL 28
SRR1766448.3725473 chr3 79771313 N chr3 79771366 N DEL 28
SRR1766462.7069828 chr4 180390417 N chr4 180390886 N DEL 22
SRR1766443.6654511 chr4 180390402 N chr4 180390477 N DUP 23
SRR1766484.7957851 chr4 180390530 N chr4 180391208 N DUP 20
SRR1766444.2556506 chr4 180390576 N chr4 180390639 N DUP 21
SRR1766447.8760417 chr4 180390576 N chr4 180391031 N DUP 22
SRR1766479.139386 chr4 180390522 N chr4 180390607 N DUP 20
SRR1766453.53516 chr4 180390638 N chr4 180390745 N DUP 29
SRR1766453.11134061 chr4 180390545 N chr4 180390638 N DUP 20
SRR1766461.3163747 chr4 180390538 N chr4 180390646 N DUP 21
SRR1766449.9336359 chr4 180390676 N chr4 180391146 N DEL 22
SRR1766472.3801090 chr4 180390538 N chr4 180390646 N DUP 22
SRR1766471.5533460 chr4 180390538 N chr4 180390646 N DUP 22
SRR1766455.8286378 chr4 180390640 N chr4 180390735 N DUP 20
SRR1766442.42794430 chr4 180390640 N chr4 180390735 N DUP 20
SRR1766471.7783539 chr4 180390637 N chr4 180391012 N DEL 25
SRR1766449.1749899 chr4 180390591 N chr4 180391050 N DUP 21
SRR1766454.6360892 chr4 180390935 N chr4 180391050 N DUP 21
SRR1766464.9414523 chr4 180390608 N chr4 180391214 N DEL 28
SRR1766449.1214453 chr4 180391059 N chr4 180391181 N DEL 29
SRR1766442.47067820 chr4 180390615 N chr4 180391224 N DEL 37
SRR1766482.5674698 chr4 180390607 N chr4 180391213 N DEL 23
SRR1766473.8686144 chr4 180390607 N chr4 180391213 N DEL 23
SRR1766467.1808429 chr4 180390607 N chr4 180391213 N DEL 22
SRR1766454.6324027 chr4 180390615 N chr4 180391224 N DEL 34
SRR1766449.1749899 chr4 180390615 N chr4 180391224 N DEL 34
SRR1766442.26071044 chr4 180390615 N chr4 180391224 N DEL 33
SRR1766460.7594419 chr4 180390607 N chr4 180391213 N DEL 20
SRR1766469.2793875 chr4 180390421 N chr4 180391224 N DEL 23
SRR1766458.4247491 chr4 180390421 N chr4 180391224 N DEL 23
SRR1766453.10166399 chr4 180390421 N chr4 180391224 N DEL 23
SRR1766478.6264161 chr6 162010661 N chr6 162010762 N DEL 28
SRR1766476.7743555 chr6 162010663 N chr6 162010726 N DEL 32
SRR1766469.8231917 chr6 162010640 N chr6 162010809 N DUP 23
SRR1766465.7360623 chr6 162011300 N chr6 162011378 N DUP 34
SRR1766469.10602117 chr6 162011300 N chr6 162011378 N DUP 34
SRR1766452.5136227 chr6 162011290 N chr6 162011365 N DUP 23
SRR1766448.4306549 chr6 162011471 N chr6 162011656 N DEL 30
SRR1766463.1801395 chr6 162011471 N chr6 162011656 N DEL 27
SRR1766480.7989608 chr6 162011471 N chr6 162011656 N DEL 27
SRR1766449.9442248 chr6 162011431 N chr6 162011656 N DEL 21
SRR1766443.10049907 chr21 44592020 N chr21 44592376 N DUP 35
SRR1766471.8305933 chr21 44592020 N chr21 44592376 N DUP 35
SRR1766485.10431269 chr21 44592020 N chr21 44592376 N DUP 25
SRR1766449.4765488 chr21 44592020 N chr21 44592376 N DUP 24
SRR1766442.35438280 chr21 44592020 N chr21 44592376 N DUP 30
SRR1766465.1358823 chr10 62370476 N chr10 62370609 N DEL 25
SRR1766444.5133737 chr10 62370456 N chr10 62370578 N DEL 31
SRR1766481.5667546 chr10 62370448 N chr10 62370628 N DEL 33
SRR1766483.2472541 chr10 62370448 N chr10 62370628 N DEL 36
SRR1766468.4425924 chr10 62370487 N chr10 62370602 N DEL 35
SRR1766476.5322532 chr10 62370607 N chr10 62371260 N DUP 31
SRR1766473.2857913 chr10 62370584 N chr10 62371255 N DUP 26
SRR1766471.9827554 chr10 62370750 N chr10 62370828 N DUP 22
SRR1766475.1761349 chr10 62370750 N chr10 62370828 N DUP 24
SRR1766453.874456 chr10 62370750 N chr10 62370828 N DUP 25
SRR1766477.3191317 chr10 62371045 N chr10 62371435 N DUP 27
SRR1766450.6102635 chr10 62371037 N chr10 62371190 N DUP 25
SRR1766449.9409974 chr10 62371128 N chr10 62371264 N DUP 29
SRR1766466.8289641 chr10 62371128 N chr10 62371264 N DUP 28
SRR1766455.4451455 chr10 62371128 N chr10 62371264 N DUP 25
SRR1766462.11124359 chr10 62371209 N chr10 62371293 N DUP 36
SRR1766464.7645344 chr10 62371128 N chr10 62371264 N DUP 34
SRR1766450.2799415 chr10 62371128 N chr10 62371264 N DUP 33
SRR1766460.3236897 chr10 62371200 N chr10 62371302 N DUP 26
SRR1766460.11272820 chr10 62371209 N chr10 62371293 N DUP 35
SRR1766465.4221373 chr10 62371209 N chr10 62371293 N DUP 35
SRR1766458.386574 chr10 62371209 N chr10 62371293 N DUP 35
SRR1766447.1331450 chr10 62371209 N chr10 62371293 N DUP 36
SRR1766463.2059416 chr10 62370659 N chr10 62371381 N DEL 20
SRR1766471.10937371 chr10 62371227 N chr10 62371449 N DUP 27
SRR1766476.10880071 chr10 62371227 N chr10 62371449 N DUP 27
SRR1766481.5366256 chr10 62371419 N chr10 62371509 N DUP 20
SRR1766485.6959853 chr10 62371419 N chr10 62371509 N DUP 25
SRR1766466.186680 chr10 62371362 N chr10 62371499 N DEL 20
SRR1766473.389348 chr10 62371367 N chr10 62371522 N DEL 21
SRR1766442.35009943 chr10 62371367 N chr10 62371522 N DEL 21
SRR1766460.11272820 chr10 62371367 N chr10 62371522 N DEL 21
SRR1766444.3315944 chr10 62371368 N chr10 62371523 N DEL 21
SRR1766442.13338086 chr9 89254496 N chr9 89254617 N DEL 20
SRR1766474.1220066 chr9 89254491 N chr9 89254612 N DEL 20
SRR1766444.525149 chr9 89254425 N chr9 89254483 N DEL 20
SRR1766477.9737244 chr9 89254418 N chr9 89254660 N DEL 30
SRR1766468.4967917 chr3 101891496 N chr3 101891710 N DEL 27
SRR1766471.4290421 chr13 83380731 N chr13 83380782 N DEL 21
SRR1766463.9696539 chr13 83380731 N chr13 83380782 N DEL 27
SRR1766484.1831171 chr21 41806228 N chr21 41806665 N DUP 27
SRR1766482.360597 chr21 41806361 N chr21 41806541 N DUP 21
SRR1766451.1777787 chr21 41806230 N chr21 41806599 N DUP 20
SRR1766453.5408994 chr21 41806302 N chr21 41806454 N DEL 22
SRR1766442.16985810 chr21 41806333 N chr21 41806521 N DEL 21
SRR1766449.3083375 chr21 41806168 N chr21 41806317 N DUP 26
SRR1766473.9285030 chr21 41806421 N chr21 41806814 N DUP 20
SRR1766465.8040727 chr21 41806341 N chr21 41806454 N DEL 20
SRR1766450.1600464 chr21 41806218 N chr21 41806288 N DEL 20
SRR1766467.6563996 chr21 41806396 N chr21 41806753 N DEL 23
SRR1766473.11526555 chr21 41689406 N chr21 41689463 N DEL 23
SRR1766448.2749749 chr21 41689413 N chr21 41689470 N DEL 30
SRR1766454.7733584 chr21 41689406 N chr21 41689463 N DEL 30
SRR1766442.29266828 chr1 143252863 N chr1 143252933 N DUP 31
SRR1766479.2922720 chr5 43032078 N chr5 43032199 N DUP 30
SRR1766448.7722582 chr5 43032027 N chr5 43032211 N DUP 30
SRR1766463.9215058 chr5 43032090 N chr5 43032148 N DEL 27
SRR1766450.10915952 chr5 43032027 N chr5 43032211 N DUP 31
SRR1766469.6876778 chr5 43032027 N chr5 43032211 N DUP 31
SRR1766453.1629404 chr5 43032027 N chr5 43032211 N DUP 33
SRR1766483.7341588 chr5 43032027 N chr5 43032211 N DUP 33
SRR1766446.8876971 chr5 43032189 N chr5 43032295 N DUP 27
SRR1766448.10120210 chr5 43032181 N chr5 43032262 N DUP 21
SRR1766449.6650428 chr5 43032189 N chr5 43032295 N DUP 24
SRR1766461.8829494 chr5 43032189 N chr5 43032295 N DUP 29
SRR1766475.7592665 chr5 43032181 N chr5 43032262 N DUP 23
SRR1766479.8454088 chr5 43032407 N chr5 43032458 N DEL 29
SRR1766473.7931566 chr5 43032407 N chr5 43032458 N DEL 31
SRR1766476.5470935 chr5 43032407 N chr5 43032458 N DEL 31
SRR1766448.3464580 chr5 43032166 N chr5 43032447 N DUP 24
SRR1766476.3704795 chr5 43032125 N chr5 43032414 N DUP 29
SRR1766453.3669188 chr5 43032367 N chr5 43032450 N DEL 32
SRR1766479.11598357 chr5 43032462 N chr5 43032526 N DUP 35
SRR1766474.191719 chr5 43032462 N chr5 43032526 N DUP 29
SRR1766454.10361147 chr18 57510089 N chr18 57510405 N DEL 25
SRR1766482.3349832 chr18 57510089 N chr18 57510405 N DEL 25
SRR1766442.27638210 chr18 57510089 N chr18 57510405 N DEL 25
SRR1766449.8983745 chr18 57510089 N chr18 57510405 N DEL 25
SRR1766450.646054 chr18 57510102 N chr18 57510418 N DEL 29
SRR1766467.5930255 chr18 57510089 N chr18 57510405 N DEL 30
SRR1766485.3130853 chr18 57510089 N chr18 57510405 N DEL 31
SRR1766455.4905559 chr18 57510089 N chr18 57510405 N DEL 38
SRR1766442.21132551 chr4 1828648 N chr4 1828701 N DEL 27
SRR1766442.11419759 chr4 1828648 N chr4 1828701 N DEL 21
SRR1766467.2018974 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766447.90772 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766471.5742663 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766467.1640808 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766442.22141324 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766478.11147337 chr1 189818463 N chr1 189818544 N DEL 32
SRR1766480.7377951 chr1 189818463 N chr1 189818544 N DEL 34
SRR1766442.23091358 chr1 189818463 N chr1 189818544 N DEL 34
SRR1766447.8843032 chr1 189818463 N chr1 189818544 N DEL 26
SRR1766479.12461066 chr1 189818463 N chr1 189818544 N DEL 21
SRR1766459.8411973 chr1 189818463 N chr1 189818544 N DEL 25
SRR1766474.10036292 chr1 189818463 N chr1 189818544 N DEL 28
SRR1766478.7644474 chr1 189818463 N chr1 189818544 N DEL 21
SRR1766476.10166012 chr7 156439918 N chr7 156440012 N DUP 20
SRR1766465.7270031 chr1 248841102 N chr1 248841157 N DEL 20
SRR1766467.6717490 chr5 10346474 N chr5 10346553 N DEL 38
SRR1766483.7742663 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766483.2867780 chr5 10346474 N chr5 10346553 N DEL 35
SRR1766476.6734492 chr5 10346474 N chr5 10346553 N DEL 35
SRR1766447.1785407 chr5 10347422 N chr5 10347479 N DUP 20
SRR1766466.1535782 chr5 10347096 N chr5 10347406 N DEL 20
SRR1766442.30459796 chr5 10346474 N chr5 10346553 N DEL 24
SRR1766447.1632621 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766468.8046972 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766442.17812002 chr5 10346474 N chr5 10346553 N DEL 38
SRR1766442.4704186 chr5 10347117 N chr5 10347398 N DEL 21
SRR1766457.5205264 chr5 10347422 N chr5 10347479 N DUP 21
SRR1766478.4509846 chr5 10346474 N chr5 10346553 N DEL 38
SRR1766443.243909 chr5 10346474 N chr5 10346553 N DEL 22
SRR1766483.5677680 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766472.1814641 chr5 10346474 N chr5 10346553 N DEL 38
SRR1766470.4139289 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766478.546252 chr19 9948187 N chr19 9948492 N DEL 33
SRR1766459.9770674 chr13 62019547 N chr13 62019606 N DEL 25
SRR1766462.9835446 chr13 62019547 N chr13 62019606 N DEL 29
SRR1766470.214716 chr13 62019547 N chr13 62019606 N DEL 27
SRR1766481.10670481 chr13 62019789 N chr13 62019848 N DUP 30
SRR1766456.6025753 chr13 62019789 N chr13 62019848 N DUP 27
SRR1766453.6644475 chr13 62019789 N chr13 62019848 N DUP 27
SRR1766469.7787499 chr13 62019789 N chr13 62019848 N DUP 32
SRR1766442.11096501 chr14 56355314 N chr14 56355425 N DUP 23
SRR1766476.4309794 chr14 56355314 N chr14 56355425 N DUP 24
SRR1766466.86738 chr14 56355314 N chr14 56355425 N DUP 23
SRR1766442.352658 chr14 56355331 N chr14 56355452 N DEL 20
SRR1766443.4673862 chr14 56355331 N chr14 56355452 N DEL 20
SRR1766445.8577450 chr14 56355331 N chr14 56355452 N DEL 20
SRR1766476.8144751 chr14 56355331 N chr14 56355452 N DEL 20
SRR1766479.7700020 chr8 29667260 N chr8 29667315 N DUP 21
SRR1766470.7687355 chr16 75059351 N chr16 75059403 N DUP 20
SRR1766485.3761545 chr10 15149605 N chr10 15149706 N DUP 24
SRR1766463.1853415 chr10 15149592 N chr10 15149657 N DUP 29
SRR1766453.3546593 chr10 15149592 N chr10 15149657 N DUP 26
SRR1766458.7380679 chr10 15149577 N chr10 15149738 N DUP 25
SRR1766457.6195757 chr7 61903967 N chr7 61904479 N DUP 20
SRR1766467.7554517 chr7 61904411 N chr7 61904927 N DEL 30
SRR1766477.3996881 chr9 134422431 N chr9 134422760 N DEL 20
SRR1766456.1207086 chr9 136308524 N chr9 136308782 N DEL 26
SRR1766445.4657924 chr19 14002233 N chr19 14002583 N DEL 30
SRR1766474.10648682 chr10 100525783 N chr10 100525866 N DUP 23
SRR1766454.10202566 chr20 7435687 N chr20 7435800 N DUP 21
SRR1766461.585810 chr20 7435687 N chr20 7435800 N DUP 21
SRR1766475.5692948 chr20 7435687 N chr20 7435800 N DUP 21
SRR1766453.5504645 chr20 7435687 N chr20 7435800 N DUP 21
SRR1766482.11599982 chr3 184414763 N chr3 184414888 N DEL 25
SRR1766459.6091257 chrX 532358 N chrX 532698 N DUP 25
SRR1766461.6522231 chrX 532736 N chrX 532905 N DEL 20
SRR1766477.8092036 chrX 532736 N chrX 532905 N DEL 20
SRR1766442.31760687 chrX 532358 N chrX 532698 N DUP 25
SRR1766470.10824691 chrX 532736 N chrX 532905 N DEL 20
SRR1766457.9194010 chrX 532736 N chrX 532905 N DEL 20
SRR1766442.4712355 chrX 532736 N chrX 532905 N DEL 20
SRR1766448.7771131 chrX 532736 N chrX 532905 N DEL 20
SRR1766460.9147976 chrX 532492 N chrX 532846 N DEL 21
SRR1766459.408763 chrX 532492 N chrX 532846 N DEL 25
SRR1766464.5201002 chrX 532334 N chrX 532489 N DUP 38
SRR1766477.4200360 chrX 532358 N chrX 532698 N DUP 25
SRR1766447.6321340 chrX 532358 N chrX 532698 N DUP 25
SRR1766470.6796442 chrX 532358 N chrX 532698 N DUP 25
SRR1766442.45090361 chrX 532358 N chrX 532698 N DUP 25
SRR1766448.8150322 chrX 532358 N chrX 532698 N DUP 25
SRR1766450.3143119 chrX 532358 N chrX 532698 N DUP 25
SRR1766474.4455774 chrX 532358 N chrX 532698 N DUP 25
SRR1766479.12130205 chrX 532358 N chrX 532698 N DUP 30
SRR1766484.10425771 chrX 532358 N chrX 532698 N DUP 30
SRR1766483.2085544 chrX 532358 N chrX 532698 N DUP 31
SRR1766485.8417833 chrX 532358 N chrX 532698 N DUP 31
SRR1766443.9657364 chrX 532358 N chrX 532698 N DUP 32
SRR1766442.34448767 chrX 532358 N chrX 532698 N DUP 32
SRR1766459.7002795 chrX 532814 N chrX 532984 N DUP 21
SRR1766478.9997886 chrX 532846 N chrX 533001 N DUP 27
SRR1766471.11981734 chrX 532846 N chrX 533001 N DUP 27
SRR1766472.6611511 chrX 532846 N chrX 533001 N DUP 27
SRR1766476.9652760 chrX 532814 N chrX 532984 N DUP 21
SRR1766483.9362901 chrX 532814 N chrX 532984 N DUP 21
SRR1766457.624091 chrX 532846 N chrX 533001 N DUP 27
SRR1766486.9501071 chrX 532814 N chrX 532984 N DUP 21
SRR1766468.7416564 chrX 532846 N chrX 533001 N DUP 24
SRR1766469.2266229 chrX 532846 N chrX 533001 N DUP 24
SRR1766442.17972795 chrX 532814 N chrX 532987 N DUP 21
SRR1766452.9736373 chrX 532358 N chrX 532698 N DUP 28
SRR1766485.7632539 chrX 532736 N chrX 532905 N DEL 23
SRR1766465.10786183 chrX 532736 N chrX 532905 N DEL 20
SRR1766449.5255823 chrX 532736 N chrX 532905 N DEL 20
SRR1766477.11445418 chrX 532846 N chrX 533001 N DUP 33
SRR1766481.7843412 chrX 532846 N chrX 533001 N DUP 33
SRR1766457.2827369 chrX 532814 N chrX 532984 N DUP 23
SRR1766481.10632956 chrX 532846 N chrX 533001 N DUP 32
SRR1766477.11106464 chrX 532814 N chrX 532987 N DUP 25
SRR1766462.4664999 chrX 532814 N chrX 532987 N DUP 25
SRR1766443.5911404 chrX 532814 N chrX 532987 N DUP 25
SRR1766447.4543671 chrX 532334 N chrX 533004 N DUP 20
SRR1766451.4329360 chrX 532334 N chrX 533004 N DUP 20
SRR1766442.35315888 chr13 27998968 N chr13 27999019 N DUP 24
SRR1766475.4958283 chr13 27998968 N chr13 27999019 N DUP 25
SRR1766484.9177243 chr13 27998968 N chr13 27999019 N DUP 27
SRR1766449.7027146 chr13 27998968 N chr13 27999019 N DUP 28
SRR1766472.11307815 chr13 27998968 N chr13 27999019 N DUP 30
SRR1766463.6908159 chr13 27998968 N chr13 27999019 N DUP 30
SRR1766483.6258830 chr13 27998983 N chr13 27999041 N DEL 21
SRR1766442.29273071 chr13 27998968 N chr13 27999019 N DUP 22
SRR1766447.5182355 chr13 27998962 N chr13 27999066 N DUP 28
SRR1766477.5162579 chr13 27998968 N chr13 27999019 N DUP 26
SRR1766448.3961823 chr13 27998968 N chr13 27999019 N DUP 27
SRR1766481.1593684 chr13 27998968 N chr13 27999019 N DUP 30
SRR1766463.10567222 chr13 27999013 N chr13 27999149 N DUP 26
SRR1766473.3699132 chr13 27999047 N chr13 27999112 N DUP 22
SRR1766452.7910045 chr13 27998967 N chr13 27999171 N DUP 23
SRR1766453.3680967 chr13 27998950 N chr13 27999150 N DUP 27
SRR1766470.6193709 chr13 27999305 N chr13 27999364 N DUP 27
SRR1766449.7959744 chr13 27999291 N chr13 27999368 N DEL 20
SRR1766477.4812811 chr8 141107639 N chr8 141107774 N DUP 23
SRR1766475.9833552 chr2 41747401 N chr2 41747610 N DUP 26
SRR1766460.651924 chr14 103896736 N chr14 103896870 N DEL 32
SRR1766462.8889482 chr14 103896737 N chr14 103896902 N DUP 27
SRR1766464.7045650 chr17 32027469 N chr17 32027546 N DEL 33
SRR1766480.4291630 chr10 127017132 N chr10 127017347 N DEL 27
SRR1766485.7632539 chrX 532905 N chrX 533078 N DUP 20
SRR1766477.11445418 chrX 532846 N chrX 533001 N DUP 33
SRR1766481.7843412 chrX 532846 N chrX 533001 N DUP 33
SRR1766457.2827369 chrX 532832 N chrX 533002 N DUP 23
SRR1766481.10632956 chrX 532846 N chrX 533001 N DUP 32
SRR1766477.11106464 chrX 532832 N chrX 533005 N DUP 25
SRR1766462.4664999 chrX 532832 N chrX 533005 N DUP 25
SRR1766443.5911404 chrX 532832 N chrX 533005 N DUP 25
SRR1766462.1476549 chr10 132335460 N chr10 132335657 N DEL 26
SRR1766450.607182 chr10 132335582 N chr10 132335782 N DEL 20
SRR1766443.3564480 chr1 193588279 N chr1 193588366 N DUP 20
SRR1766453.1152432 chr1 193588279 N chr1 193588366 N DUP 25
SRR1766470.610446 chr1 193588279 N chr1 193588366 N DUP 20
SRR1766444.1016580 chr19 32954938 N chr19 32955259 N DEL 24
SRR1766452.7683969 chr22 32565007 N chr22 32565128 N DEL 22
SRR1766470.9687831 chr8 144513945 N chr8 144514004 N DUP 24
SRR1766468.4218410 chr20 61173396 N chr20 61173575 N DEL 20
SRR1766481.10486062 chr2 108765460 N chr2 108765989 N DEL 24
SRR1766445.2550083 chr4 9981210 N chr4 9981460 N DEL 20
SRR1766444.130694 chr3 126008563 N chr3 126008665 N DEL 23
SRR1766462.37377 chr5 125632894 N chr5 125633008 N DUP 21
SRR1766445.1525882 chr5 125632894 N chr5 125633007 N DUP 20
SRR1766486.4586852 chr9 37918523 N chr9 37918584 N DEL 26
SRR1766484.288518 chr9 37918523 N chr9 37918584 N DEL 26
SRR1766475.5294056 chr19 39153429 N chr19 39153611 N DUP 20
SRR1766442.35551343 chr19 39153429 N chr19 39153611 N DUP 34
SRR1766452.5236743 chr19 39153429 N chr19 39153611 N DUP 36
SRR1766468.2261208 chr12 86502818 N chr12 86502946 N DEL 25
SRR1766442.31006958 chr5 1422521 N chr5 1422598 N DEL 20
SRR1766452.3373823 chr5 1423394 N chr5 1423531 N DUP 22
SRR1766444.2682053 chr5 1423121 N chr5 1423394 N DEL 26
SRR1766463.7541807 chr5 1422640 N chr5 1423199 N DEL 23
SRR1766448.5245341 chr5 1422628 N chr5 1423225 N DEL 25
SRR1766455.8397902 chr5 1422971 N chr5 1423356 N DEL 20
SRR1766452.3551185 chr5 1423356 N chr5 1423419 N DUP 26
SRR1766442.32985031 chr7 79625404 N chr7 79625731 N DEL 20
SRR1766448.4254032 chr7 79625404 N chr7 79625731 N DEL 20
SRR1766442.8894332 chr7 79625289 N chr7 79625731 N DEL 20
SRR1766473.10770663 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766452.1963307 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766482.608962 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766485.7101525 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766475.5230133 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766444.1004140 chr9 65463999 N chr9 65464292 N DEL 20
SRR1766454.4028571 chr19 40377443 N chr19 40377511 N DUP 30
SRR1766442.6322403 chr12 130843991 N chr12 130844094 N DEL 34
SRR1766442.7020145 chr18 72700585 N chr18 72700676 N DUP 21
SRR1766442.30657527 chr18 72700585 N chr18 72700676 N DUP 25
SRR1766448.3275279 chr18 72700585 N chr18 72700676 N DUP 25
SRR1766470.8099070 chr18 72700585 N chr18 72700676 N DUP 25
SRR1766447.1740189 chr18 72700585 N chr18 72700676 N DUP 33
SRR1766486.8736913 chr18 72700713 N chr18 72700768 N DUP 21
SRR1766446.5312837 chr18 72700723 N chr18 72700802 N DUP 20
SRR1766471.9090486 chr18 72700723 N chr18 72700802 N DUP 20
SRR1766473.4480261 chr18 72700713 N chr18 72700768 N DUP 24
SRR1766475.5339645 chr18 72700649 N chr18 72700824 N DUP 27
SRR1766454.10850453 chr18 72700798 N chr18 72700851 N DEL 20
SRR1766442.1681150 chr18 72700798 N chr18 72700851 N DEL 24
SRR1766474.8554568 chr18 72700798 N chr18 72700851 N DEL 24
SRR1766483.12153215 chr18 72700798 N chr18 72700851 N DEL 22
SRR1766477.7121867 chr18 72700798 N chr18 72700851 N DEL 21
SRR1766443.10371014 chr18 72700788 N chr18 72700851 N DEL 24
SRR1766477.10723407 chr18 72700788 N chr18 72700851 N DEL 23
SRR1766476.4863783 chr18 72700788 N chr18 72700851 N DEL 24
SRR1766467.4006965 chr18 72700799 N chr18 72700852 N DEL 21
SRR1766486.2793190 chr18 72700794 N chr18 72700857 N DEL 24
SRR1766448.9225421 chr18 72700672 N chr18 72700851 N DEL 20
SRR1766473.585183 chr18 72700727 N chr18 72700856 N DEL 22
SRR1766460.9078900 chr18 72700752 N chr18 72700851 N DEL 22
SRR1766465.1660947 chr18 72700752 N chr18 72700851 N DEL 21
SRR1766444.5777634 chr2 219217455 N chr2 219217749 N DEL 24
SRR1766444.937925 chr13 112913168 N chr13 112913367 N DEL 26
SRR1766452.5371918 chr1 4332502 N chr1 4332590 N DEL 20
SRR1766442.25037148 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766480.789992 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766469.1790376 chr1 4332556 N chr1 4332992 N DEL 22
SRR1766471.256383 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766443.3753855 chr1 4332556 N chr1 4333518 N DEL 20
SRR1766471.8142180 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766450.6375570 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766455.6174278 chr1 4332671 N chr1 4333223 N DEL 20
SRR1766460.9406510 chr1 4332556 N chr1 4332963 N DEL 20
SRR1766453.704886 chr5 2082196 N chr5 2082951 N DUP 20
SRR1766449.2189563 chr5 2082209 N chr5 2082964 N DUP 34
SRR1766459.10980685 chr5 2082196 N chr5 2082447 N DUP 20
SRR1766484.1156189 chr5 2082209 N chr5 2082964 N DUP 20
SRR1766478.1860006 chr5 2082209 N chr5 2082964 N DUP 30
SRR1766450.2008726 chr5 2082209 N chr5 2082964 N DUP 30
SRR1766443.610151 chr5 2082209 N chr5 2082964 N DUP 22
SRR1766485.7238556 chr5 2082906 N chr5 2082968 N DUP 21
SRR1766459.10336075 chr4 38880239 N chr4 38880295 N DEL 20
SRR1766449.5204186 chr16 22939935 N chr16 22940395 N DEL 25
SRR1766460.2025712 chr14 85847842 N chr14 85848173 N DEL 26
SRR1766467.11107955 chr14 85847842 N chr14 85848173 N DEL 26
SRR1766482.7098379 chr14 85847842 N chr14 85848173 N DEL 20
SRR1766477.3232805 chr14 85847948 N chr14 85848239 N DEL 20
SRR1766448.9952925 chr17 83172689 N chr17 83173481 N DEL 28
SRR1766463.7038479 chr17 83172689 N chr17 83173367 N DEL 20
SRR1766446.2336436 chr10 46136103 N chr10 46136168 N DEL 21
SRR1766465.8064377 chr13 18944529 N chr13 18945170 N DEL 20
SRR1766482.1963407 chr5 175050953 N chr5 175051008 N DUP 25
SRR1766449.1821551 chr5 175050953 N chr5 175051008 N DUP 36
SRR1766482.12957866 chr5 175050969 N chr5 175051024 N DUP 27
SRR1766455.3355411 chr5 175050969 N chr5 175051024 N DUP 27
SRR1766442.39217338 chr5 175050953 N chr5 175051008 N DUP 37
SRR1766461.5058047 chr5 175050953 N chr5 175051008 N DUP 37
SRR1766475.3288234 chr5 175050955 N chr5 175051037 N DUP 26
SRR1766454.8584461 chr5 175050955 N chr5 175051037 N DUP 28
SRR1766467.11469131 chr5 175050955 N chr5 175051037 N DUP 24
SRR1766459.7085575 chr5 175050955 N chr5 175051037 N DUP 30
SRR1766458.4133442 chr5 175050945 N chr5 175051029 N DUP 34
SRR1766447.4007054 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766447.9114426 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766448.4957899 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766448.7792711 chr5 175050955 N chr5 175051037 N DUP 39
SRR1766452.10321710 chr5 175050945 N chr5 175051029 N DUP 38
SRR1766455.6790559 chr5 175050953 N chr5 175051008 N DUP 31
SRR1766472.4827124 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766479.9037325 chr5 175050945 N chr5 175051029 N DUP 38
SRR1766481.11873666 chr5 175050945 N chr5 175051029 N DUP 36
SRR1766447.4007054 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766451.1959023 chr5 175050945 N chr5 175051029 N DUP 38
SRR1766454.6574963 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766456.4092508 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766457.8785463 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766470.7788759 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766472.2327221 chr5 175050955 N chr5 175051037 N DUP 38
SRR1766447.413892 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766452.6976528 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766457.4840642 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766470.7313587 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766478.6602309 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766484.10286372 chr5 175050944 N chr5 175051028 N DUP 33
SRR1766442.35734643 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766450.5203004 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766461.5058047 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766455.1892458 chr5 175050945 N chr5 175051029 N DUP 34
SRR1766472.39408 chr5 175050945 N chr5 175051029 N DUP 34
SRR1766480.8347342 chr5 175050945 N chr5 175051029 N DUP 34
SRR1766461.7579894 chr5 175050953 N chr5 175051008 N DUP 25
SRR1766451.8483047 chr5 175050944 N chr5 175051028 N DUP 34
SRR1766447.9114426 chr5 175050953 N chr5 175051008 N DUP 24
SRR1766462.9281737 chr5 175050953 N chr5 175051008 N DUP 24
SRR1766467.2137023 chr5 175050953 N chr5 175051008 N DUP 30
SRR1766469.8261633 chr5 175050944 N chr5 175051028 N DUP 34
SRR1766474.9737249 chr5 175050944 N chr5 175051028 N DUP 29
SRR1766468.7190526 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766475.10314943 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766453.5373669 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766468.82812 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766450.6205861 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.8470335 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766470.4308219 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.46260196 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.17570005 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766453.9692498 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.11277883 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766463.7644666 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.43724364 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766446.2875471 chr14 48710753 N chr14 48710986 N DUP 22
SRR1766450.2967389 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766472.10603905 chr14 48710753 N chr14 48710986 N DUP 23
SRR1766462.2861715 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766465.9454850 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766443.6859543 chr14 48710753 N chr14 48710986 N DUP 20
SRR1766446.7779737 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766483.3811038 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766457.5768050 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766467.3768663 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766448.2507356 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766442.31012994 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766463.5102635 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766470.5233128 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766483.7327647 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766453.10379217 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766445.3167664 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766460.6129341 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766474.1487035 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766485.2389651 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766468.5267218 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766479.2762163 chr14 48710814 N chr14 48710959 N DEL 25
SRR1766452.9985132 chr4 48104421 N chr4 48104514 N DEL 21
SRR1766451.311775 chr4 48104421 N chr4 48104514 N DEL 22
SRR1766442.15647221 chr4 48104420 N chr4 48104625 N DEL 23
SRR1766442.32996336 chr4 48104464 N chr4 48104691 N DEL 21
SRR1766476.10020416 chr4 48104420 N chr4 48104625 N DEL 24
SRR1766486.5629839 chr4 48104464 N chr4 48104691 N DEL 24
SRR1766454.1951430 chr4 48104420 N chr4 48104625 N DEL 27
SRR1766451.821205 chr4 48104420 N chr4 48104625 N DEL 28
SRR1766477.5593298 chr4 48104464 N chr4 48104691 N DEL 27
SRR1766453.3320851 chr4 48104464 N chr4 48104691 N DEL 27
SRR1766459.2554158 chr4 48104420 N chr4 48104625 N DEL 27
SRR1766481.10027804 chr4 48104420 N chr4 48104625 N DEL 26
SRR1766442.26239820 chr4 48104464 N chr4 48104691 N DEL 33
SRR1766442.36144754 chr4 48104464 N chr4 48104691 N DEL 33
SRR1766456.1433357 chr4 48104417 N chr4 48104684 N DEL 28
SRR1766456.955390 chr4 48104682 N chr4 48104739 N DUP 20
SRR1766442.496214 chr11 86732407 N chr11 86732741 N DUP 20
SRR1766477.9656294 chr2 57548108 N chr2 57548161 N DEL 29
SRR1766442.19056028 chr2 57548108 N chr2 57548161 N DEL 27
SRR1766470.6887218 chr2 57548108 N chr2 57548161 N DEL 24
SRR1766462.10334310 chrX 136451220 N chrX 136451269 N DUP 21
SRR1766451.5315885 chr5 180297012 N chr5 180297105 N DEL 24
SRR1766472.5620055 chr5 180297012 N chr5 180297105 N DEL 23
SRR1766462.7149598 chr16 7229912 N chr16 7230179 N DUP 25
SRR1766452.2071920 chr16 7229912 N chr16 7230179 N DUP 25
SRR1766453.10549147 chr16 7230002 N chr16 7230179 N DUP 20
SRR1766442.1922502 chr14 89567556 N chr14 89567720 N DUP 27
SRR1766473.6022383 chr14 89567556 N chr14 89567654 N DUP 27
SRR1766460.9566402 chr14 89567589 N chr14 89567654 N DUP 30
SRR1766449.3225221 chr14 89567589 N chr14 89567654 N DUP 30
SRR1766449.4399257 chr14 89567556 N chr14 89567654 N DUP 25
SRR1766454.6520794 chr14 89567556 N chr14 89567654 N DUP 25
SRR1766458.3737403 chr14 89567556 N chr14 89567654 N DUP 25
SRR1766442.43692910 chr14 89567621 N chr14 89567688 N DEL 30
SRR1766475.9134706 chr14 86443422 N chr14 86443494 N DEL 20
SRR1766465.9250892 chr14 86443422 N chr14 86443494 N DEL 25
SRR1766460.8005540 chr14 86443460 N chr14 86443513 N DUP 24
SRR1766466.10372861 chr14 86443460 N chr14 86443513 N DUP 27
SRR1766472.8052251 chr14 86443460 N chr14 86443552 N DUP 37
SRR1766442.7367609 chr14 86443460 N chr14 86443513 N DUP 33
SRR1766442.28998354 chr14 86443476 N chr14 86443573 N DUP 32
SRR1766486.5411664 chr14 86443460 N chr14 86443513 N DUP 34
SRR1766481.12920665 chr14 86443460 N chr14 86443513 N DUP 35
SRR1766448.2943442 chr14 86443460 N chr14 86443584 N DUP 36
SRR1766452.6550543 chr14 86443478 N chr14 86443548 N DUP 31
SRR1766470.5723466 chr14 86443460 N chr14 86443584 N DUP 36
SRR1766463.6288637 chr14 86443460 N chr14 86443584 N DUP 35
SRR1766475.4870310 chr14 86443478 N chr14 86443548 N DUP 30
SRR1766442.34630070 chr14 86443460 N chr14 86443513 N DUP 26
SRR1766461.11011897 chr14 86443478 N chr14 86443548 N DUP 30
SRR1766470.611993 chr14 86443478 N chr14 86443548 N DUP 33
SRR1766442.7954196 chr14 86443478 N chr14 86443548 N DUP 34
SRR1766459.6923307 chr14 86443478 N chr14 86443548 N DUP 28
SRR1766467.7149342 chr14 86443460 N chr14 86443513 N DUP 23
SRR1766460.2752859 chr14 86443478 N chr14 86443548 N DUP 24
SRR1766464.2892468 chr14 86443478 N chr14 86443548 N DUP 25
SRR1766454.1807925 chr14 86443635 N chr14 86443737 N DEL 29
SRR1766462.2928365 chr14 86443577 N chr14 86443685 N DEL 22
SRR1766461.3674012 chr14 86443635 N chr14 86443737 N DEL 34
SRR1766483.3498350 chr14 86443635 N chr14 86443737 N DEL 34
SRR1766486.3612478 chr14 86443635 N chr14 86443737 N DEL 34
SRR1766463.349530 chr14 86443635 N chr14 86443737 N DEL 20
SRR1766448.10153681 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766471.4194 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766449.8655581 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766454.4271292 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766482.7644767 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766473.751926 chr14 86443763 N chr14 86443844 N DUP 24
SRR1766476.939331 chr14 86444059 N chr14 86444112 N DEL 20
SRR1766470.2305340 chr14 86444059 N chr14 86444112 N DEL 23
SRR1766464.4151464 chr14 86444059 N chr14 86444112 N DEL 27
SRR1766442.7259017 chr14 86444059 N chr14 86444112 N DEL 33
SRR1766442.30329864 chr14 86444059 N chr14 86444112 N DEL 36
SRR1766452.6844358 chr14 86443884 N chr14 86444112 N DEL 23
SRR1766447.6390002 chr14 86443884 N chr14 86444112 N DEL 23
SRR1766461.3674012 chr14 86443884 N chr14 86444112 N DEL 23
SRR1766461.1350871 chr12 127166359 N chr12 127166438 N DUP 35
SRR1766482.4679794 chr12 127166345 N chr12 127166404 N DUP 29
SRR1766454.8431121 chr12 127166359 N chr12 127166438 N DUP 32
SRR1766464.783149 chr12 127166359 N chr12 127166438 N DUP 33
SRR1766472.51397 chr12 127166359 N chr12 127166468 N DUP 31
SRR1766479.12580237 chr3 93470409 N chr3 93470458 N DUP 37
SRR1766483.573341 chr3 93470409 N chr3 93470458 N DUP 38
SRR1766478.228532 chr3 93470409 N chr3 93470458 N DUP 38
SRR1766442.33326029 chr3 93470408 N chr3 93470457 N DUP 32
SRR1766448.8458862 chr3 93470409 N chr3 93470458 N DUP 30
SRR1766449.8704930 chr3 93470409 N chr3 93470458 N DUP 27
SRR1766450.6321970 chr3 93470409 N chr3 93470458 N DUP 39
SRR1766479.2916449 chr4 163894706 N chr4 163894774 N DUP 27
SRR1766482.8152960 chr4 163894706 N chr4 163894774 N DUP 27
SRR1766447.11446666 chr4 163894706 N chr4 163894774 N DUP 28
SRR1766471.5449216 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766478.1121405 chr4 163894706 N chr4 163894774 N DUP 34
SRR1766442.13216659 chr4 163894706 N chr4 163894774 N DUP 28
SRR1766442.23537322 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766459.9368097 chr4 163894706 N chr4 163894774 N DUP 34
SRR1766460.10824500 chr4 163894706 N chr4 163894774 N DUP 31
SRR1766467.6722339 chr4 163894706 N chr4 163894774 N DUP 30
SRR1766471.1311902 chr4 163894706 N chr4 163894774 N DUP 34
SRR1766471.6440397 chr4 163894706 N chr4 163894774 N DUP 33
SRR1766472.9948279 chr4 163894706 N chr4 163894774 N DUP 31
SRR1766479.8815481 chr4 163894706 N chr4 163894774 N DUP 34
SRR1766442.10322986 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766442.12261298 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766443.6385912 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766449.6458596 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766472.2736243 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766449.6186756 chr4 163894706 N chr4 163894774 N DUP 27
SRR1766446.3686635 chr4 163894706 N chr4 163894774 N DUP 27
SRR1766447.771987 chr4 163894706 N chr4 163894774 N DUP 28
SRR1766446.2422617 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766471.1652729 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766477.9359985 chr4 163894706 N chr4 163894774 N DUP 30
SRR1766469.4720168 chr4 163894706 N chr4 163894774 N DUP 32
SRR1766469.6241735 chr4 163894706 N chr4 163894774 N DUP 32
SRR1766466.9190665 chr4 163894780 N chr4 163894840 N DEL 22
SRR1766457.4566415 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766468.5657479 chr4 163894780 N chr4 163894840 N DEL 27
SRR1766470.5628948 chr4 163894757 N chr4 163894840 N DEL 25
SRR1766463.1287744 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766464.10859506 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766469.5846318 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766455.3996277 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766442.2394403 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766469.5548198 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766484.11020182 chrX 57698188 N chrX 57698702 N DUP 27
SRR1766463.1756856 chrX 57698191 N chrX 57698743 N DUP 22
SRR1766442.22382523 chrX 57698352 N chrX 57698793 N DEL 20
SRR1766445.8343522 chr2 131754041 N chr2 131755478 N DUP 20
SRR1766461.803893 chr9 128439918 N chr9 128440214 N DEL 20
SRR1766442.15552778 chr19 34534847 N chr19 34534916 N DUP 21
SRR1766470.5214552 chr19 34534869 N chr19 34534942 N DUP 31
SRR1766472.2362149 chr19 34534867 N chr19 34534928 N DUP 32
SRR1766455.9153626 chr3 159680839 N chr3 159680899 N DUP 21
SRR1766476.7357564 chr3 159680839 N chr3 159680899 N DUP 21
SRR1766448.10566826 chr11 112324043 N chr11 112325032 N DEL 29
SRR1766473.523687 chrX 72179191 N chrX 72179359 N DEL 20
SRR1766485.6598329 chr3 143449252 N chr3 143449760 N DEL 28
SRR1766452.939341 chr3 143449536 N chr3 143449697 N DUP 26
SRR1766486.2874702 chr3 143449617 N chr3 143449670 N DEL 22
SRR1766479.8359576 chr3 143449794 N chr3 143449872 N DUP 34
SRR1766479.5543580 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766481.7765743 chr3 143449760 N chr3 143449866 N DUP 33
SRR1766484.691538 chr3 143449201 N chr3 143449794 N DEL 22
SRR1766472.441327 chr3 143449763 N chr3 143449874 N DUP 23
SRR1766447.9621093 chr3 143449763 N chr3 143449874 N DUP 23
SRR1766477.4764861 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766462.3480851 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766465.11120355 chr3 143449763 N chr3 143449846 N DUP 22
SRR1766475.2600938 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766484.2298927 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766460.1120946 chr3 143449806 N chr3 143449860 N DUP 24
SRR1766465.928632 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766442.22868292 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766446.3454657 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766482.12637828 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766449.8666212 chr18 54780375 N chr18 54780531 N DEL 32
SRR1766453.4893866 chr18 54780375 N chr18 54780531 N DEL 32
SRR1766469.10985631 chr18 54780375 N chr18 54780531 N DEL 32
SRR1766460.4061683 chr18 54780375 N chr18 54780531 N DEL 25
SRR1766471.5538539 chr6 169957126 N chr6 169957298 N DEL 32
SRR1766485.9785545 chr6 169957309 N chr6 169957483 N DEL 22
SRR1766454.3516641 chr7 100995098 N chr7 100995846 N DEL 20
SRR1766479.7732507 chr7 100994654 N chr7 100995408 N DEL 25
SRR1766442.26434261 chr10 126947600 N chr10 126947697 N DEL 21
SRR1766461.6115088 chr10 126947489 N chr10 126948593 N DEL 22
SRR1766475.5677341 chr10 52834289 N chr10 52834484 N DEL 23
SRR1766468.3609739 chr10 52834246 N chr10 52834302 N DUP 25
SRR1766473.1894817 chr10 52834617 N chr10 52834964 N DEL 26
SRR1766471.3025623 chr10 52834265 N chr10 52834466 N DUP 27
SRR1766465.4275800 chr10 52834306 N chr10 52834544 N DEL 22
SRR1766484.4009 chr10 52835393 N chr10 52835520 N DUP 23
SRR1766468.5156569 chr10 52834486 N chr10 52834698 N DUP 21
SRR1766467.824677 chr10 52834481 N chr10 52834553 N DUP 24
SRR1766470.10552302 chr10 52834192 N chr10 52834339 N DUP 21
SRR1766486.4689209 chr10 52834961 N chr10 52835471 N DUP 27
SRR1766466.10643060 chr10 52834584 N chr10 52834705 N DEL 27
SRR1766477.6829744 chr10 52834231 N chr10 52834896 N DEL 24
SRR1766457.538449 chr10 52834215 N chr10 52834348 N DEL 22
SRR1766483.4245322 chr10 52834329 N chr10 52834501 N DEL 22
SRR1766473.4486536 chr10 52834377 N chr10 52834998 N DUP 20
SRR1766471.11790596 chr10 52834246 N chr10 52834302 N DUP 25
SRR1766476.7922702 chr10 52834262 N chr10 52834452 N DUP 24
SRR1766484.12078672 chr10 52834348 N chr10 52834996 N DUP 21
SRR1766450.7046305 chr10 52834882 N chr10 52835011 N DUP 25
SRR1766452.5302509 chr10 52834377 N chr10 52834998 N DUP 20
SRR1766460.7474422 chr10 52834265 N chr10 52834466 N DUP 22
SRR1766472.2495678 chr10 52835012 N chr10 52835442 N DEL 20
SRR1766476.10022101 chr10 52834262 N chr10 52834452 N DUP 23
SRR1766475.11081218 chr10 52834282 N chr10 52834479 N DEL 23
SRR1766485.2973743 chr10 52834212 N chr10 52834357 N DEL 25
SRR1766471.430497 chr10 52834845 N chr10 52834903 N DEL 24
SRR1766465.887054 chr10 52834584 N chr10 52834705 N DEL 27
SRR1766478.6423002 chr10 52834265 N chr10 52834466 N DUP 22
SRR1766447.7849046 chr10 52834348 N chr10 52834996 N DUP 22
SRR1766467.9335405 chr10 52834963 N chr10 52835230 N DUP 23
SRR1766461.4203167 chr10 52834888 N chr10 52834982 N DUP 23
SRR1766452.7871041 chr10 52834592 N chr10 52834953 N DUP 22
SRR1766447.9225541 chr10 52834348 N chr10 52834444 N DUP 20
SRR1766442.28290693 chr10 52834974 N chr10 52835037 N DUP 20
SRR1766443.2792696 chr10 52834212 N chr10 52834357 N DEL 24
SRR1766464.6711284 chr10 52834300 N chr10 52834541 N DEL 20
SRR1766468.4012834 chr10 52834584 N chr10 52834705 N DEL 22
SRR1766456.1725809 chr10 52834966 N chr10 52835029 N DUP 29
SRR1766446.2319339 chr10 52834845 N chr10 52834903 N DEL 23
SRR1766483.2483593 chr10 52834171 N chr10 52834689 N DUP 29
SRR1766461.2464575 chr10 52834192 N chr10 52834318 N DUP 26
SRR1766484.3548182 chr10 52834592 N chr10 52834953 N DUP 22
SRR1766453.2168285 chr10 52834882 N chr10 52835011 N DUP 27
SRR1766461.8160401 chr18 1747179 N chr18 1747240 N DUP 20
SRR1766459.5551605 chr5 38832251 N chr5 38832338 N DEL 20
SRR1766452.9628770 chr17 83120204 N chr17 83120258 N DEL 25
SRR1766449.3155568 chr3 50076518 N chr3 50076824 N DEL 26
SRR1766480.2808339 chr10 6413623 N chr10 6413738 N DEL 22
SRR1766481.6314684 chr10 6413628 N chr10 6413686 N DUP 21
SRR1766471.10342797 chr10 6413627 N chr10 6413787 N DEL 33
SRR1766485.5284021 chr10 6413627 N chr10 6413787 N DEL 35
SRR1766486.2323722 chr10 6413700 N chr10 6413787 N DEL 30
SRR1766445.9976419 chr3 195710745 N chr3 195710881 N DEL 23
SRR1766442.30048324 chr3 195710777 N chr3 195711138 N DEL 20
SRR1766442.19902109 chr3 195710637 N chr3 195711221 N DUP 20
SRR1766474.9856445 chr3 195711182 N chr3 195711453 N DEL 22
SRR1766453.2806591 chr3 195710745 N chr3 195710836 N DEL 20
SRR1766460.5415474 chr3 195710745 N chr3 195710836 N DEL 25
SRR1766460.1511398 chr3 195710789 N chr3 195711373 N DUP 20
SRR1766453.5877578 chr3 195710573 N chr3 195710799 N DEL 23
SRR1766454.10630146 chr3 195710778 N chr3 195711409 N DEL 21
SRR1766477.1346454 chr3 195710700 N chr3 195710836 N DEL 20
SRR1766479.12792430 chr3 195710781 N chr3 195711578 N DEL 25
SRR1766464.8428911 chr3 195710745 N chr3 195710836 N DEL 23
SRR1766449.2039271 chr3 195710833 N chr3 195710922 N DUP 20
SRR1766459.6172648 chr3 195710656 N chr3 195710745 N DUP 20
SRR1766466.2910937 chr3 195710788 N chr3 195710879 N DEL 20
SRR1766445.5415585 chr3 195711047 N chr3 195711574 N DEL 25
SRR1766447.11284297 chr3 195710574 N chr3 195710888 N DUP 25
SRR1766451.7640748 chr3 195710745 N chr3 195711286 N DEL 20
SRR1766451.7364049 chr3 195710833 N chr3 195710967 N DUP 23
SRR1766446.3317050 chr3 195711089 N chr3 195711405 N DEL 26
SRR1766482.8002010 chr3 195710777 N chr3 195711138 N DEL 21
SRR1766457.8733614 chr3 195710878 N chr3 195711372 N DUP 20
SRR1766479.9603242 chr3 195710925 N chr3 195711151 N DEL 20
SRR1766466.2795537 chr3 195711047 N chr3 195711574 N DEL 28
SRR1766471.4813397 chr3 195710789 N chr3 195711373 N DUP 22
SRR1766467.9044595 chr3 195710788 N chr3 195710879 N DEL 20
SRR1766471.10686592 chr3 195710472 N chr3 195710833 N DEL 20
SRR1766454.63412 chr3 195710788 N chr3 195710879 N DEL 20
SRR1766464.416862 chr3 195710833 N chr3 195710922 N DUP 20
SRR1766450.9241373 chr3 195710818 N chr3 195711613 N DUP 20
SRR1766456.2591922 chr7 1384768 N chr7 1384842 N DEL 28
SRR1766453.6868035 chr8 138805065 N chr8 138806007 N DEL 30
SRR1766477.2720172 chr8 138806218 N chr8 138806279 N DEL 21
SRR1766483.5259067 chr8 138806218 N chr8 138806279 N DEL 24
SRR1766453.10004252 chr8 138806218 N chr8 138806279 N DEL 24
SRR1766473.1844425 chr19 14314279 N chr19 14314430 N DEL 20
SRR1766481.2524873 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766442.42263299 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766448.11007892 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766463.9881219 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766462.4506747 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766453.2777982 chr21 30210371 N chr21 30210421 N DUP 21
SRR1766478.9624827 chr21 30210371 N chr21 30210421 N DUP 25
SRR1766477.5047197 chr1 152910459 N chr1 152910910 N DEL 35
SRR1766484.7504615 chr1 152910444 N chr1 152910715 N DEL 20
SRR1766442.1937426 chr1 152910562 N chr1 152910713 N DEL 20
SRR1766464.2543136 chr1 152910530 N chr1 152910801 N DEL 20
SRR1766448.115485 chr1 152910590 N chr1 152911011 N DEL 29
SRR1766448.5359956 chr1 152910573 N chr1 152911375 N DEL 38
SRR1766468.7180568 chr1 152910873 N chr1 152911375 N DEL 22
SRR1766475.10239803 chr8 53948571 N chr8 53949132 N DEL 20
SRR1766448.3359006 chr8 53949358 N chr8 53949423 N DUP 23
SRR1766444.7125359 chr8 53949351 N chr8 53949416 N DUP 22
SRR1766460.6027258 chr8 53949349 N chr8 53949414 N DUP 20
SRR1766473.1960105 chr8 53949349 N chr8 53949414 N DUP 26
SRR1766442.4347839 chr8 53949349 N chr8 53949414 N DUP 25
SRR1766481.1865092 chr8 53949349 N chr8 53949414 N DUP 25
SRR1766461.10896229 chr8 53949349 N chr8 53949414 N DUP 21
SRR1766451.3608378 chr8 53949349 N chr8 53949414 N DUP 22
SRR1766474.3445500 chr8 53949349 N chr8 53949414 N DUP 23
SRR1766485.9463329 chr8 53949349 N chr8 53949414 N DUP 22
SRR1766460.441049 chr8 53949349 N chr8 53949414 N DUP 21
SRR1766477.635213 chr8 53949349 N chr8 53949414 N DUP 22
SRR1766486.8335902 chr8 53949349 N chr8 53949414 N DUP 22
SRR1766448.4220291 chr8 53949349 N chr8 53949414 N DUP 24
SRR1766463.2129608 chr8 53949349 N chr8 53949414 N DUP 24
SRR1766469.8102695 chr8 53949349 N chr8 53949414 N DUP 24
SRR1766453.2819308 chr8 53949349 N chr8 53949414 N DUP 25
SRR1766486.3462545 chr1 193564094 N chr1 193564157 N DUP 20
SRR1766471.8347138 chr1 193564152 N chr1 193564215 N DUP 24
SRR1766476.3882521 chr1 193564152 N chr1 193564215 N DUP 21
SRR1766479.11486539 chr4 47123656 N chr4 47123728 N DEL 32
SRR1766468.7902720 chr4 47123656 N chr4 47123728 N DEL 28
SRR1766469.668495 chr4 47123656 N chr4 47123728 N DEL 29
SRR1766476.461666 chr7 98548123 N chr7 98548208 N DEL 20
SRR1766461.8064668 chr7 98548235 N chr7 98548690 N DUP 21
SRR1766458.1981564 chr7 98548225 N chr7 98548276 N DUP 22
SRR1766484.11219731 chr7 98548225 N chr7 98548276 N DUP 28
SRR1766462.1249024 chr7 98548200 N chr7 98548307 N DUP 22
SRR1766448.2205439 chr7 98548218 N chr7 98548525 N DUP 22
SRR1766475.3967999 chr7 98548245 N chr7 98548466 N DEL 26
SRR1766452.3016551 chr7 98548186 N chr7 98548645 N DUP 31
SRR1766442.7191805 chr7 98548235 N chr7 98548690 N DUP 29
SRR1766466.2797376 chr19 51944903 N chr19 51945156 N DEL 25
SRR1766485.9605830 chr6 59360896 N chr6 59361217 N DEL 20
SRR1766484.9393062 chr11 131265291 N chr11 131265465 N DEL 22
SRR1766442.22279736 chr11 131265291 N chr11 131265465 N DEL 24
SRR1766448.674019 chr11 131265291 N chr11 131265465 N DEL 24
SRR1766476.7224224 chr11 131265291 N chr11 131265465 N DEL 24
SRR1766485.10255151 chr11 131265325 N chr11 131265447 N DEL 30
SRR1766445.8661391 chr11 131265291 N chr11 131265465 N DEL 26
SRR1766458.1558429 chr11 131265291 N chr11 131265465 N DEL 26
SRR1766475.1156443 chr11 131265325 N chr11 131265447 N DEL 30
SRR1766448.6456425 chr11 131265325 N chr11 131265447 N DEL 30
SRR1766451.9100705 chr11 131265291 N chr11 131265465 N DEL 26
SRR1766485.9338154 chr11 131265291 N chr11 131265465 N DEL 26
SRR1766479.3546291 chr11 131265325 N chr11 131265447 N DEL 30
SRR1766467.219304 chr11 131265291 N chr11 131265465 N DEL 30
SRR1766451.4150346 chr11 131265352 N chr11 131265544 N DUP 21
SRR1766466.292360 chr8 142205166 N chr8 142205237 N DEL 22
SRR1766476.535031 chr4 43451137 N chr4 43451231 N DEL 34
SRR1766479.10388521 chr1 2960156 N chr1 2960277 N DEL 25
SRR1766442.26579387 chr6 4895507 N chr6 4895622 N DEL 21
SRR1766444.1029360 chr20 63871760 N chr20 63872045 N DEL 32
SRR1766470.2305551 chr1 143218205 N chr1 143218298 N DUP 22
SRR1766470.2298968 chr1 143218118 N chr1 143218283 N DUP 23
SRR1766452.746458 chr1 143218118 N chr1 143218283 N DUP 24
SRR1766467.9996857 chr6 169924033 N chr6 169924140 N DUP 28
SRR1766442.17343206 chr6 169924033 N chr6 169924254 N DUP 24
SRR1766468.3918415 chr6 169923954 N chr6 169924136 N DUP 20
SRR1766482.4613517 chr6 169923954 N chr6 169924136 N DUP 22
SRR1766467.2115205 chr6 169924004 N chr6 169924105 N DUP 24
SRR1766474.10375373 chr10 2392620 N chr10 2392783 N DUP 28
SRR1766447.460340 chr10 60240162 N chr10 60240282 N DUP 31
SRR1766457.6485003 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766461.10565373 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766451.8173222 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766443.2558803 chr10 60240271 N chr10 60240402 N DUP 20
SRR1766461.34003 chr21 8464792 N chr21 8464898 N DUP 21
SRR1766473.3235767 chr21 8464715 N chr21 8464897 N DUP 24
SRR1766451.6536886 chr21 8464792 N chr21 8464894 N DUP 20
SRR1766442.620304 chr21 8464833 N chr21 8464942 N DUP 21
SRR1766459.1611681 chr21 8464457 N chr21 8464830 N DEL 21
SRR1766446.6490081 chr21 8464792 N chr21 8464900 N DUP 25
SRR1766453.7794336 chr21 8464794 N chr21 8464902 N DUP 34
SRR1766486.3641391 chrX 107204870 N chrX 107205043 N DEL 21
SRR1766468.1757784 chrX 107204870 N chrX 107205043 N DEL 24
SRR1766462.2979910 chrX 107204870 N chrX 107205043 N DEL 26
SRR1766478.3051211 chrX 107204827 N chrX 107204882 N DUP 26
SRR1766442.9865723 chrX 107204827 N chrX 107204882 N DUP 26
SRR1766443.4347326 chrX 107204827 N chrX 107205110 N DUP 33
SRR1766454.3763868 chrX 107204827 N chrX 107205110 N DUP 30
SRR1766471.9933313 chrX 107204827 N chrX 107205110 N DUP 31
SRR1766486.1230929 chrX 107204847 N chrX 107204902 N DUP 26
SRR1766463.2942810 chrX 107204827 N chrX 107204882 N DUP 26
SRR1766473.3981399 chrX 107204922 N chrX 107205043 N DEL 20
SRR1766457.6266848 chrX 107204827 N chrX 107205110 N DUP 34
SRR1766466.4236866 chrX 107204898 N chrX 107205043 N DEL 27
SRR1766485.724969 chrX 107204898 N chrX 107205043 N DEL 27
SRR1766465.2348161 chrX 107204898 N chrX 107205043 N DEL 26
SRR1766447.6559092 chrX 107204898 N chrX 107205043 N DEL 26
SRR1766467.9269252 chrX 107204922 N chrX 107205043 N DEL 21
SRR1766454.4028571 chr19 40377443 N chr19 40377511 N DUP 30
SRR1766484.5433352 chr1 34102766 N chr1 34102824 N DEL 34
SRR1766453.3143994 chr1 34102766 N chr1 34102824 N DEL 30
SRR1766443.8046965 chr1 34102766 N chr1 34102824 N DEL 28
SRR1766475.5642958 chr1 34102722 N chr1 34102818 N DEL 20
SRR1766452.4723694 chr1 34102766 N chr1 34102824 N DEL 25
SRR1766478.3716221 chr1 34102766 N chr1 34102824 N DEL 25
SRR1766481.5713646 chr1 34102766 N chr1 34102824 N DEL 21
SRR1766486.9056919 chr5 1272674 N chr5 1273724 N DEL 25
SRR1766464.9101210 chr5 1272674 N chr5 1273724 N DEL 33
SRR1766476.8657152 chr5 1272674 N chr5 1273724 N DEL 28
SRR1766474.6306011 chr5 1272828 N chr5 1273738 N DEL 20
SRR1766462.1593480 chr5 1272950 N chr5 1273940 N DEL 33
SRR1766453.8101317 chr5 1272844 N chr5 1273940 N DEL 29
SRR1766460.8119854 chr5 1272950 N chr5 1273940 N DEL 36
SRR1766459.4436321 chr5 1272844 N chr5 1273940 N DEL 29
SRR1766483.2079340 chr5 1272950 N chr5 1273940 N DEL 36
SRR1766472.437435 chr5 1272950 N chr5 1273940 N DEL 36
SRR1766461.10590260 chr5 1272950 N chr5 1273940 N DEL 35
SRR1766452.1640759 chr5 1272844 N chr5 1273940 N DEL 24
SRR1766476.9508035 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766480.5186410 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766442.12661975 chr5 1272817 N chr5 1273951 N DEL 27
SRR1766442.43499975 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766468.5427890 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766480.8591848 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766460.8119854 chr5 1272772 N chr5 1273940 N DEL 27
SRR1766449.7348751 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766481.1203964 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766485.4631770 chr7 1295512 N chr7 1295592 N DEL 22
SRR1766482.9747560 chr3 198168406 N chr3 198168752 N DEL 23
SRR1766447.9259204 chr21 14261871 N chr21 14261948 N DUP 23
SRR1766442.33116854 chr21 45502086 N chr21 45502218 N DEL 22
SRR1766447.3396728 chr21 45502086 N chr21 45502218 N DEL 31
SRR1766456.4267116 chr21 45502086 N chr21 45502218 N DEL 30
SRR1766474.2654014 chr21 45502086 N chr21 45502218 N DEL 24
SRR1766454.6352513 chr21 45502086 N chr21 45502218 N DEL 23
SRR1766471.12028313 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766477.4370754 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766461.5320310 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766473.7606447 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766448.840955 chr21 45502108 N chr21 45502239 N DEL 38
SRR1766443.9979007 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766472.8823673 chr21 45502108 N chr21 45502239 N DEL 38
SRR1766452.863021 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766454.7710972 chr21 45502108 N chr21 45502239 N DEL 38
SRR1766469.4529495 chr21 45502108 N chr21 45502239 N DEL 22
SRR1766464.4951487 chr21 45502108 N chr21 45502239 N DEL 22
SRR1766448.9862027 chr21 45502108 N chr21 45502239 N DEL 22
SRR1766483.8762190 chr21 45502108 N chr21 45502239 N DEL 22
SRR1766485.3080118 chr19 621074 N chr19 621137 N DEL 22
SRR1766449.3144827 chr19 621074 N chr19 621137 N DEL 23
SRR1766458.1133797 chr19 621074 N chr19 621137 N DEL 26
SRR1766461.2564736 chr12 132317140 N chr12 132317242 N DUP 36
SRR1766448.9099191 chr6 1542134 N chr6 1542359 N DEL 36
SRR1766456.3063338 chr1 11522690 N chr1 11522911 N DEL 20
SRR1766471.4990592 chr1 11522701 N chr1 11522790 N DEL 25
SRR1766462.9815771 chr1 11522701 N chr1 11522834 N DEL 23
SRR1766459.6434565 chr1 11522701 N chr1 11522790 N DEL 37
SRR1766442.13372194 chr1 11522672 N chr1 11522981 N DEL 20
SRR1766482.3461498 chr1 11522745 N chr1 11522944 N DEL 21
SRR1766444.3020589 chr1 11522932 N chr1 11522997 N DUP 20
SRR1766459.11097738 chr1 11522789 N chr1 11522964 N DUP 26
SRR1766448.8745751 chr1 11522680 N chr1 11522976 N DUP 32
SRR1766442.36692428 chr1 11522778 N chr1 11523008 N DUP 20
SRR1766472.1438968 chr1 11522673 N chr1 11522914 N DUP 20
SRR1766481.3241932 chr1 11522878 N chr1 11523042 N DUP 25
SRR1766467.2534300 chr1 11522789 N chr1 11522887 N DUP 20
SRR1766458.598827 chr1 11522759 N chr1 11522958 N DEL 20
SRR1766468.1363934 chr1 11522833 N chr1 11522898 N DUP 25
SRR1766476.7871370 chr1 11522673 N chr1 11522892 N DUP 20
SRR1766482.7986008 chr1 11522833 N chr1 11522920 N DUP 20
SRR1766449.318750 chr1 11522811 N chr1 11522909 N DUP 20
SRR1766460.1744327 chr1 11522844 N chr1 11522900 N DEL 20
SRR1766482.1406693 chr1 11522733 N chr1 11522864 N DUP 31
SRR1766468.1363934 chr1 11522789 N chr1 11522964 N DUP 20
SRR1766447.966989 chr1 11522789 N chr1 11522898 N DUP 20
SRR1766461.2232196 chr1 11522757 N chr1 11522921 N DUP 21
SRR1766478.4754 chr1 11522877 N chr1 11522955 N DEL 20
SRR1766447.9072749 chr1 11522878 N chr1 11523009 N DUP 20
SRR1766483.3694014 chr1 11522801 N chr1 11522899 N DUP 20
SRR1766448.2677992 chr1 11522778 N chr1 11523010 N DEL 20
SRR1766449.9867223 chr1 11522723 N chr1 11522977 N DEL 20
SRR1766447.9072749 chr1 11522680 N chr1 11522976 N DUP 26
SRR1766469.1635488 chr1 11522779 N chr1 11523042 N DUP 20
SRR1766483.8843556 chr1 11522783 N chr1 11523103 N DEL 25
SRR1766477.6118014 chr1 11522768 N chr1 11523053 N DUP 25
SRR1766442.10152581 chr1 11522783 N chr1 11523103 N DEL 20
SRR1766475.2047625 chr1 11522871 N chr1 11523136 N DEL 26
SRR1766444.4167185 chr8 1912377 N chr8 1912659 N DEL 22
SRR1766458.5797418 chr4 6512034 N chr4 6512659 N DEL 26
SRR1766462.7526382 chr4 6511915 N chr4 6512055 N DUP 25
SRR1766443.5814116 chr4 6511768 N chr4 6512007 N DUP 21
SRR1766473.7629812 chr4 6511991 N chr4 6512443 N DUP 25
SRR1766453.7211894 chr4 6512049 N chr4 6512641 N DEL 20
SRR1766442.26404495 chr4 6512051 N chr4 6512712 N DEL 21
SRR1766462.1106642 chr4 6511695 N chr4 6511870 N DEL 20
SRR1766473.7629812 chr4 6512154 N chr4 6512515 N DEL 23
SRR1766470.1436507 chr4 6511773 N chr4 6512806 N DEL 24
SRR1766465.5187428 chr4 6511714 N chr4 6511863 N DUP 23
SRR1766442.17603216 chr4 6511789 N chr4 6512079 N DUP 26
SRR1766464.7167864 chr4 6512163 N chr4 6512662 N DEL 21
SRR1766444.2166882 chr4 6511719 N chr4 6512233 N DEL 26
SRR1766481.8785133 chr4 6511659 N chr4 6512053 N DUP 25
SRR1766455.4043507 chr4 6511719 N chr4 6511840 N DEL 20
SRR1766463.7471291 chr4 6512034 N chr4 6512803 N DEL 30
SRR1766454.1081355 chr4 6511859 N chr4 6512074 N DUP 20
SRR1766479.5221559 chr4 6511719 N chr4 6512728 N DEL 20
SRR1766442.21849030 chr4 6511794 N chr4 6512069 N DUP 21
SRR1766476.7413809 chr4 6511689 N chr4 6512509 N DEL 20
SRR1766467.924225 chr4 6511666 N chr4 6511971 N DUP 20
SRR1766444.1067630 chr4 6511948 N chr4 6512442 N DUP 20
SRR1766473.9112661 chr4 6511751 N chr4 6512551 N DUP 21
SRR1766447.6177714 chr4 6512603 N chr4 6512832 N DEL 26
SRR1766483.9989377 chr4 6511719 N chr4 6512311 N DEL 23
SRR1766471.3979794 chr4 6512051 N chr4 6512682 N DEL 25
SRR1766442.22389402 chr4 6511751 N chr4 6512062 N DUP 20
SRR1766480.1267692 chr4 6512040 N chr4 6512695 N DEL 20
SRR1766442.6046883 chr4 6512010 N chr4 6512695 N DEL 33
SRR1766467.3829509 chr4 6511718 N chr4 6512238 N DEL 25
SRR1766476.5210159 chr4 6511987 N chr4 6512040 N DUP 20
SRR1766464.1447890 chr11 134738880 N chr11 134739013 N DEL 24
SRR1766466.97568 chr11 134738880 N chr11 134739013 N DEL 24
SRR1766472.7390616 chr11 134738880 N chr11 134739013 N DEL 24
SRR1766460.1648769 chr11 134738880 N chr11 134739013 N DEL 24
SRR1766485.412779 chrX 142126133 N chrX 142126203 N DEL 23
SRR1766442.22059425 chr18 41349926 N chr18 41350003 N DUP 22
SRR1766485.9523507 chr18 41349926 N chr18 41350003 N DUP 22
SRR1766484.11242492 chr18 41349885 N chr18 41349953 N DUP 24
SRR1766482.3731191 chr18 41349926 N chr18 41350003 N DUP 21
SRR1766450.1825494 chr18 41349886 N chr18 41349996 N DUP 28
SRR1766467.5983629 chr18 41349886 N chr18 41349996 N DUP 28
SRR1766442.7309810 chr18 41349926 N chr18 41350003 N DUP 20
SRR1766446.2070074 chr18 41349926 N chr18 41350003 N DUP 29
SRR1766442.1331155 chr18 41349926 N chr18 41350003 N DUP 30
SRR1766470.9433185 chr18 41349926 N chr18 41350003 N DUP 32
SRR1766471.8057925 chr5 173128934 N chr5 173129271 N DEL 30
SRR1766461.10990412 chr5 173129209 N chr5 173129546 N DEL 20
SRR1766453.10133426 chr9 69340816 N chr9 69340939 N DUP 24
SRR1766460.3848292 chr9 69340870 N chr9 69340939 N DEL 23
SRR1766467.324415 chr9 69340843 N chr9 69340950 N DEL 38
SRR1766442.11735860 chr2 118305297 N chr2 118305361 N DEL 22
SRR1766450.9287962 chr2 118305695 N chr2 118305758 N DUP 21
SRR1766444.1566573 chr1 248522890 N chr1 248522991 N DEL 25
SRR1766476.4894098 chr18 79236837 N chr18 79237427 N DEL 25
SRR1766453.4199231 chr18 79237129 N chr18 79237508 N DEL 30
SRR1766456.3210256 chr3 127154860 N chr3 127155071 N DEL 33
SRR1766470.10505792 chr19 53990620 N chr19 53990838 N DUP 21
SRR1766471.6330094 chr19 53991104 N chr19 53991210 N DUP 22
SRR1766474.6870307 chr22 41643842 N chr22 41644169 N DEL 35
SRR1766464.6445769 chr17 82009753 N chr17 82009807 N DUP 26
SRR1766485.7290112 chr17 44984359 N chr17 44984657 N DEL 26
SRR1766456.1143039 chr17 44984734 N chr17 44985257 N DEL 30
SRR1766463.7510430 chr10 102637739 N chr10 102637791 N DUP 20
SRR1766477.7700857 chr10 102637701 N chr10 102637790 N DUP 35
SRR1766442.7307863 chr10 102637739 N chr10 102637791 N DUP 23
SRR1766449.10509094 chr10 102637739 N chr10 102637833 N DUP 21
SRR1766461.2338778 chr10 102637739 N chr10 102637791 N DUP 31
SRR1766477.4480609 chr11 101629020 N chr11 101629084 N DUP 22
SRR1766475.756274 chr2 152590090 N chr2 152590157 N DUP 22
SRR1766442.27533844 chr11 71362343 N chr11 71363366 N DEL 20
SRR1766453.2986693 chr11 71362343 N chr11 71363159 N DEL 25
SRR1766459.9383911 chr11 71362527 N chr11 71363436 N DUP 22
SRR1766474.6302661 chr11 71362527 N chr11 71363436 N DUP 22
SRR1766484.9064412 chr11 71362529 N chr11 71363207 N DUP 24
SRR1766446.4771634 chr11 71362526 N chr11 71362836 N DUP 20
SRR1766480.2108999 chr11 71362560 N chr11 71362687 N DUP 23
SRR1766485.7538658 chr11 71362652 N chr11 71363058 N DUP 25
SRR1766469.1259714 chr11 71362639 N chr11 71362893 N DUP 20
SRR1766477.11320401 chr11 71362459 N chr11 71362795 N DEL 22
SRR1766466.1682812 chr11 71362862 N chr11 71362975 N DEL 20
SRR1766466.5005942 chr11 71362698 N chr11 71362938 N DEL 20
SRR1766463.5234507 chr11 71362886 N chr11 71363047 N DEL 20
SRR1766454.4259208 chr11 71362990 N chr11 71363167 N DEL 31
SRR1766486.1892815 chr11 71363159 N chr11 71363214 N DUP 26
SRR1766442.33072783 chr11 71362866 N chr11 71363163 N DEL 26
SRR1766477.6075709 chr11 71362814 N chr11 71363181 N DUP 22
SRR1766444.5716179 chr11 71362965 N chr11 71363332 N DUP 32
SRR1766442.2535608 chr6 95502075 N chr6 95502146 N DUP 20
SRR1766445.7045337 chr6 95502145 N chr6 95502198 N DEL 34
SRR1766477.2963336 chr6 95502145 N chr6 95502198 N DEL 34
SRR1766454.2697701 chr6 95502109 N chr6 95502198 N DEL 34
SRR1766473.4780268 chr6 95502356 N chr6 95502417 N DEL 21
SRR1766455.9427814 chr6 95502060 N chr6 95502129 N DUP 25
SRR1766478.5601427 chr6 95502040 N chr6 95502569 N DUP 26
SRR1766463.4611848 chr6 95502629 N chr6 95503099 N DEL 24
SRR1766464.9675500 chr6 95502629 N chr6 95503099 N DEL 21
SRR1766468.5301496 chr6 95502629 N chr6 95503099 N DEL 21
SRR1766449.4949800 chr6 95502629 N chr6 95503099 N DEL 21
SRR1766454.9052230 chr6 95502629 N chr6 95503099 N DEL 21
SRR1766443.8918103 chr6 95503164 N chr6 95503230 N DUP 21
SRR1766442.7162371 chr6 95503164 N chr6 95503230 N DUP 26
SRR1766477.10290181 chr6 95502629 N chr6 95503099 N DEL 25
SRR1766483.10054416 chr6 95503164 N chr6 95503267 N DUP 25
SRR1766486.2662318 chr1 24907883 N chr1 24908334 N DEL 29
SRR1766450.9369944 chr1 24907883 N chr1 24908384 N DEL 24
SRR1766460.115271 chr1 24907883 N chr1 24908409 N DEL 26
SRR1766471.10855959 chr1 24907858 N chr1 24908409 N DEL 25
SRR1766470.7748660 chr1 24907864 N chr1 24908440 N DEL 20
SRR1766476.2639533 chr7 205405 N chr7 205496 N DUP 27
SRR1766466.11305139 chr7 205394 N chr7 205485 N DUP 22
SRR1766447.6251263 chr7 205394 N chr7 205485 N DUP 27
SRR1766478.4488520 chr1 125179352 N chr1 125179428 N DEL 20
SRR1766445.6516164 chr1 125179352 N chr1 125179428 N DEL 32
SRR1766467.2287342 chr1 125179358 N chr1 125179434 N DEL 23
SRR1766444.2249590 chr9 80232120 N chr9 80232234 N DEL 29
SRR1766447.10208748 chr2 3171063 N chr2 3171180 N DEL 23
SRR1766462.8992315 chr11 134760064 N chr11 134760197 N DUP 24
SRR1766466.10149980 chr11 134760067 N chr11 134760200 N DUP 24
SRR1766467.3018696 chr11 134760067 N chr11 134760200 N DUP 24
SRR1766456.3047089 chr11 134759990 N chr11 134760197 N DUP 31
SRR1766465.10897309 chr11 134760143 N chr11 134760202 N DUP 20
SRR1766467.3838176 chr11 134760143 N chr11 134760202 N DUP 37
SRR1766478.4310245 chr3 197518840 N chr3 197519251 N DEL 28
SRR1766442.23128855 chr22 18418152 N chr22 18418273 N DUP 28
SRR1766448.5933464 chr22 18418152 N chr22 18418273 N DUP 27
SRR1766472.9672541 chr22 18418214 N chr22 18418326 N DUP 20
SRR1766465.3728799 chr22 18418189 N chr22 18418266 N DUP 39
SRR1766464.5510248 chr22 18418189 N chr22 18418266 N DUP 32
SRR1766471.11937713 chr22 18418189 N chr22 18418266 N DUP 32
SRR1766447.7280118 chr22 18418189 N chr22 18418266 N DUP 26
SRR1766442.37538566 chr22 18418189 N chr22 18418266 N DUP 26
SRR1766476.9848852 chr22 18418189 N chr22 18418266 N DUP 21
SRR1766466.6327549 chr22 18418189 N chr22 18418266 N DUP 26
SRR1766458.9247823 chr22 18418189 N chr22 18418266 N DUP 22
SRR1766442.11164701 chr22 18418189 N chr22 18418266 N DUP 27
SRR1766470.5908973 chr22 18418152 N chr22 18418273 N DUP 25
SRR1766463.259549 chr18 59233851 N chr18 59233900 N DUP 25
SRR1766442.45297134 chr18 59233810 N chr18 59233931 N DUP 22
SRR1766461.10703115 chr18 59234185 N chr18 59234258 N DEL 24
SRR1766472.5458148 chr18 59234185 N chr18 59234258 N DEL 20
SRR1766446.5257225 chr12 122093067 N chr12 122093251 N DEL 21
SRR1766474.892858 chr21 5329574 N chr21 5329703 N DUP 21
SRR1766465.3153599 chr21 5329602 N chr21 5329755 N DUP 27
SRR1766457.7733511 chr11 473723 N chr11 473858 N DUP 20
SRR1766485.5375791 chr11 473723 N chr11 473858 N DUP 20
SRR1766461.8911752 chr11 473777 N chr11 473844 N DUP 24
SRR1766483.6063020 chr11 473723 N chr11 473858 N DUP 20
SRR1766463.966182 chr11 473723 N chr11 473858 N DUP 22
SRR1766446.6455652 chr2 241011227 N chr2 241011291 N DEL 28
SRR1766468.2737368 chr2 241011227 N chr2 241011291 N DEL 28
SRR1766465.9371366 chr2 241011261 N chr2 241011388 N DEL 28
SRR1766442.30844760 chr2 90383099 N chr2 90383170 N DUP 35
SRR1766454.9242232 chr2 90383099 N chr2 90383170 N DUP 35
SRR1766460.10535913 chr2 90383099 N chr2 90383170 N DUP 26
SRR1766466.6694867 chr2 90383099 N chr2 90383170 N DUP 26
SRR1766463.10078175 chr2 90383099 N chr2 90383170 N DUP 29
SRR1766484.10631252 chr2 90383099 N chr2 90383170 N DUP 30
SRR1766450.7941652 chr2 90383099 N chr2 90383170 N DUP 24
SRR1766461.3283016 chr2 90383099 N chr2 90383170 N DUP 24
SRR1766447.11136813 chr2 90383099 N chr2 90383170 N DUP 23
SRR1766475.459621 chr2 90383099 N chr2 90383170 N DUP 20
SRR1766453.8932800 chr2 90383062 N chr2 90383135 N DEL 35
SRR1766463.7684069 chr2 90383062 N chr2 90383135 N DEL 35
SRR1766481.10654764 chr2 90383062 N chr2 90383135 N DEL 35
SRR1766464.8116009 chr2 90383062 N chr2 90383135 N DEL 33
SRR1766446.2714963 chr1 3176302 N chr1 3176436 N DUP 20
SRR1766460.7839088 chr1 3176212 N chr1 3176438 N DUP 32
SRR1766444.2675616 chr6 54310807 N chr6 54310873 N DEL 20
SRR1766484.7499008 chr6 54310807 N chr6 54310873 N DEL 20
SRR1766442.7384271 chr6 54310807 N chr6 54310873 N DEL 25
SRR1766484.1628542 chr6 54310807 N chr6 54310873 N DEL 36
SRR1766444.2675616 chr6 54310807 N chr6 54310873 N DEL 20
SRR1766468.997017 chr6 54310970 N chr6 54311048 N DEL 23
SRR1766457.7498004 chr7 155354508 N chr7 155354572 N DUP 24
SRR1766460.5330172 chr7 155354508 N chr7 155354572 N DUP 24
SRR1766464.437873 chr7 155354509 N chr7 155354573 N DUP 23
SRR1766472.164914 chr7 155354509 N chr7 155354573 N DUP 23
SRR1766459.5453688 chr7 155354509 N chr7 155354573 N DUP 22
SRR1766462.1485448 chr3 98836936 N chr3 98837211 N DUP 22
SRR1766474.7634086 chr3 98836936 N chr3 98837211 N DUP 22
SRR1766473.10389319 chr3 98836936 N chr3 98837211 N DUP 22
SRR1766486.10435513 chr3 98836936 N chr3 98837211 N DUP 28
SRR1766462.809999 chr10 57693309 N chr10 57693476 N DEL 29
SRR1766461.2747020 chr10 57693403 N chr10 57693470 N DUP 32
SRR1766476.3000853 chr10 57693403 N chr10 57693470 N DUP 29
SRR1766459.6753269 chr10 57693403 N chr10 57693470 N DUP 26
SRR1766442.37999359 chr10 57693403 N chr10 57693470 N DUP 24
SRR1766442.38955487 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766472.8923067 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766477.4716957 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766453.5385784 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766455.1778743 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766448.9008293 chr10 57693434 N chr10 57693573 N DUP 24
SRR1766444.2235050 chr10 57693434 N chr10 57693573 N DUP 21
SRR1766482.3689180 chr10 57693403 N chr10 57693470 N DUP 32
SRR1766451.1700638 chr10 57693403 N chr10 57693470 N DUP 29
SRR1766453.8106407 chr10 57693403 N chr10 57693470 N DUP 29
SRR1766466.8902659 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766483.9385623 chr10 57693434 N chr10 57693559 N DUP 21
SRR1766470.9922797 chr10 57693434 N chr10 57693559 N DUP 20
SRR1766463.2489223 chr10 57693434 N chr10 57693559 N DUP 20
SRR1766483.5544864 chr10 57693434 N chr10 57693559 N DUP 20
SRR1766444.4056279 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766463.10909858 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766482.3562229 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766465.1035677 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766457.1363229 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766461.552479 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766448.3340831 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766453.8992478 chr10 57693476 N chr10 57693628 N DUP 23
SRR1766443.1159957 chr10 57693472 N chr10 57693555 N DUP 24
SRR1766459.204497 chr10 57693565 N chr10 57693737 N DEL 38
SRR1766470.4773511 chr10 57693537 N chr10 57693737 N DEL 38
SRR1766444.6954974 chr10 57693537 N chr10 57693737 N DEL 38
SRR1766461.2747020 chr10 57693537 N chr10 57693737 N DEL 38
SRR1766484.1893741 chr10 57693537 N chr10 57693737 N DEL 38
SRR1766442.17174949 chr10 57693537 N chr10 57693737 N DEL 37
SRR1766463.2226648 chr10 57693537 N chr10 57693737 N DEL 33
SRR1766467.52779 chr10 57693537 N chr10 57693737 N DEL 33
SRR1766447.3931403 chr10 57693509 N chr10 57693737 N DEL 33
SRR1766483.4020392 chr10 57693509 N chr10 57693737 N DEL 33
SRR1766448.3603075 chr10 57693363 N chr10 57693737 N DEL 20
SRR1766452.2090012 chr8 93666164 N chr8 93666243 N DEL 21
SRR1766480.886026 chr18 47982842 N chr18 47982909 N DEL 29
SRR1766458.5901849 chr2 238633800 N chr2 238634029 N DEL 21
SRR1766478.1203600 chr7 44307316 N chr7 44307574 N DEL 20
SRR1766463.5329350 chr1 194303974 N chr1 194304045 N DUP 30
SRR1766474.4138833 chr1 194303974 N chr1 194304045 N DUP 27
SRR1766461.3794238 chr1 194303974 N chr1 194304045 N DUP 25
SRR1766446.2074640 chr1 194303974 N chr1 194304045 N DUP 22
SRR1766442.33491480 chr1 194303974 N chr1 194304045 N DUP 22
SRR1766484.11718702 chr1 194303979 N chr1 194304085 N DUP 24
SRR1766477.3912043 chr1 194303974 N chr1 194304045 N DUP 22
SRR1766458.2713721 chr1 194303979 N chr1 194304085 N DUP 21
SRR1766471.1897321 chr1 194303979 N chr1 194304085 N DUP 21
SRR1766462.10934262 chr1 194303979 N chr1 194304085 N DUP 24
SRR1766483.6270725 chr1 194303981 N chr1 194304087 N DUP 24
SRR1766466.9430200 chr1 194303974 N chr1 194304045 N DUP 27
SRR1766462.10318776 chr1 194303979 N chr1 194304085 N DUP 26
SRR1766478.8008826 chr1 194303979 N chr1 194304085 N DUP 27
SRR1766453.9802769 chr15 99538164 N chr15 99538234 N DUP 30
SRR1766448.1799644 chr3 60860819 N chr3 60860911 N DUP 21
SRR1766451.5226196 chr3 60860911 N chr3 60860976 N DEL 24
SRR1766474.837542 chr3 60860911 N chr3 60860976 N DEL 27
SRR1766462.2354933 chr3 60860911 N chr3 60860976 N DEL 20
SRR1766457.1737569 chr3 60860849 N chr3 60861005 N DEL 20
SRR1766443.5382570 chr3 60861325 N chr3 60861374 N DUP 23
SRR1766472.4426684 chr3 60861363 N chr3 60861418 N DUP 32
SRR1766475.7945408 chr3 60861363 N chr3 60861418 N DUP 30
SRR1766462.5828437 chr3 60861363 N chr3 60861418 N DUP 30
SRR1766478.6821376 chr9 137346675 N chr9 137346755 N DUP 25
SRR1766482.9248942 chr9 137346675 N chr9 137346755 N DUP 29
SRR1766456.5732290 chr9 137346675 N chr9 137346755 N DUP 31
SRR1766449.1322370 chr9 137346675 N chr9 137346755 N DUP 32
SRR1766442.17412559 chr9 137346675 N chr9 137346755 N DUP 34
SRR1766479.3488358 chr2 117643563 N chr2 117643630 N DUP 26
SRR1766459.3930887 chr2 117643612 N chr2 117643716 N DEL 22
SRR1766478.2952910 chr2 117643563 N chr2 117643630 N DUP 26
SRR1766475.72241 chr7 98242729 N chr7 98243136 N DUP 23
SRR1766446.3423439 chr7 98242729 N chr7 98243136 N DUP 26
SRR1766452.5261696 chr7 98242901 N chr7 98243073 N DUP 23
SRR1766477.7985835 chr14 105693773 N chr14 105693850 N DUP 30
SRR1766485.5430354 chr14 105693685 N chr14 105693776 N DUP 23
SRR1766452.9897100 chr1 2977693 N chr1 2977772 N DUP 34
SRR1766450.1049268 chr7 62442454 N chr7 62442698 N DUP 21
SRR1766471.2210920 chr7 62442660 N chr7 62442734 N DUP 25
SRR1766467.9128986 chr2 64375753 N chr2 64376213 N DEL 24
SRR1766443.179353 chr2 64375753 N chr2 64376213 N DEL 29
SRR1766461.8014131 chr2 64375795 N chr2 64376208 N DEL 24
SRR1766480.2497720 chr2 64375813 N chr2 64376039 N DEL 24
SRR1766455.3924306 chr2 64375967 N chr2 64376219 N DEL 29
SRR1766478.9075524 chr2 64375947 N chr2 64376018 N DEL 22
SRR1766471.8460006 chrX 35692462 N chrX 35692559 N DUP 31
SRR1766483.6209409 chrX 35692537 N chrX 35692610 N DUP 31
SRR1766477.7315024 chrX 35692492 N chrX 35692559 N DUP 28
SRR1766475.7968703 chrX 35692492 N chrX 35692559 N DUP 34
SRR1766455.386080 chrX 35692492 N chrX 35692559 N DUP 31
SRR1766477.943855 chrX 35692503 N chrX 35692560 N DUP 20
SRR1766468.1854140 chr1 8301316 N chr1 8301597 N DEL 34
SRR1766468.1854140 chr1 8301301 N chr1 8301582 N DEL 21
SRR1766480.6327103 chr1 8301521 N chr1 8301634 N DEL 20
SRR1766445.7914758 chr1 8301785 N chr1 8301952 N DUP 30
SRR1766477.4719669 chr1 8301483 N chr1 8301848 N DEL 25
SRR1766472.6181988 chr1 8301851 N chr1 8301934 N DUP 30
SRR1766461.8633633 chr1 8301486 N chr1 8301851 N DEL 20
SRR1766460.2163640 chr8 132187901 N chr8 132187983 N DEL 25
SRR1766484.7138450 chr5 180615503 N chr5 180615562 N DEL 22
SRR1766455.198855 chr5 180615465 N chr5 180615624 N DUP 30
SRR1766444.6610758 chr5 180615317 N chr5 180615522 N DUP 20
SRR1766481.6316063 chr5 180615420 N chr5 180615611 N DUP 24
SRR1766465.6219816 chr22 18370651 N chr22 18370706 N DEL 25
SRR1766478.11701309 chr10 2871852 N chr10 2871910 N DEL 37
SRR1766442.17362191 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766450.2437205 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766451.10089738 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766485.9023809 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766456.4442558 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766461.388165 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766449.9118484 chr10 83585241 N chr10 83585319 N DEL 31
SRR1766484.2236619 chr10 83585233 N chr10 83585348 N DUP 21
SRR1766456.5063869 chr22 32329881 N chr22 32330167 N DUP 21
SRR1766451.6534568 chr22 32330100 N chr22 32331304 N DEL 29
SRR1766461.6554851 chr9 89671689 N chr9 89671819 N DEL 32
SRR1766442.27168270 chr9 89671692 N chr9 89671871 N DUP 20
SRR1766453.6777803 chr9 89671710 N chr9 89671868 N DUP 27
SRR1766455.4344450 chr9 89671692 N chr9 89671937 N DUP 23
SRR1766464.1845413 chr9 89671770 N chr9 89671877 N DUP 20
SRR1766473.5048874 chr9 89671713 N chr9 89671871 N DUP 27
SRR1766481.97153 chr9 89671770 N chr9 89671826 N DUP 23
SRR1766459.10678798 chr9 89671692 N chr9 89671837 N DUP 24
SRR1766455.1511834 chr9 89671818 N chr9 89671874 N DUP 22
SRR1766475.9514433 chr9 89671772 N chr9 89671849 N DUP 20
SRR1766473.5048874 chr9 89671770 N chr9 89671877 N DUP 24
SRR1766450.7868999 chr9 89671729 N chr9 89671833 N DUP 23
SRR1766481.10663315 chr9 89671770 N chr9 89671877 N DUP 22
SRR1766450.5021997 chr9 89671692 N chr9 89671802 N DUP 23
SRR1766478.9056447 chr9 89671770 N chr9 89671877 N DUP 26
SRR1766449.1978826 chr9 89671818 N chr9 89671874 N DUP 27
SRR1766471.4303433 chr9 89671738 N chr9 89671893 N DUP 24
SRR1766447.443044 chr9 89671770 N chr9 89671877 N DUP 28
SRR1766482.5794508 chr9 89671692 N chr9 89671853 N DUP 31
SRR1766474.7663017 chr22 36434342 N chr22 36434399 N DUP 22
SRR1766448.9788747 chr1 96153244 N chr1 96153309 N DUP 25
SRR1766450.8675057 chr1 96153244 N chr1 96153309 N DUP 32
SRR1766444.6197180 chr1 96153244 N chr1 96153309 N DUP 30
SRR1766445.10309417 chr1 96153244 N chr1 96153309 N DUP 29
SRR1766481.11244748 chr1 96153244 N chr1 96153309 N DUP 25
SRR1766443.9470226 chr1 96153244 N chr1 96153309 N DUP 25
SRR1766442.9972324 chr1 96153244 N chr1 96153309 N DUP 25
SRR1766475.5016149 chr1 96153244 N chr1 96153309 N DUP 23
SRR1766476.10068121 chr1 96153244 N chr1 96153309 N DUP 20
SRR1766482.12656170 chr1 96153244 N chr1 96153309 N DUP 26
SRR1766471.11558901 chr1 96153244 N chr1 96153309 N DUP 30
SRR1766479.8424729 chr1 96153244 N chr1 96153309 N DUP 30
SRR1766479.11251285 chr20 22378581 N chr20 22378638 N DEL 20
SRR1766469.8627368 chr20 22378581 N chr20 22378638 N DEL 25
SRR1766467.375395 chr7 72255269 N chr7 72255599 N DEL 20
SRR1766482.8965201 chr4 1652601 N chr4 1652972 N DEL 22
SRR1766463.5418275 chr6 104424259 N chr6 104424400 N DEL 25
SRR1766457.7759522 chr3 181743053 N chr3 181743112 N DUP 25
SRR1766447.1495805 chr19 108019 N chr19 108076 N DUP 20
SRR1766461.3872695 chr19 107980 N chr19 108037 N DUP 25
SRR1766462.8314030 chr19 108019 N chr19 108076 N DUP 23
SRR1766475.1018103 chr19 107980 N chr19 108037 N DUP 28
SRR1766472.10946882 chr19 107980 N chr19 108081 N DUP 20
SRR1766461.7452503 chr19 107980 N chr19 108081 N DUP 22
SRR1766445.5725495 chr19 107980 N chr19 108081 N DUP 28
SRR1766448.6909808 chr19 108001 N chr19 108106 N DUP 27
SRR1766445.641220 chr19 108001 N chr19 108106 N DUP 28
SRR1766477.9531331 chr19 108014 N chr19 108167 N DUP 24
SRR1766472.8870166 chr19 108014 N chr19 108167 N DUP 29
SRR1766460.1082899 chr6 38103619 N chr6 38103674 N DEL 37
SRR1766483.1665888 chr6 38103619 N chr6 38103674 N DEL 33
SRR1766448.7012654 chr6 38103619 N chr6 38103674 N DEL 32
SRR1766474.7268480 chr6 38103619 N chr6 38103674 N DEL 30
SRR1766442.11322981 chr6 38103619 N chr6 38103674 N DEL 30
SRR1766455.3486668 chr6 25206656 N chr6 25206733 N DUP 24
SRR1766451.4105653 chr6 25206681 N chr6 25206731 N DUP 27
SRR1766469.1862069 chr6 25206656 N chr6 25206733 N DUP 24
SRR1766465.9915501 chr6 25206713 N chr6 25206784 N DUP 27
SRR1766457.2866596 chr6 25206713 N chr6 25206784 N DUP 25
SRR1766461.6166102 chrX 114387045 N chrX 114387676 N DUP 23
SRR1766450.6626251 chrX 114387120 N chrX 114387406 N DEL 20
SRR1766455.3927219 chrX 114387148 N chrX 114387240 N DEL 20
SRR1766445.2706233 chrX 114387199 N chrX 114387641 N DUP 28
SRR1766454.9028196 chrX 114387199 N chrX 114387641 N DUP 26
SRR1766445.9650319 chrX 114387221 N chrX 114387385 N DUP 20
SRR1766479.6862988 chrX 114387308 N chrX 114387474 N DUP 21
SRR1766453.5861128 chrX 114387059 N chrX 114387183 N DUP 20
SRR1766447.986226 chrX 114387221 N chrX 114387385 N DUP 20
SRR1766481.5985479 chrX 114387221 N chrX 114387385 N DUP 21
SRR1766477.10961291 chrX 114387199 N chrX 114387641 N DUP 23
SRR1766467.1549694 chrX 114387386 N chrX 114387585 N DUP 22
SRR1766447.11354775 chr12 132621012 N chr12 132621074 N DEL 24
SRR1766442.25929985 chr19 480906 N chr19 481059 N DEL 23
SRR1766459.10428478 chr19 480788 N chr19 481623 N DEL 20
SRR1766442.29871329 chr19 481321 N chr19 481648 N DEL 20
SRR1766486.9812069 chr11 131680938 N chr11 131681523 N DUP 20
SRR1766471.9004494 chr11 131680960 N chr11 131681797 N DEL 20
SRR1766443.2736729 chr20 18023106 N chr20 18023460 N DEL 20
SRR1766469.8867015 chr19 16379957 N chr19 16380289 N DEL 20
SRR1766484.8151235 chr19 16379850 N chr19 16380293 N DEL 25
SRR1766458.332714 chr3 134701429 N chr3 134701482 N DUP 22
SRR1766483.5989940 chr3 134701429 N chr3 134701482 N DUP 22
SRR1766473.3623053 chr3 134701427 N chr3 134701504 N DUP 34
SRR1766457.7995779 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766477.7775706 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766459.4379318 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766470.6180568 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766474.10151694 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766471.9587337 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766452.1432668 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766442.41086000 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766445.5422077 chr3 134701427 N chr3 134701504 N DUP 36
SRR1766480.293217 chr20 60501332 N chr20 60501533 N DEL 20
