SRR1766473.9568686 chr6 40209174 N chr6 40209625 N DEL 10
SRR1766462.670452 chr6 40209145 N chr6 40209198 N DUP 14
SRR1766473.4075371 chr6 40209145 N chr6 40209198 N DUP 14
SRR1766477.890951 chr6 40209145 N chr6 40209198 N DUP 14
SRR1766457.549986 chr6 40209145 N chr6 40209198 N DUP 14
SRR1766447.3435014 chr6 40209145 N chr6 40209198 N DUP 10
SRR1766446.7051739 chr6 40209154 N chr6 40209913 N DUP 18
SRR1766447.9882624 chr6 40209134 N chr6 40209197 N DUP 14
SRR1766457.4275394 chr6 40209138 N chr6 40209275 N DUP 11
SRR1766460.3882408 chr6 40209227 N chr6 40209914 N DUP 17
SRR1766456.5530273 chr6 40209275 N chr6 40209364 N DEL 17
SRR1766486.8209297 chr6 40209227 N chr6 40209606 N DUP 14
SRR1766457.4145131 chr6 40209161 N chr6 40209718 N DUP 10
SRR1766462.7242706 chr6 40209314 N chr6 40209409 N DEL 16
SRR1766485.9634000 chr6 40209227 N chr6 40209606 N DUP 11
SRR1766478.7536017 chr6 40209309 N chr6 40209422 N DEL 13
SRR1766447.9326736 chr6 40209275 N chr6 40209364 N DEL 17
SRR1766463.815128 chr6 40209192 N chr6 40209273 N DEL 15
SRR1766454.1184692 chr6 40209226 N chr6 40209693 N DEL 11
SRR1766453.3507462 chr6 40209389 N chr6 40209866 N DEL 19
SRR1766453.1306798 chr6 40209557 N chr6 40209782 N DUP 17
SRR1766479.11915969 chr6 40209557 N chr6 40209782 N DUP 17
SRR1766482.13049617 chr6 40209435 N chr6 40209568 N DUP 11
SRR1766447.9305880 chr6 40209172 N chr6 40209646 N DEL 14
SRR1766455.1378690 chr6 40209699 N chr6 40209910 N DUP 17
SRR1766455.7600844 chr6 40209710 N chr6 40209933 N DUP 17
SRR1766461.225301 chr6 40209766 N chr6 40209863 N DUP 19
SRR1766473.9568686 chr6 40209766 N chr6 40209863 N DUP 19
SRR1766454.7893747 chr6 40209767 N chr6 40209864 N DUP 17
SRR1766454.2849246 chr6 40209810 N chr6 40209905 N DUP 12
SRR1766460.7018530 chr6 40209521 N chr6 40209914 N DUP 17
SRR1766482.5377961 chr6 40209566 N chr6 40209751 N DEL 16
SRR1766466.1461148 chr6 40209513 N chr6 40209900 N DUP 14
SRR1766451.3569801 chr6 40209440 N chr6 40209555 N DUP 17
SRR1766449.601789 chr6 40209545 N chr6 40209792 N DEL 10
SRR1766451.3864695 chr6 40209512 N chr6 40209899 N DUP 11
SRR1766476.2995335 chr6 40209512 N chr6 40209899 N DUP 11
SRR1766472.10092431 chr6 40209486 N chr6 40209883 N DUP 17
SRR1766467.2602274 chr6 40209520 N chr6 40209921 N DUP 11
SRR1766484.202117 chr6 40209545 N chr6 40209792 N DEL 10
SRR1766442.25191808 chr6 40209521 N chr6 40209914 N DUP 17
SRR1766445.4999125 chr6 40209512 N chr6 40209899 N DUP 16
SRR1766458.1050790 chr6 40209513 N chr6 40209900 N DUP 12
SRR1766484.3925706 chr6 40209513 N chr6 40209900 N DUP 13
SRR1766442.12541431 chr6 40209810 N chr6 40209913 N DUP 19
SRR1766473.6636659 chr6 40209605 N chr6 40209864 N DEL 18
SRR1766450.8524 chr6 40209605 N chr6 40209864 N DEL 18
SRR1766442.20536606 chr6 40209605 N chr6 40209864 N DEL 17
SRR1766471.2270222 chr6 40209161 N chr6 40209864 N DEL 14
SRR1766442.27668881 chr6 40209535 N chr6 40209864 N DEL 12
SRR1766443.296974 chr6 40209787 N chr6 40209912 N DEL 13
SRR1766473.9221763 chr6 40209554 N chr6 40209889 N DEL 11
SRR1766442.37302361 chr6 40209744 N chr6 40209903 N DEL 19
SRR1766460.3882408 chr6 40209744 N chr6 40209903 N DEL 18
SRR1766455.1329637 chr6 40209744 N chr6 40209903 N DEL 18
SRR1766475.10669225 chr6 40209765 N chr6 40209908 N DEL 16
SRR1766442.26017208 chr6 40209744 N chr6 40209903 N DEL 18
SRR1766473.680692 chr6 40209744 N chr6 40209903 N DEL 18
SRR1766470.8625940 chr6 40209491 N chr6 40209896 N DEL 14
SRR1766444.2979777 chr6 40209154 N chr6 40209913 N DEL 18
SRR1766482.2261671 chr6 40209154 N chr6 40209913 N DEL 18
SRR1766467.5781574 chr6 40209144 N chr6 40209913 N DEL 15
SRR1766442.21006621 chr6 40209144 N chr6 40209913 N DEL 12
SRR1766454.1072266 chr10 1409628 N chr10 1409861 N DUP 10
SRR1766480.2458580 chr7 57927384 N chr7 57928234 N DUP 14
SRR1766485.3726830 chr7 57928293 N chr7 57928807 N DEL 17
SRR1766472.10424680 chr7 57927521 N chr7 57928541 N DEL 11
SRR1766458.1129689 chr7 57927457 N chr7 57928646 N DUP 13
SRR1766454.9642876 chr7 57928584 N chr7 57928756 N DEL 15
SRR1766461.10244698 chr7 57928741 N chr7 57928913 N DEL 13
SRR1766443.5158616 chr2 10015574 N chr2 10015631 N DUP 10
SRR1766442.39674558 chr2 10015560 N chr2 10015648 N DEL 10
SRR1766442.22180632 chr2 10015549 N chr2 10015724 N DEL 10
SRR1766444.5811458 chr2 10015461 N chr2 10015820 N DUP 14
SRR1766453.2312095 chr2 10015549 N chr2 10015724 N DEL 10
SRR1766482.3981777 chr2 10015503 N chr2 10015874 N DUP 10
SRR1766461.3630218 chr2 10015560 N chr2 10015834 N DEL 10
SRR1766455.6460420 chr2 10015856 N chr2 10016256 N DUP 10
SRR1766450.387849 chr2 10015545 N chr2 10015889 N DEL 12
SRR1766472.2917252 chr2 10015538 N chr2 10015911 N DEL 10
SRR1766483.12509417 chr2 10015665 N chr2 10015893 N DEL 11
SRR1766448.3180146 chr2 10015562 N chr2 10015935 N DEL 10
SRR1766450.7506182 chr2 10015632 N chr2 10015918 N DEL 18
SRR1766461.10190401 chr2 10015480 N chr2 10015940 N DEL 12
SRR1766484.4623757 chr5 92251214 N chr5 92251265 N DUP 13
SRR1766442.10696079 chr5 92251214 N chr5 92251265 N DUP 13
SRR1766485.4612852 chr5 92251214 N chr5 92251265 N DUP 13
SRR1766442.36759277 chr5 92251454 N chr5 92251513 N DUP 12
SRR1766482.6350970 chr5 92251454 N chr5 92251513 N DUP 13
SRR1766450.10885329 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766484.8893486 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766447.9303687 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766477.6271903 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766476.4404715 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766472.6831349 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766470.6645822 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766443.2272923 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766471.11106732 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766475.9824406 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766459.7837757 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766454.5150949 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766442.39144130 chr5 92251472 N chr5 92251567 N DUP 11
SRR1766481.7325313 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766476.166040 chr5 92251472 N chr5 92251567 N DUP 11
SRR1766447.4120250 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766484.2954826 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766479.9735463 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766477.9224121 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766471.3081370 chr5 92251472 N chr5 92251567 N DUP 11
SRR1766442.15349372 chr5 92251472 N chr5 92251533 N DUP 11
SRR1766458.8518665 chr10 36190353 N chr10 36190404 N DEL 11
SRR1766470.8866232 chr10 36190358 N chr10 36190409 N DEL 10
SRR1766458.9133773 chr15 21777133 N chr15 21777482 N DEL 10
SRR1766464.10702561 chr15 21777136 N chr15 21777485 N DEL 15
SRR1766461.1182085 chr2 208177089 N chr2 208177164 N DEL 19
SRR1766472.3314723 chr2 208177089 N chr2 208177164 N DEL 19
SRR1766443.212780 chr19 40350033 N chr19 40350336 N DEL 15
SRR1766484.2812032 chr19 40349896 N chr19 40350199 N DEL 10
SRR1766442.17693725 chr19 40349973 N chr19 40350276 N DEL 10
SRR1766473.7750635 chr19 40349984 N chr19 40350287 N DEL 19
SRR1766445.7894087 chr4 95192460 N chr4 95192556 N DEL 10
SRR1766471.6046448 chr19 36796431 N chr19 36796482 N DEL 11
SRR1766456.1922052 chr9 65398366 N chr9 65398565 N DEL 12
SRR1766475.8026983 chr2 216226465 N chr2 216226563 N DUP 12
SRR1766444.728493 chrX 21731630 N chrX 21731720 N DEL 16
SRR1766442.8330757 chrX 21731713 N chrX 21731848 N DUP 11
SRR1766479.957156 chrX 21731713 N chrX 21731848 N DUP 14
SRR1766481.4382009 chr9 43335699 N chr9 43335824 N DEL 15
SRR1766475.7535635 chr9 43335699 N chr9 43335824 N DEL 15
SRR1766486.1965635 chr9 43335699 N chr9 43335824 N DEL 15
SRR1766470.10134647 chr8 121201380 N chr8 121201459 N DUP 10
SRR1766456.643668 chr8 121201378 N chr8 121201457 N DUP 15
SRR1766448.8348723 chr8 121201479 N chr8 121201666 N DUP 10
SRR1766474.2896056 chr8 121201769 N chr8 121201834 N DEL 18
SRR1766479.3003673 chr8 121201769 N chr8 121201834 N DEL 15
SRR1766460.3454021 chr8 121201770 N chr8 121201835 N DEL 14
SRR1766453.7944451 chr8 121201770 N chr8 121201835 N DEL 14
SRR1766442.21275634 chr2 205380379 N chr2 205380612 N DEL 13
SRR1766470.1516395 chr2 205380379 N chr2 205380612 N DEL 13
SRR1766464.9212812 chr2 205380379 N chr2 205380612 N DEL 17
SRR1766474.8397851 chr2 205380379 N chr2 205380612 N DEL 18
SRR1766444.6049303 chr2 205380379 N chr2 205380612 N DEL 18
SRR1766483.5358359 chr2 205380533 N chr2 205380633 N DUP 12
SRR1766448.3783836 chr2 205380387 N chr2 205380751 N DUP 10
SRR1766465.2096849 chr2 205380489 N chr2 205380622 N DEL 15
SRR1766474.4326775 chr2 205380379 N chr2 205380612 N DEL 17
SRR1766484.291650 chr2 205380384 N chr2 205380617 N DEL 10
SRR1766472.3022630 chr2 205380379 N chr2 205380612 N DEL 17
SRR1766469.5152683 chr2 205380453 N chr2 205380688 N DUP 10
SRR1766457.1764423 chr2 205381058 N chr2 205381115 N DEL 12
SRR1766471.4466941 chr2 205380388 N chr2 205381064 N DUP 14
SRR1766459.1387881 chr2 205380418 N chr2 205381046 N DEL 15
SRR1766461.3065168 chr2 201283099 N chr2 201283548 N DEL 12
SRR1766458.8789487 chr2 201283099 N chr2 201283548 N DEL 12
SRR1766479.6378661 chr2 201283099 N chr2 201283548 N DEL 12
SRR1766461.3065168 chr2 201283100 N chr2 201283549 N DEL 11
SRR1766475.7774262 chr7 157994720 N chr7 157995450 N DUP 12
SRR1766454.6011466 chr7 157994771 N chr7 157994852 N DUP 18
SRR1766462.1996092 chr7 157994867 N chr7 157995235 N DEL 10
SRR1766456.4570169 chr7 157994892 N chr7 157995219 N DEL 12
SRR1766466.4874667 chr7 157994850 N chr7 157995218 N DEL 12
SRR1766461.5777529 chr7 157994809 N chr7 157995218 N DEL 12
SRR1766478.1115482 chr7 157994858 N chr7 157995226 N DEL 12
SRR1766476.6885246 chr7 157994850 N chr7 157995218 N DEL 11
SRR1766478.6885597 chr7 157994835 N chr7 157995244 N DEL 11
SRR1766442.12778434 chr7 157994870 N chr7 157995278 N DEL 10
SRR1766442.16096874 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766447.1575509 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766453.8522873 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766445.9125244 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766471.1777261 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766442.45549660 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766455.2898692 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766462.4787455 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766459.2785444 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766451.2213510 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766470.4532228 chr2 36182231 N chr2 36182304 N DEL 10
SRR1766449.1846243 chr2 36182257 N chr2 36182400 N DUP 10
SRR1766467.665054 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766478.4081387 chr2 36182309 N chr2 36182414 N DUP 12
SRR1766447.1916193 chr2 36182257 N chr2 36182400 N DUP 10
SRR1766467.7387588 chrX 738954 N chrX 739063 N DEL 10
SRR1766444.610448 chr21 45452872 N chr21 45453134 N DUP 12
SRR1766467.3745615 chr21 45452872 N chr21 45453134 N DUP 12
SRR1766462.7819178 chr20 53837892 N chr20 53837947 N DUP 18
SRR1766451.2412593 chr20 53837892 N chr20 53837947 N DUP 13
SRR1766463.9996456 chr1 42324194 N chr1 42324285 N DEL 15
SRR1766481.9989619 chr1 42324217 N chr1 42324308 N DEL 10
SRR1766448.19336 chr1 42324204 N chr1 42324293 N DUP 18
SRR1766485.648402 chr1 42324204 N chr1 42324293 N DUP 18
SRR1766455.5763460 chr1 42324204 N chr1 42324293 N DUP 10
SRR1766444.5503561 chr1 42324204 N chr1 42324293 N DUP 12
SRR1766442.5989375 chr6 65443284 N chr6 65443347 N DUP 11
SRR1766442.3554828 chr6 65443311 N chr6 65443378 N DEL 11
SRR1766443.6485012 chr6 65443311 N chr6 65443378 N DEL 11
SRR1766442.31688981 chr6 65443311 N chr6 65443378 N DEL 11
SRR1766457.2957956 chr6 65443311 N chr6 65443378 N DEL 10
SRR1766453.7950980 chr6 65443311 N chr6 65443378 N DEL 10
SRR1766455.6205566 chr2 238769437 N chr2 238769550 N DEL 13
SRR1766450.7920914 chr4 3919305 N chr4 3919454 N DEL 11
SRR1766480.7368196 chr5 158582707 N chr5 158583006 N DUP 10
SRR1766452.72925 chr5 158582999 N chr5 158583323 N DEL 10
SRR1766456.6188695 chr5 158583151 N chr5 158583375 N DUP 15
SRR1766472.930962 chr5 158582986 N chr5 158583582 N DUP 10
SRR1766449.8637137 chrX 62523322 N chrX 62523832 N DEL 10
SRR1766485.6609093 chrX 62523940 N chrX 62524112 N DEL 10
SRR1766480.1648543 chrX 62523355 N chrX 62523525 N DUP 10
SRR1766460.3028012 chr15 78373872 N chr15 78373925 N DUP 10
SRR1766442.18635948 chr5 145742265 N chr5 145742354 N DEL 12
SRR1766461.4868162 chr5 145742264 N chr5 145742353 N DEL 13
SRR1766457.5094193 chr7 155932809 N chr7 155933018 N DEL 13
SRR1766467.402072 chr7 155932809 N chr7 155933018 N DEL 19
SRR1766482.5016453 chr7 155932809 N chr7 155933018 N DEL 16
SRR1766451.7273075 chr21 42349289 N chr21 42349366 N DUP 10
SRR1766480.219519 chr5 117993527 N chr5 117993580 N DEL 12
SRR1766446.1599666 chr5 117993527 N chr5 117993580 N DEL 13
SRR1766457.2030254 chr1 154714109 N chr1 154714339 N DUP 14
SRR1766477.749271 chr1 154714331 N chr1 154714762 N DUP 17
SRR1766455.3191781 chr1 154714319 N chr1 154714691 N DUP 10
SRR1766444.1959785 chr1 154714375 N chr1 154714618 N DUP 10
SRR1766469.2821435 chr1 154714381 N chr1 154714432 N DUP 11
SRR1766442.40563046 chr1 154714349 N chr1 154714427 N DEL 10
SRR1766486.2104134 chr1 154714468 N chr1 154714535 N DUP 15
SRR1766468.2370654 chr1 154714451 N chr1 154714631 N DUP 16
SRR1766453.2898949 chr1 154714526 N chr1 154714703 N DUP 11
SRR1766475.6450498 chr1 154714290 N chr1 154714532 N DEL 11
SRR1766485.75103 chr1 154714183 N chr1 154714580 N DEL 13
SRR1766448.9273968 chr1 154714195 N chr1 154714762 N DEL 11
SRR1766470.2783005 chr1 154714599 N chr1 154714784 N DEL 12
SRR1766478.504357 chr1 154714352 N chr1 154714749 N DEL 10
SRR1766462.8055582 chr16 34696431 N chr16 34696482 N DUP 10
SRR1766442.12016444 chr16 34696431 N chr16 34696482 N DUP 12
SRR1766465.2750913 chr16 34696431 N chr16 34696482 N DUP 16
SRR1766480.2862494 chr18 76587059 N chr18 76587281 N DEL 15
SRR1766442.29225713 chr18 76587139 N chr18 76587293 N DEL 10
SRR1766467.3619138 chr18 76587029 N chr18 76587319 N DEL 11
SRR1766446.1731880 chr16 89995295 N chr16 89995441 N DUP 10
SRR1766442.13571049 chr13 108258351 N chr13 108258400 N DUP 10
SRR1766478.8389258 chr13 108258351 N chr13 108258400 N DUP 10
SRR1766482.3535483 chr13 108258351 N chr13 108258400 N DUP 11
SRR1766476.11208833 chr13 108258351 N chr13 108258400 N DUP 12
SRR1766482.2054380 chr13 108258351 N chr13 108258400 N DUP 14
SRR1766462.6406353 chr13 108258355 N chr13 108258404 N DUP 11
SRR1766462.7163229 chr6 87128940 N chr6 87129013 N DEL 10
SRR1766463.9171038 chr6 87128940 N chr6 87129013 N DEL 10
SRR1766483.10743055 chr6 87129128 N chr6 87129195 N DEL 11
SRR1766443.3975051 chr6 87129128 N chr6 87129195 N DEL 13
SRR1766486.447320 chr6 87129198 N chr6 87129265 N DUP 14
SRR1766449.1395501 chr17 79709889 N chr17 79710414 N DEL 17
SRR1766464.3869662 chr17 79709801 N chr17 79710414 N DEL 10
SRR1766484.9346968 chr1 3502173 N chr1 3502251 N DUP 17
SRR1766454.8844611 chr1 243480544 N chr1 243480982 N DUP 19
SRR1766483.6288009 chr1 243480793 N chr1 243481044 N DUP 18
SRR1766470.6972473 chr1 243480740 N chr1 243480906 N DEL 14
SRR1766462.7343981 chr1 243480580 N chr1 243480923 N DEL 10
SRR1766448.10728698 chr1 243480839 N chr1 243481059 N DEL 12
SRR1766472.3168133 chr9 24739245 N chr9 24739363 N DUP 10
SRR1766467.321575 chr17 68001923 N chr17 68002228 N DEL 10
SRR1766474.4290743 chr17 68002099 N chr17 68002400 N DEL 11
SRR1766442.25779218 chr17 68002245 N chr17 68002555 N DEL 10
SRR1766471.6344186 chr17 68002451 N chr17 68003116 N DEL 10
SRR1766479.4092345 chr17 68002232 N chr17 68003204 N DUP 10
SRR1766470.8696700 chr1 1192538 N chr1 1192755 N DEL 10
SRR1766479.13223392 chr1 1192538 N chr1 1192926 N DEL 10
SRR1766443.1267782 chr1 1192725 N chr1 1192921 N DEL 10
SRR1766469.2894144 chr1 1192610 N chr1 1192827 N DEL 10
SRR1766471.1972827 chr1 1192617 N chr1 1192834 N DEL 15
SRR1766449.8500478 chr1 1192593 N chr1 1192834 N DEL 15
SRR1766462.4778579 chr1 1192617 N chr1 1192858 N DEL 11
SRR1766442.13628522 chr10 132605310 N chr10 132605568 N DUP 10
SRR1766456.4023159 chr16 89074320 N chr16 89074555 N DEL 16
SRR1766450.3307004 chr16 89074290 N chr16 89074555 N DEL 10
SRR1766442.29339462 chr10 132965341 N chr10 132965854 N DEL 10
SRR1766466.2426217 chr13 58176976 N chr13 58177042 N DUP 12
SRR1766462.10163603 chr17 2034659 N chr17 2034891 N DEL 10
SRR1766481.13234930 chr19 52554561 N chr19 52555318 N DEL 10
SRR1766446.2265413 chr19 52554136 N chr19 52554809 N DEL 12
SRR1766459.8336534 chr5 40697200 N chr5 40697301 N DEL 12
SRR1766479.99536 chr5 40697251 N chr5 40697306 N DUP 10
SRR1766443.9554326 chr5 40697251 N chr5 40697306 N DUP 10
SRR1766442.31258665 chr5 40697251 N chr5 40697306 N DUP 10
SRR1766467.8179777 chr5 40697251 N chr5 40697306 N DUP 10
SRR1766477.8398286 chr5 40697252 N chr5 40697307 N DUP 10
SRR1766459.4474013 chr10 26811890 N chr10 26811945 N DEL 10
SRR1766460.9439543 chr10 26811890 N chr10 26811945 N DEL 10
SRR1766475.7417461 chr9 43326702 N chr9 43326951 N DEL 11
SRR1766451.9390055 chr6 1054136 N chr6 1054188 N DUP 16
SRR1766453.9027704 chr22 48757290 N chr22 48757507 N DUP 12
SRR1766450.387174 chr22 48757463 N chr22 48757566 N DUP 17
SRR1766458.6284656 chr22 48757304 N chr22 48757482 N DUP 10
SRR1766476.3236244 chr22 48757482 N chr22 48757549 N DUP 15
SRR1766451.7704511 chr22 48757482 N chr22 48757549 N DUP 15
SRR1766483.9939486 chr22 48757482 N chr22 48757588 N DUP 10
SRR1766442.12723009 chr1 55662714 N chr1 55662790 N DUP 10
SRR1766482.8429665 chr1 55662714 N chr1 55662790 N DUP 11
SRR1766467.9973048 chr1 55662714 N chr1 55662790 N DUP 17
SRR1766471.415555 chr8 93833420 N chr8 93833802 N DEL 10
SRR1766476.11267475 chr8 93833416 N chr8 93833798 N DEL 19
SRR1766469.4498363 chr8 93833457 N chr8 93833802 N DEL 11
SRR1766454.10260786 chr8 93833694 N chr8 93833808 N DEL 10
SRR1766457.2120505 chr8 93833788 N chr8 93834010 N DEL 15
SRR1766442.12588855 chr8 93833857 N chr8 93834409 N DEL 10
SRR1766444.4475118 chr8 93833718 N chr8 93834053 N DEL 17
SRR1766478.7566217 chr8 93834418 N chr8 93834525 N DUP 11
SRR1766445.2625664 chr8 93834566 N chr8 93834645 N DUP 10
SRR1766478.6747538 chr8 93834691 N chr8 93834883 N DEL 10
SRR1766442.13569260 chr8 93834718 N chr8 93834833 N DEL 16
SRR1766478.11142125 chr18 29511662 N chr18 29511838 N DEL 15
SRR1766476.7549764 chr18 29511662 N chr18 29511838 N DEL 12
SRR1766484.5172379 chr18 29511787 N chr18 29512116 N DEL 12
SRR1766476.2134445 chr18 29511761 N chr18 29512116 N DEL 12
SRR1766442.3639045 chr18 29511761 N chr18 29512116 N DEL 11
SRR1766455.7116177 chr18 29512204 N chr18 29512344 N DUP 13
SRR1766467.292615 chr18 29512204 N chr18 29512344 N DUP 14
SRR1766450.9692300 chr18 29511751 N chr18 29512205 N DEL 12
SRR1766466.1942525 chr18 29511666 N chr18 29512204 N DEL 14
SRR1766475.5918332 chr18 29511666 N chr18 29512204 N DEL 18
SRR1766485.12004081 chr18 29511666 N chr18 29512230 N DEL 14
SRR1766484.9098791 chr4 162764116 N chr4 162764199 N DEL 12
SRR1766456.815454 chr4 162764125 N chr4 162764199 N DEL 14
SRR1766447.7595681 chr4 162764125 N chr4 162764199 N DEL 14
SRR1766470.9437047 chr14 67700868 N chr14 67701174 N DEL 11
SRR1766480.878275 chr10 68503004 N chr10 68503089 N DEL 12
SRR1766461.10562237 chr6 994146 N chr6 994210 N DUP 10
SRR1766473.7978047 chr7 157324697 N chr7 157325009 N DEL 15
SRR1766442.13136366 chr7 157324697 N chr7 157325009 N DEL 10
SRR1766464.561889 chr7 157324385 N chr7 157325030 N DEL 12
SRR1766483.8244552 chr14 34735123 N chr14 34735250 N DEL 11
SRR1766453.10892011 chr14 34735123 N chr14 34735288 N DEL 11
SRR1766480.1702292 chr9 134524046 N chr9 134524175 N DUP 10
SRR1766479.7397739 chr9 134524128 N chr9 134524187 N DUP 10
SRR1766445.6411802 chr9 134523932 N chr9 134524191 N DUP 10
SRR1766466.6111114 chr6 522354 N chr6 522748 N DEL 15
SRR1766486.9232122 chr13 113375300 N chr13 113375981 N DEL 10
SRR1766442.16716254 chr13 113375340 N chr13 113376001 N DEL 10
SRR1766466.8833002 chr13 113375420 N chr13 113376001 N DEL 10
SRR1766453.1685489 chr13 113375367 N chr13 113375608 N DEL 10
SRR1766442.18034647 chr13 113375420 N chr13 113376001 N DEL 10
SRR1766483.1007781 chr13 113375420 N chr13 113376001 N DEL 10
SRR1766458.824786 chr13 113375289 N chr13 113375598 N DUP 16
SRR1766463.8563728 chr13 113375602 N chr13 113375921 N DUP 10
SRR1766442.7748246 chr13 113376001 N chr13 113376080 N DUP 15
SRR1766473.5647016 chr13 113376001 N chr13 113376080 N DUP 15
SRR1766446.8369414 chr13 113375580 N chr13 113376001 N DEL 10
SRR1766463.8786286 chr13 113375839 N chr13 113375998 N DUP 15
SRR1766458.824786 chr13 113375337 N chr13 113375958 N DEL 13
SRR1766452.381912 chr13 113376041 N chr13 113376349 N DEL 10
SRR1766460.5768967 chr6 71316412 N chr6 71316473 N DUP 10
SRR1766476.5189228 chr6 71316412 N chr6 71316473 N DUP 10
SRR1766483.1945455 chr18 3113373 N chr18 3113486 N DEL 15
SRR1766482.12819358 chr3 77323092 N chr3 77323144 N DUP 14
SRR1766470.5413413 chr3 77323092 N chr3 77323144 N DUP 10
SRR1766475.3383508 chr3 77323092 N chr3 77323231 N DUP 14
SRR1766460.8179183 chr3 77323072 N chr3 77323153 N DUP 10
SRR1766453.6593551 chr3 77323092 N chr3 77323144 N DUP 14
SRR1766478.4434323 chr3 77323092 N chr3 77323202 N DUP 10
SRR1766475.10073472 chr3 77323094 N chr3 77323146 N DUP 10
SRR1766480.1027218 chr3 77323092 N chr3 77323144 N DUP 12
SRR1766465.6317734 chr3 77323072 N chr3 77323211 N DUP 10
SRR1766464.7925165 chr3 77323092 N chr3 77323231 N DUP 12
SRR1766475.1021030 chr3 77323092 N chr3 77323144 N DUP 18
SRR1766459.1207565 chr3 77323068 N chr3 77323236 N DUP 12
SRR1766450.6971141 chr3 77323094 N chr3 77323204 N DUP 12
SRR1766475.7501766 chr3 77323068 N chr3 77323236 N DUP 13
SRR1766451.7845618 chrY 10790402 N chrY 10790643 N DEL 12
SRR1766452.2963636 chr2 38479868 N chr2 38480021 N DEL 11
SRR1766450.3678986 chr19 14636173 N chr19 14636299 N DEL 15
SRR1766453.9491509 chr19 14636175 N chr19 14636301 N DEL 13
SRR1766466.6225683 chr19 14636176 N chr19 14636302 N DEL 12
SRR1766442.21322860 chr19 14636177 N chr19 14636303 N DEL 11
SRR1766476.2570549 chr18 22740477 N chr18 22740571 N DUP 11
SRR1766461.3979564 chr18 22740477 N chr18 22740571 N DUP 12
SRR1766470.11076688 chr18 22740478 N chr18 22740572 N DUP 11
SRR1766479.7642685 chr18 22740480 N chr18 22740574 N DUP 13
SRR1766479.13293243 chr12 7197426 N chr12 7197528 N DUP 12
SRR1766444.4710132 chr12 7197426 N chr12 7197528 N DUP 12
SRR1766453.3652266 chr12 7197426 N chr12 7197528 N DUP 17
SRR1766478.5771996 chr12 7197490 N chr12 7197541 N DUP 10
SRR1766484.5798433 chr12 7197515 N chr12 7197588 N DUP 11
SRR1766475.7449761 chr12 7197454 N chr12 7197582 N DEL 11
SRR1766454.6180553 chr12 7197454 N chr12 7197582 N DEL 10
SRR1766449.8470532 chr12 7197454 N chr12 7197582 N DEL 10
SRR1766470.4351337 chr10 82098397 N chr10 82098473 N DEL 13
SRR1766449.1348248 chr10 82098400 N chr10 82098476 N DEL 12
SRR1766453.2639819 chr1 167806412 N chr1 167806490 N DEL 10
SRR1766473.4912186 chr1 167806409 N chr1 167806487 N DEL 10
SRR1766450.2462552 chrX 1581852 N chrX 1582057 N DUP 14
SRR1766471.3529461 chrX 1581677 N chrX 1582162 N DEL 10
SRR1766471.11551969 chrX 1581686 N chrX 1582373 N DEL 10
SRR1766456.6043241 chr6 166824827 N chr6 166824926 N DEL 14
SRR1766461.1932987 chr6 166824810 N chr6 166824903 N DEL 15
SRR1766468.2685443 chr6 166824860 N chr6 166824957 N DEL 11
SRR1766475.10985322 chr6 166824795 N chr6 166824860 N DUP 13
SRR1766469.44660 chr6 166824926 N chr6 166824989 N DUP 18
SRR1766479.5464903 chr6 166824776 N chr6 166824967 N DEL 12
SRR1766459.3169022 chr6 166824776 N chr6 166824967 N DEL 12
SRR1766485.7585292 chr7 61610125 N chr7 61610543 N DEL 13
SRR1766454.6379474 chr5 21344829 N chr5 21344912 N DEL 17
SRR1766453.551323 chr5 21344829 N chr5 21344912 N DEL 17
SRR1766449.3101329 chr5 21344829 N chr5 21344912 N DEL 17
SRR1766485.4826104 chr10 16646011 N chr10 16646070 N DUP 11
SRR1766477.3528578 chr10 16646011 N chr10 16646070 N DUP 12
SRR1766442.21891090 chr10 16646011 N chr10 16646070 N DUP 15
SRR1766447.10488370 chr10 16646011 N chr10 16646112 N DUP 11
SRR1766448.1342968 chr10 16646011 N chr10 16646112 N DUP 16
SRR1766464.1106556 chr10 16646073 N chr10 16646156 N DEL 13
SRR1766464.7789299 chr17 77885469 N chr17 77885665 N DEL 10
SRR1766468.495698 chr13 87990186 N chr13 87990243 N DEL 18
SRR1766479.9892609 chr13 87990186 N chr13 87990243 N DEL 15
SRR1766475.4352322 chr13 87990186 N chr13 87990243 N DEL 13
SRR1766449.3646662 chr13 87990186 N chr13 87990243 N DEL 13
SRR1766458.1705585 chr13 87990186 N chr13 87990243 N DEL 12
SRR1766442.10766529 chr3 197877336 N chr3 197877661 N DEL 10
SRR1766459.4277807 chr3 197877063 N chr3 197877712 N DEL 10
SRR1766470.6113389 chr8 142116253 N chr8 142116746 N DEL 15
SRR1766460.879122 chr8 142116186 N chr8 142116269 N DUP 10
SRR1766461.9765918 chr8 142116267 N chr8 142116736 N DEL 19
SRR1766474.5479588 chr8 142116194 N chr8 142116309 N DUP 13
SRR1766442.45343044 chr8 142116268 N chr8 142116345 N DEL 10
SRR1766442.23242165 chr8 142116109 N chr8 142116433 N DEL 13
SRR1766459.136911 chr8 142115961 N chr8 142116570 N DEL 10
SRR1766460.879122 chr8 142116628 N chr8 142116783 N DUP 18
SRR1766457.1348101 chr19 7640147 N chr19 7640632 N DEL 14
SRR1766461.9420238 chr19 7640206 N chr19 7640505 N DEL 11
SRR1766482.7113450 chr19 7640356 N chr19 7640645 N DUP 12
SRR1766471.11517789 chr19 7640290 N chr19 7640369 N DEL 10
SRR1766442.14653607 chr19 7640438 N chr19 7640687 N DUP 13
SRR1766463.1473794 chr19 7640335 N chr19 7640538 N DEL 18
SRR1766447.4780252 chr19 7640293 N chr19 7640542 N DEL 11
SRR1766483.7795068 chr19 7640600 N chr19 7640661 N DUP 10
SRR1766457.1348101 chr19 7640327 N chr19 7640618 N DEL 15
SRR1766446.2767360 chr19 7640291 N chr19 7640628 N DEL 11
SRR1766462.6250909 chr6 167575839 N chr6 167575987 N DEL 10
SRR1766446.588066 chr8 1698487 N chr8 1698631 N DUP 10
SRR1766477.10707876 chr8 1698652 N chr8 1699088 N DEL 15
SRR1766477.2277245 chr8 1698518 N chr8 1698664 N DEL 10
SRR1766484.93610 chr8 1698664 N chr8 1698808 N DUP 10
SRR1766478.6232040 chr8 1698752 N chr8 1698808 N DUP 10
SRR1766447.3412355 chr8 1698440 N chr8 1698788 N DEL 15
SRR1766459.8806486 chr8 1698808 N chr8 1698923 N DEL 15
SRR1766448.3198592 chr8 1698473 N chr8 1698935 N DEL 10
SRR1766457.1967128 chr8 1698561 N chr8 1699023 N DEL 15
SRR1766442.29334801 chr18 78755796 N chr18 78755972 N DUP 12
SRR1766471.2193416 chr18 78755792 N chr18 78755968 N DUP 10
SRR1766442.40012687 chr9 137861493 N chr9 137861710 N DEL 13
SRR1766442.742115 chrY 10773275 N chrY 10773371 N DEL 13
SRR1766464.2190590 chr8 79730478 N chr8 79730609 N DUP 10
SRR1766477.3911342 chr5 49687 N chr5 49778 N DEL 11
SRR1766481.4145111 chr5 49687 N chr5 49778 N DEL 11
SRR1766442.22613791 chr4 117740053 N chr4 117740136 N DEL 14
SRR1766455.4700077 chr4 117740055 N chr4 117740138 N DEL 12
SRR1766465.5813673 chr4 117740055 N chr4 117740138 N DEL 12
SRR1766477.1375051 chr4 117740054 N chr4 117740137 N DEL 13
SRR1766471.2358954 chr4 117740226 N chr4 117740320 N DEL 10
SRR1766442.10497564 chr4 117740226 N chr4 117740320 N DEL 11
SRR1766453.2545477 chr4 117740228 N chr4 117740322 N DEL 13
SRR1766465.762195 chr4 117740227 N chr4 117740321 N DEL 14
SRR1766465.211241 chr16 89342136 N chr16 89342227 N DEL 19
SRR1766462.8886384 chr16 89342136 N chr16 89342227 N DEL 18
SRR1766472.10773969 chrX 1297339 N chrX 1297452 N DUP 10
SRR1766476.10407791 chrX 1297415 N chrX 1297473 N DEL 10
SRR1766445.5498862 chrX 1297273 N chrX 1297443 N DUP 10
SRR1766443.1933880 chrX 1297340 N chrX 1297453 N DUP 10
SRR1766442.20723698 chrX 1297339 N chrX 1297452 N DUP 10
SRR1766470.10770788 chrX 1297409 N chrX 1297465 N DUP 10
SRR1766445.8876915 chrX 1297263 N chrX 1297547 N DUP 12
SRR1766474.4541691 chrX 1297473 N chrX 1297529 N DUP 10
SRR1766454.8963487 chrX 1297486 N chrX 1297542 N DUP 10
SRR1766463.3610676 chr3 60860390 N chr3 60860455 N DUP 11
SRR1766479.13600969 chr3 60860390 N chr3 60860455 N DUP 11
SRR1766472.3986952 chr3 60860390 N chr3 60860455 N DUP 11
SRR1766473.817752 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766454.2085433 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766444.1734587 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766448.7267246 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766460.10344168 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766477.10564264 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766465.5888777 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766483.7088928 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766448.9888280 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766444.1734587 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766473.9139992 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766479.13726865 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766452.6164498 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766471.697922 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766462.4032350 chr13 35124778 N chr13 35124915 N DEL 12
SRR1766467.11041177 chr13 35124778 N chr13 35124915 N DEL 12
SRR1766456.1892722 chr12 39713610 N chr12 39713759 N DUP 10
SRR1766465.2601458 chr8 123315143 N chr8 123315495 N DEL 19
SRR1766463.10957138 chr8 123315143 N chr8 123315495 N DEL 15
SRR1766461.9696750 chr8 123315298 N chr8 123315957 N DEL 10
SRR1766461.9696750 chr8 123315305 N chr8 123315757 N DUP 10
SRR1766485.4406859 chr8 123315190 N chr8 123315591 N DEL 13
SRR1766466.4885941 chr8 123315673 N chr8 123316106 N DUP 10
SRR1766480.1413409 chr8 123315203 N chr8 123315960 N DEL 10
SRR1766443.2470571 chr8 123315730 N chr8 123316060 N DUP 11
SRR1766442.23239024 chr7 157439769 N chr7 157439825 N DEL 12
SRR1766471.2054337 chr7 157439596 N chr7 157440124 N DEL 10
SRR1766454.618763 chrY 10976009 N chrY 10976111 N DEL 10
SRR1766455.6011185 chrY 10976009 N chrY 10976111 N DEL 10
SRR1766449.10556070 chrX 818457 N chrX 818546 N DEL 15
SRR1766472.7772488 chrX 818428 N chrX 818546 N DEL 15
SRR1766446.1074889 chrX 818457 N chrX 818546 N DEL 17
SRR1766475.976711 chr22 46609045 N chr22 46609164 N DEL 10
SRR1766455.4851743 chr8 139997414 N chr8 139997732 N DUP 10
SRR1766469.5150890 chr8 139997342 N chr8 139997640 N DEL 10
SRR1766445.3513444 chr19 57138016 N chr19 57138178 N DUP 14
SRR1766465.6743129 chr19 57138060 N chr19 57138116 N DUP 13
SRR1766475.7586315 chr19 57137986 N chr19 57138146 N DUP 12
SRR1766469.10762129 chr19 57138052 N chr19 57138155 N DUP 10
SRR1766474.60635 chr19 57138024 N chr19 57138099 N DUP 13
SRR1766463.3412795 chr19 57138057 N chr19 57138133 N DUP 12
SRR1766442.35089032 chr19 57138028 N chr19 57138152 N DUP 12
SRR1766442.38839232 chr19 57138011 N chr19 57138242 N DUP 14
SRR1766470.9249561 chr19 57138052 N chr19 57138231 N DUP 15
SRR1766472.2081827 chr22 42087844 N chr22 42088450 N DEL 10
SRR1766471.6319322 chr22 42087820 N chr22 42088424 N DUP 15
SRR1766443.2575371 chr22 42087670 N chr22 42087976 N DEL 13
SRR1766453.5082174 chr22 42087726 N chr22 42088332 N DEL 10
SRR1766475.405940 chr5 95360576 N chr5 95360665 N DUP 14
SRR1766479.12623699 chr9 20417278 N chr9 20417443 N DEL 10
SRR1766479.4174472 chrX 2166513 N chrX 2166576 N DEL 19
SRR1766473.6198366 chr9 119250198 N chr9 119250259 N DEL 12
SRR1766456.708743 chr5 15935502 N chr5 15935787 N DEL 11
SRR1766466.7598979 chr14 34350232 N chr14 34350323 N DEL 10
SRR1766469.9186669 chr14 34349958 N chr14 34350472 N DEL 10
SRR1766474.1345334 chr14 34350188 N chr14 34350247 N DUP 10
SRR1766484.11739419 chr14 34350188 N chr14 34350247 N DUP 10
SRR1766461.6617292 chr14 34350232 N chr14 34350293 N DEL 10
SRR1766466.6752984 chr4 2430240 N chr4 2430302 N DUP 10
SRR1766457.1214383 chr4 2430240 N chr4 2430302 N DUP 10
SRR1766462.3980863 chr4 2430240 N chr4 2430302 N DUP 10
SRR1766449.21631 chr4 2430230 N chr4 2430609 N DEL 10
SRR1766473.782496 chr4 2430337 N chr4 2430464 N DEL 10
SRR1766457.8278912 chr4 2430230 N chr4 2430672 N DEL 10
SRR1766444.679140 chr4 2430410 N chr4 2430726 N DEL 10
SRR1766480.1687803 chr5 160504972 N chr5 160505148 N DEL 11
SRR1766472.11821186 chr5 2219487 N chr5 2219537 N DUP 10
SRR1766476.732756 chr22 46194970 N chr22 46195300 N DEL 15
SRR1766478.10327167 chr12 39712315 N chr12 39712512 N DUP 13
SRR1766442.41243329 chr12 39712252 N chr12 39712513 N DUP 14
SRR1766444.3363549 chr10 7526771 N chr10 7526828 N DUP 11
SRR1766455.6347094 chr10 7526771 N chr10 7526828 N DUP 12
SRR1766467.10990244 chr10 7526850 N chr10 7526983 N DUP 16
SRR1766462.1802173 chr10 7526781 N chr10 7526923 N DUP 12
SRR1766486.2647662 chr10 7526782 N chr10 7526924 N DUP 11
SRR1766479.10906004 chr10 7526850 N chr10 7526983 N DUP 14
SRR1766468.5144228 chr16 34583291 N chr16 34583362 N DUP 11
SRR1766469.5829954 chr16 34583299 N chr16 34583393 N DUP 10
SRR1766451.4286354 chr9 80122819 N chr9 80123403 N DUP 13
SRR1766481.9801896 chr9 80122819 N chr9 80123403 N DUP 13
SRR1766477.8275190 chr14 79471048 N chr14 79471111 N DEL 15
SRR1766473.9396436 chr14 79471048 N chr14 79471111 N DEL 15
SRR1766481.8309394 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766478.9892453 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766469.8403513 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766484.11461911 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766471.7683050 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766471.10708940 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766447.10788821 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766458.4102203 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766461.9033213 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766468.2323489 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766465.10276724 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766442.30073744 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766476.7013938 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766451.10333380 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766442.42097907 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766445.3539154 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766467.4136555 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766475.3192630 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766449.7045159 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766457.7278639 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766467.1108090 chr22 38807715 N chr22 38807941 N DUP 10
SRR1766446.10531661 chr10 92393448 N chr10 92393539 N DEL 19
SRR1766459.1943428 chr10 92393448 N chr10 92393539 N DEL 19
SRR1766460.416714 chr10 92393448 N chr10 92393539 N DEL 17
SRR1766479.6574 chr10 108880281 N chr10 108880339 N DUP 15
SRR1766442.39887904 chr10 108880281 N chr10 108880339 N DUP 16
SRR1766463.6114574 chr14 101245352 N chr14 101245911 N DEL 10
SRR1766478.1825873 chr14 101245352 N chr14 101245911 N DEL 10
SRR1766465.9327965 chr14 101245352 N chr14 101245533 N DEL 15
SRR1766484.7439924 chr14 101245362 N chr14 101245435 N DEL 11
SRR1766452.2424098 chr14 101245344 N chr14 101245831 N DEL 14
SRR1766481.8432542 chr14 101245352 N chr14 101245911 N DEL 15
SRR1766478.9702500 chr14 101245344 N chr14 101245831 N DEL 15
SRR1766446.420543 chr14 101245345 N chr14 101245544 N DEL 10
SRR1766479.13375974 chr14 101245271 N chr14 101245324 N DUP 12
SRR1766443.5828807 chr14 101245271 N chr14 101245342 N DUP 16
SRR1766462.1978821 chr14 101245345 N chr14 101245904 N DEL 15
SRR1766466.4792661 chr14 101245370 N chr14 101245821 N DEL 15
SRR1766470.1638359 chr14 101245345 N chr14 101245578 N DUP 10
SRR1766470.5716333 chr14 101245298 N chr14 101245533 N DEL 19
SRR1766485.4283071 chr14 101245423 N chr14 101245944 N DUP 15
SRR1766474.3378948 chr14 101245273 N chr14 101245902 N DUP 15
SRR1766442.1229275 chr14 101245291 N chr14 101245902 N DUP 10
SRR1766470.1825605 chr14 101245273 N chr14 101245470 N DUP 14
SRR1766450.7194758 chr14 101245332 N chr14 101245423 N DEL 13
SRR1766449.8007059 chr14 101245892 N chr14 101246379 N DEL 15
SRR1766465.1116988 chr14 101245308 N chr14 101245435 N DEL 15
SRR1766484.2331466 chr14 101245281 N chr14 101245426 N DEL 14
SRR1766486.8858851 chr14 101245318 N chr14 101245515 N DUP 10
SRR1766446.2136184 chr14 101245290 N chr14 101245435 N DEL 13
SRR1766476.1774820 chr14 101245221 N chr14 101245438 N DEL 12
SRR1766442.30835632 chr14 101245536 N chr14 101246203 N DEL 15
SRR1766442.38613342 chr14 101245281 N chr14 101245532 N DUP 10
SRR1766466.8893021 chr14 101245303 N chr14 101246454 N DUP 13
SRR1766473.5689713 chr14 101245435 N chr14 101245542 N DUP 10
SRR1766460.8212328 chr14 101245496 N chr14 101245821 N DEL 14
SRR1766462.8603687 chr14 101245548 N chr14 101246215 N DEL 10
SRR1766479.13375974 chr14 101245453 N chr14 101245508 N DEL 10
SRR1766447.5452777 chr14 101245435 N chr14 101245614 N DUP 10
SRR1766458.6651298 chr14 101245271 N chr14 101245558 N DUP 15
SRR1766465.11064262 chr14 101245273 N chr14 101245578 N DUP 16
SRR1766454.2135611 chr14 101246005 N chr14 101246708 N DEL 15
SRR1766442.15262427 chr14 101245221 N chr14 101245528 N DEL 10
SRR1766442.42286057 chr14 101245452 N chr14 101245543 N DEL 10
SRR1766445.4212652 chr14 101245591 N chr14 101245896 N DUP 15
SRR1766470.2488826 chr14 101245597 N chr14 101245904 N DEL 13
SRR1766481.1297127 chr14 101245482 N chr14 101245591 N DEL 10
SRR1766478.2367219 chr14 101245623 N chr14 101246864 N DUP 15
SRR1766477.3098970 chr14 101245380 N chr14 101245451 N DUP 18
SRR1766442.5700407 chr14 101245533 N chr14 101245658 N DUP 15
SRR1766447.7848055 chr14 101245640 N chr14 101245821 N DEL 18
SRR1766472.6341740 chr14 101245314 N chr14 101245621 N DEL 15
SRR1766485.8047111 chr14 101245314 N chr14 101245621 N DEL 15
SRR1766451.3254329 chr14 101245633 N chr14 101245686 N DUP 10
SRR1766450.4364560 chr14 101245358 N chr14 101245431 N DEL 10
SRR1766463.5282942 chr14 101245623 N chr14 101245694 N DUP 15
SRR1766469.6404545 chr14 101245280 N chr14 101245623 N DEL 15
SRR1766442.36906202 chr14 101245633 N chr14 101245686 N DUP 15
SRR1766442.2944098 chr14 101245723 N chr14 101245904 N DEL 10
SRR1766452.2250233 chr14 101245274 N chr14 101245507 N DUP 15
SRR1766464.1808613 chr14 101245282 N chr14 101245713 N DUP 10
SRR1766471.10588742 chr14 101245307 N chr14 101246100 N DEL 15
SRR1766447.8209277 chr14 101245624 N chr14 101246829 N DUP 14
SRR1766442.21797007 chr14 101245282 N chr14 101245713 N DUP 10
SRR1766463.6114574 chr14 101245401 N chr14 101245726 N DEL 15
SRR1766486.6495742 chr14 101245706 N chr14 101245903 N DUP 10
SRR1766446.1672006 chr14 101245309 N chr14 101245812 N DUP 10
SRR1766454.7690490 chr14 101245281 N chr14 101245748 N DUP 15
SRR1766459.8727129 chr14 101245289 N chr14 101245792 N DUP 15
SRR1766464.8372563 chr14 101245352 N chr14 101245749 N DEL 10
SRR1766483.1597335 chr14 101245298 N chr14 101245749 N DEL 12
SRR1766454.2060420 chr14 101245767 N chr14 101245892 N DUP 14
SRR1766481.8432542 chr14 101245298 N chr14 101245749 N DEL 10
SRR1766446.6150418 chr14 101245298 N chr14 101246487 N DEL 15
SRR1766465.5700396 chr14 101245282 N chr14 101245785 N DUP 10
SRR1766446.6150418 chr14 101245829 N chr14 101246316 N DEL 10
SRR1766465.439369 chr14 101245317 N chr14 101245460 N DUP 10
SRR1766454.8144665 chr14 101245298 N chr14 101245821 N DEL 15
SRR1766447.5452777 chr14 101245294 N chr14 101245817 N DEL 10
SRR1766467.2066155 chr14 101245823 N chr14 101246830 N DUP 11
SRR1766477.2321932 chr14 101245346 N chr14 101245527 N DEL 17
SRR1766481.10341623 chr14 101245290 N chr14 101245831 N DEL 13
SRR1766466.4792661 chr14 101245352 N chr14 101246487 N DEL 19
SRR1766466.10752342 chr14 101245333 N chr14 101246324 N DEL 10
SRR1766459.5305497 chr14 101245821 N chr14 101246036 N DUP 10
SRR1766478.9074782 chr14 101245275 N chr14 101245886 N DUP 10
SRR1766463.10018286 chr14 101245271 N chr14 101245378 N DUP 18
SRR1766450.4428949 chr14 101245271 N chr14 101245378 N DUP 17
SRR1766453.6407873 chr14 101245274 N chr14 101245903 N DUP 10
SRR1766442.5693907 chr14 101245362 N chr14 101245453 N DEL 14
SRR1766473.5689713 chr14 101245271 N chr14 101245360 N DUP 10
SRR1766469.5260493 chr14 101245271 N chr14 101245378 N DUP 17
SRR1766462.2601057 chr14 101245279 N chr14 101245908 N DUP 10
SRR1766453.6407873 chr14 101245496 N chr14 101245911 N DEL 15
SRR1766479.6506790 chr14 101245278 N chr14 101245349 N DUP 15
SRR1766449.9274970 chr14 101245586 N chr14 101245911 N DEL 10
SRR1766486.1210980 chr14 101245370 N chr14 101245911 N DEL 15
SRR1766477.3098970 chr14 101245332 N chr14 101246089 N DEL 10
SRR1766454.7375551 chr14 101245271 N chr14 101245954 N DUP 10
SRR1766484.7439924 chr14 101245344 N chr14 101245939 N DEL 10
SRR1766450.7194758 chr14 101245425 N chr14 101245964 N DUP 15
SRR1766463.7734475 chr14 101245460 N chr14 101245911 N DEL 10
SRR1766466.3621639 chr14 101245974 N chr14 101246101 N DEL 10
SRR1766449.1277676 chr14 101245831 N chr14 101245992 N DUP 19
SRR1766486.11512295 chr14 101245821 N chr14 101246000 N DUP 16
SRR1766450.8037774 chr14 101245317 N chr14 101245442 N DUP 12
SRR1766470.10752330 chr14 101245308 N chr14 101245939 N DEL 10
SRR1766442.10000842 chr14 101245281 N chr14 101245948 N DEL 10
SRR1766483.4238392 chr14 101245974 N chr14 101246101 N DEL 10
SRR1766468.31014 chr14 101245271 N chr14 101245378 N DUP 15
SRR1766443.11096063 chr14 101245308 N chr14 101245453 N DEL 14
SRR1766450.3353896 chr14 101245913 N chr14 101246074 N DUP 10
SRR1766465.11064262 chr14 101245536 N chr14 101246707 N DEL 10
SRR1766443.6819343 chr14 101246087 N chr14 101246214 N DEL 15
SRR1766470.396866 chr14 101246076 N chr14 101246473 N DEL 10
SRR1766479.11943828 chr14 101245819 N chr14 101246088 N DUP 10
SRR1766455.5129217 chr14 101246163 N chr14 101246560 N DEL 10
SRR1766447.10219899 chr14 101245831 N chr14 101246136 N DUP 15
SRR1766484.761616 chr14 101245307 N chr14 101246100 N DEL 10
SRR1766468.5097685 chr14 101245325 N chr14 101246100 N DEL 10
SRR1766445.1207403 chr14 101245460 N chr14 101246379 N DEL 15
SRR1766486.11512295 chr14 101246100 N chr14 101246603 N DUP 15
SRR1766470.1895312 chr14 101245325 N chr14 101246100 N DEL 10
SRR1766445.7569450 chr14 101245442 N chr14 101246379 N DEL 10
SRR1766463.4513275 chr14 101245946 N chr14 101246379 N DEL 15
SRR1766442.33696470 chr14 101245289 N chr14 101246100 N DEL 13
SRR1766470.396866 chr14 101245442 N chr14 101246379 N DEL 10
SRR1766464.6546876 chr14 101245442 N chr14 101246379 N DEL 10
SRR1766484.2989722 chr14 101245271 N chr14 101245378 N DUP 15
SRR1766471.9908205 chr14 101245579 N chr14 101246174 N DEL 10
SRR1766442.42250094 chr14 101245368 N chr14 101246215 N DEL 10
SRR1766458.3178253 chr14 101245318 N chr14 101245515 N DUP 10
SRR1766453.6240820 chr14 101245587 N chr14 101246182 N DEL 15
SRR1766453.879915 chr14 101245694 N chr14 101246217 N DEL 15
SRR1766457.8017718 chr14 101245370 N chr14 101246217 N DEL 16
SRR1766449.6654833 chr14 101245296 N chr14 101246215 N DEL 10
SRR1766455.5129217 chr14 101245932 N chr14 101246473 N DEL 16
SRR1766468.2840145 chr14 101245904 N chr14 101246281 N DUP 15
SRR1766477.6709766 chr14 101245327 N chr14 101246298 N DUP 10
SRR1766461.3588899 chr14 101245334 N chr14 101246289 N DEL 10
SRR1766482.4872556 chr14 101245821 N chr14 101246306 N DUP 19
SRR1766449.5020930 chr14 101245334 N chr14 101245533 N DEL 10
SRR1766454.11030453 chr14 101245271 N chr14 101245468 N DUP 10
SRR1766454.7690490 chr14 101245314 N chr14 101246287 N DEL 10
SRR1766443.7847574 chr14 101245345 N chr14 101245452 N DUP 15
SRR1766484.5382012 chr14 101245300 N chr14 101246291 N DEL 10
SRR1766451.3254329 chr14 101245326 N chr14 101246317 N DEL 17
SRR1766475.8846686 chr14 101245344 N chr14 101246317 N DEL 19
SRR1766456.3516764 chr14 101245478 N chr14 101246379 N DEL 15
SRR1766457.6100005 chr14 101245496 N chr14 101246379 N DEL 10
SRR1766468.6715708 chr14 101245283 N chr14 101246452 N DUP 15
SRR1766471.7528543 chr14 101245290 N chr14 101246011 N DEL 10
SRR1766482.4872556 chr14 101245273 N chr14 101245902 N DUP 10
SRR1766464.2378079 chr14 101245889 N chr14 101246178 N DEL 10
SRR1766473.6728132 chr14 101245452 N chr14 101246425 N DEL 10
SRR1766479.5642890 chr14 101245579 N chr14 101246444 N DEL 10
SRR1766479.9225617 chr14 101245453 N chr14 101246444 N DEL 10
SRR1766442.42250094 chr14 101245692 N chr14 101246485 N DEL 15
SRR1766481.11495774 chr14 101245314 N chr14 101246485 N DEL 12
SRR1766486.4776314 chr14 101245921 N chr14 101246550 N DUP 10
SRR1766465.4071350 chr14 101245309 N chr14 101246550 N DUP 15
SRR1766479.11943828 chr14 101245676 N chr14 101246487 N DEL 10
SRR1766444.5740043 chr14 101245328 N chr14 101246551 N DUP 15
SRR1766459.2447632 chr14 101245320 N chr14 101246473 N DEL 10
SRR1766442.33647476 chr14 101245296 N chr14 101246485 N DEL 10
SRR1766442.36720550 chr14 101246281 N chr14 101246552 N DEL 15
SRR1766469.9614842 chr14 101246295 N chr14 101246546 N DUP 10
SRR1766480.6181736 chr14 101246299 N chr14 101246552 N DEL 10
SRR1766461.7594490 chr14 101245865 N chr14 101246604 N DEL 10
SRR1766477.6589584 chr14 101246570 N chr14 101246623 N DUP 16
SRR1766442.466758 chr14 101245471 N chr14 101246552 N DEL 10
SRR1766442.31600668 chr14 101245481 N chr14 101246580 N DEL 15
SRR1766481.9721316 chr14 101245865 N chr14 101246604 N DEL 10
SRR1766459.424307 chr14 101245691 N chr14 101246610 N DEL 11
SRR1766444.5740043 chr14 101245973 N chr14 101246604 N DEL 14
SRR1766485.11852955 chr14 101245291 N chr14 101246570 N DEL 13
SRR1766479.6506790 chr14 101245865 N chr14 101246604 N DEL 10
SRR1766463.3487261 chr14 101245865 N chr14 101246604 N DEL 10
SRR1766457.7217813 chr14 101245361 N chr14 101246604 N DEL 13
SRR1766456.1886143 chr14 101245273 N chr14 101246676 N DUP 15
SRR1766483.7188093 chr14 101246100 N chr14 101246603 N DUP 15
SRR1766452.6714314 chr14 101245533 N chr14 101246342 N DUP 10
SRR1766447.10219899 chr14 101245219 N chr14 101246642 N DEL 10
SRR1766484.7193371 chr14 101245920 N chr14 101246695 N DEL 10
SRR1766469.5943272 chr14 101245758 N chr14 101246731 N DEL 10
SRR1766464.937969 chr14 101245632 N chr14 101246497 N DEL 15
SRR1766479.11989098 chr14 101245460 N chr14 101245749 N DEL 12
SRR1766484.962215 chr14 101245921 N chr14 101246802 N DUP 10
SRR1766472.1116421 chr14 105570216 N chr14 105570792 N DEL 10
SRR1766457.9137224 chr14 105570133 N chr14 105570729 N DEL 10
SRR1766464.7136723 chr4 186043601 N chr4 186043666 N DUP 15
SRR1766475.7816568 chr4 186043304 N chr4 186043437 N DEL 10
SRR1766467.5874479 chr4 186043437 N chr4 186043700 N DUP 10
SRR1766463.3158830 chr4 186043518 N chr4 186043651 N DEL 10
SRR1766455.9305778 chr4 186043260 N chr4 186043523 N DUP 10
SRR1766462.6306000 chr4 186043259 N chr4 186043524 N DEL 10
SRR1766480.8697591 chr4 186043386 N chr4 186043585 N DEL 10
SRR1766464.10779901 chr4 186043383 N chr4 186043714 N DEL 10
SRR1766450.2393247 chr4 186043679 N chr4 186043746 N DEL 15
SRR1766486.8748168 chr2 60467221 N chr2 60467274 N DUP 11
SRR1766443.7941489 chr2 60467221 N chr2 60467337 N DUP 15
SRR1766471.5731134 chr2 60468151 N chr2 60468228 N DUP 13
SRR1766486.91312 chr2 60467296 N chr2 60467598 N DUP 12
SRR1766480.8030291 chr2 60467281 N chr2 60467583 N DUP 15
SRR1766471.1687300 chr2 60467307 N chr2 60467588 N DUP 16
SRR1766445.3464120 chr2 60467296 N chr2 60467598 N DUP 12
SRR1766446.4705664 chr2 60467408 N chr2 60467617 N DUP 16
SRR1766460.11092820 chr2 60467402 N chr2 60467605 N DUP 17
SRR1766465.2042980 chr2 60467297 N chr2 60467755 N DUP 18
SRR1766478.11860608 chr2 60467311 N chr2 60467744 N DEL 10
SRR1766450.4600800 chr2 60467335 N chr2 60467765 N DEL 12
SRR1766445.7527810 chr2 60467353 N chr2 60467825 N DEL 15
SRR1766464.5980845 chr2 60467297 N chr2 60467920 N DUP 19
SRR1766461.4846002 chr2 60467242 N chr2 60467879 N DEL 17
SRR1766481.10885226 chr2 60467555 N chr2 60467874 N DEL 10
SRR1766459.7325521 chr2 60467275 N chr2 60467816 N DEL 15
SRR1766483.5691955 chr2 60467286 N chr2 60468019 N DEL 10
SRR1766452.7151758 chr2 60467332 N chr2 60468056 N DEL 18
SRR1766478.8676184 chr2 60467221 N chr2 60468156 N DUP 16
SRR1766459.890083 chr2 60467244 N chr2 60468199 N DEL 10
SRR1766442.30954513 chr2 60467242 N chr2 60468227 N DEL 14
SRR1766443.7941489 chr2 60467314 N chr2 60468227 N DEL 10
SRR1766450.4837751 chr2 60467314 N chr2 60468272 N DEL 15
SRR1766482.10514975 chr2 60468190 N chr2 60468242 N DEL 13
SRR1766465.7484885 chr2 60468192 N chr2 60468262 N DEL 15
SRR1766485.3801890 chr2 60467256 N chr2 60468262 N DEL 10
SRR1766459.4304213 chr2 60467331 N chr2 60468271 N DEL 16
SRR1766443.871209 chr2 60467306 N chr2 60468261 N DEL 15
SRR1766484.770940 chr2 60467244 N chr2 60468271 N DEL 18
SRR1766455.3902386 chr2 60467241 N chr2 60468271 N DEL 15
SRR1766467.899119 chr2 60467313 N chr2 60468271 N DEL 15
SRR1766484.10722202 chr2 60467241 N chr2 60468271 N DEL 15
SRR1766461.4443736 chr2 60467268 N chr2 60468271 N DEL 10
SRR1766478.1923593 chr9 129339964 N chr9 129340017 N DEL 10
SRR1766457.1002041 chr17 402226 N chr17 402302 N DUP 12
SRR1766444.2198687 chr17 402226 N chr17 402302 N DUP 10
SRR1766477.1418828 chr17 402226 N chr17 402302 N DUP 12
SRR1766455.8706326 chr17 402226 N chr17 402302 N DUP 13
SRR1766480.219519 chr5 117993527 N chr5 117993580 N DEL 12
SRR1766446.1599666 chr5 117993527 N chr5 117993580 N DEL 13
SRR1766448.3767833 chr12 120021332 N chr12 120021636 N DEL 18
SRR1766447.5736528 chr12 120021396 N chr12 120021698 N DUP 10
SRR1766461.520360 chr12 120021719 N chr12 120022038 N DEL 19
SRR1766442.4211080 chr22 26736381 N chr22 26736598 N DEL 15
SRR1766449.7094048 chr1 83013731 N chr1 83013787 N DEL 10
SRR1766445.8204391 chr1 83013731 N chr1 83013787 N DEL 11
SRR1766461.2771859 chr1 83013731 N chr1 83013787 N DEL 17
SRR1766476.3864456 chr1 83013731 N chr1 83013787 N DEL 19
SRR1766479.8992341 chr1 83013731 N chr1 83013787 N DEL 16
SRR1766470.2374739 chr1 83013736 N chr1 83013787 N DEL 10
SRR1766446.372013 chr1 83013731 N chr1 83013787 N DEL 10
SRR1766453.9248675 chr1 83013731 N chr1 83013787 N DEL 10
SRR1766443.4637349 chr1 83013726 N chr1 83013787 N DEL 10
SRR1766485.11030020 chr1 83013698 N chr1 83013789 N DEL 15
SRR1766459.10635134 chr1 83013696 N chr1 83013787 N DEL 10
SRR1766469.8401615 chr1 83013698 N chr1 83013789 N DEL 15
SRR1766445.4701610 chr1 83013699 N chr1 83013790 N DEL 14
SRR1766443.8533574 chr1 83013700 N chr1 83013791 N DEL 13
SRR1766459.365250 chr1 83013702 N chr1 83013793 N DEL 11
SRR1766472.6607448 chr21 8594954 N chr21 8595147 N DEL 11
SRR1766466.7092978 chr3 180459351 N chr3 180459494 N DEL 14
SRR1766442.22467875 chr19 40648154 N chr19 40648409 N DEL 10
SRR1766469.1686096 chr19 40648188 N chr19 40648394 N DEL 10
SRR1766459.4715714 chr19 40648404 N chr19 40648454 N DUP 14
SRR1766451.3828811 chr19 40648404 N chr19 40648453 N DUP 16
SRR1766444.439063 chr12 122164137 N chr12 122164432 N DEL 10
SRR1766465.11018805 chr12 122164148 N chr12 122164746 N DEL 15
SRR1766486.3963338 chr9 9845197 N chr9 9845270 N DEL 12
SRR1766483.9943874 chr9 9845197 N chr9 9845270 N DEL 16
SRR1766476.8604135 chr9 9845211 N chr9 9845282 N DUP 17
SRR1766444.4430820 chr19 2973963 N chr19 2974261 N DEL 15
SRR1766442.44837182 chr19 2974059 N chr19 2974357 N DEL 10
SRR1766457.6197943 chr6 78554080 N chr6 78554135 N DEL 15
SRR1766470.5203252 chr6 78554078 N chr6 78554200 N DEL 10
SRR1766483.11966298 chr6 78554078 N chr6 78554200 N DEL 10
SRR1766479.9531288 chr12 14179718 N chr12 14179847 N DEL 11
SRR1766484.17580 chr12 14179718 N chr12 14179847 N DEL 13
SRR1766457.5758255 chr12 14179718 N chr12 14179847 N DEL 13
SRR1766471.11701813 chr12 14179718 N chr12 14179847 N DEL 16
SRR1766446.5787655 chr12 14179718 N chr12 14179927 N DEL 17
SRR1766481.11031130 chr12 14179718 N chr12 14179927 N DEL 17
SRR1766475.5335324 chr12 14179718 N chr12 14179927 N DEL 17
SRR1766442.36783829 chr12 14179755 N chr12 14179873 N DUP 10
SRR1766460.9014412 chr7 67850050 N chr7 67850103 N DEL 10
SRR1766454.6465392 chr6 82306852 N chr6 82306941 N DUP 11
SRR1766454.3230512 chr6 82306920 N chr6 82306999 N DEL 12
SRR1766458.6858572 chr6 82306996 N chr6 82307055 N DEL 17
SRR1766478.11040264 chr6 82306996 N chr6 82307055 N DEL 17
SRR1766450.10261164 chr6 82306998 N chr6 82307077 N DEL 16
SRR1766460.3745333 chr6 82306998 N chr6 82307077 N DEL 15
SRR1766458.3474171 chr6 82306998 N chr6 82307077 N DEL 15
SRR1766486.6220893 chr6 82306998 N chr6 82307077 N DEL 15
SRR1766463.5288650 chr6 82306998 N chr6 82307077 N DEL 15
SRR1766442.80768 chr12 131327113 N chr12 131327181 N DEL 12
SRR1766464.9519003 chr12 131327322 N chr12 131327392 N DUP 10
SRR1766476.7566276 chr12 131327117 N chr12 131327347 N DEL 13
SRR1766479.7246577 chr12 131327115 N chr12 131327345 N DEL 11
SRR1766481.10731177 chr13 106570720 N chr13 106570783 N DUP 12
SRR1766486.1896406 chr12 132518400 N chr12 132519012 N DEL 16
SRR1766476.9916818 chr12 132518635 N chr12 132518727 N DEL 15
SRR1766462.730940 chr12 132518680 N chr12 132518803 N DUP 10
SRR1766482.8161618 chr12 132518966 N chr12 132519110 N DEL 10
SRR1766467.10119278 chr2 236491181 N chr2 236491278 N DUP 10
SRR1766484.159036 chr2 236491181 N chr2 236491278 N DUP 11
SRR1766463.1122541 chr2 236491181 N chr2 236491278 N DUP 15
SRR1766469.5767519 chr2 236491181 N chr2 236491278 N DUP 15
SRR1766464.2476334 chrX 98534232 N chrX 98534439 N DUP 11
SRR1766453.8252410 chrX 98534236 N chrX 98534439 N DUP 16
SRR1766442.10833203 chr8 55767151 N chr8 55767254 N DEL 10
SRR1766485.10372490 chr8 55767153 N chr8 55767256 N DEL 13
SRR1766458.7750060 chr9 135261540 N chr9 135261799 N DUP 10
SRR1766457.3518584 chr9 135261530 N chr9 135261799 N DUP 16
SRR1766484.810925 chr9 135261535 N chr9 135261724 N DEL 12
SRR1766474.6905791 chr9 135261557 N chr9 135261726 N DEL 13
SRR1766457.1617167 chr9 135261730 N chr9 135261805 N DUP 13
SRR1766455.2612109 chr9 135261730 N chr9 135261805 N DUP 13
SRR1766482.2305095 chr9 135261785 N chr9 135261944 N DUP 10
SRR1766455.8088660 chr9 135261474 N chr9 135261805 N DEL 10
SRR1766442.11925313 chr8 142674091 N chr8 142674285 N DEL 15
SRR1766458.9032698 chr3 15163738 N chr3 15163893 N DUP 10
SRR1766442.46811603 chr7 36939434 N chr7 36939517 N DEL 15
SRR1766455.2933259 chr7 36939434 N chr7 36939517 N DEL 15
SRR1766446.2478883 chr7 36939434 N chr7 36939517 N DEL 15
SRR1766477.4994065 chr7 36939434 N chr7 36939517 N DEL 15
SRR1766450.5949375 chr7 36939437 N chr7 36939520 N DEL 12
SRR1766462.2569474 chr22 23381270 N chr22 23381411 N DEL 15
SRR1766445.8498237 chr22 23381269 N chr22 23381413 N DEL 12
SRR1766485.7849889 chr1 1056492 N chr1 1056581 N DEL 11
SRR1766454.2754508 chr10 41755895 N chr10 41756753 N DEL 17
SRR1766476.8508302 chr10 41755533 N chr10 41756390 N DEL 10
SRR1766442.42184993 chr7 14471315 N chr7 14471407 N DEL 13
SRR1766449.7626711 chr7 14471405 N chr7 14471530 N DUP 13
SRR1766469.4150726 chr7 14471405 N chr7 14471530 N DUP 14
SRR1766481.12693527 chr7 14471405 N chr7 14471530 N DUP 14
SRR1766442.15588503 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766442.37713788 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766449.1240833 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766464.10588109 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766442.40180803 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766483.78704 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766448.7831943 chr7 14471405 N chr7 14471530 N DUP 11
SRR1766454.5217581 chr7 14471405 N chr7 14471530 N DUP 11
SRR1766468.2715767 chr7 14471405 N chr7 14471530 N DUP 11
SRR1766455.8519310 chr7 14471405 N chr7 14471530 N DUP 10
SRR1766442.9179734 chr7 14471405 N chr7 14471530 N DUP 10
SRR1766449.7626711 chr7 14471405 N chr7 14471530 N DUP 10
SRR1766482.2760425 chr7 14471405 N chr7 14471530 N DUP 10
SRR1766449.7449003 chr7 14471405 N chr7 14471466 N DUP 18
SRR1766467.11600466 chr7 14471405 N chr7 14471466 N DUP 18
SRR1766446.4336791 chr7 14471405 N chr7 14471466 N DUP 18
SRR1766486.11271527 chr7 14471405 N chr7 14471466 N DUP 18
SRR1766465.6965993 chr7 14471405 N chr7 14471466 N DUP 17
SRR1766442.4927756 chr7 14471405 N chr7 14471466 N DUP 17
SRR1766443.211294 chr7 14471405 N chr7 14471466 N DUP 17
SRR1766442.233973 chr7 14471405 N chr7 14471466 N DUP 19
SRR1766450.5102090 chr7 14471405 N chr7 14471466 N DUP 19
SRR1766478.1819822 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766445.7708660 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766446.3770641 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766471.5303173 chr7 14471405 N chr7 14471466 N DUP 19
SRR1766471.7149905 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766477.9785768 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766442.44498754 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766450.1169239 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766447.8222869 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766448.9387396 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766442.2648806 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766462.5752283 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766479.9203479 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766442.12253223 chr7 14471409 N chr7 14471470 N DUP 10
SRR1766442.33750572 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766471.8974421 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766481.10609624 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766453.1051164 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766471.3005635 chr7 14471405 N chr7 14471530 N DUP 13
SRR1766472.4514954 chr7 14471405 N chr7 14471530 N DUP 13
SRR1766472.389000 chr7 14471405 N chr7 14471530 N DUP 11
SRR1766478.5212267 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766457.6265077 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766471.7205843 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766457.6265077 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766470.9529769 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766466.37817 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766442.25108929 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766443.6083702 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766458.7578535 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766482.10852768 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766442.6585063 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766456.2489751 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766451.9708365 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766445.2585395 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766480.566338 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766459.1216777 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766475.2836113 chr7 14471405 N chr7 14471466 N DUP 15
SRR1766444.1066160 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766464.709269 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766447.8222869 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766474.3356550 chr7 14471405 N chr7 14471466 N DUP 17
SRR1766456.3903884 chr17 72948351 N chr17 72948460 N DEL 10
SRR1766477.10058285 chr17 72948351 N chr17 72948460 N DEL 10
SRR1766445.6756708 chr17 72948430 N chr17 72948501 N DUP 15
SRR1766448.5056434 chr17 72948430 N chr17 72948501 N DUP 15
SRR1766455.6281613 chr17 72948430 N chr17 72948501 N DUP 15
SRR1766454.7345606 chr17 72948360 N chr17 72948433 N DEL 10
SRR1766481.4109840 chr17 72948357 N chr17 72948430 N DEL 10
SRR1766481.1686056 chr17 72948447 N chr17 72948554 N DUP 16
SRR1766452.3967246 chr21 6573044 N chr21 6573208 N DUP 12
SRR1766455.7714545 chr17 891874 N chr17 892059 N DEL 15
SRR1766472.6656346 chr17 891869 N chr17 892347 N DEL 10
SRR1766444.259232 chr17 891857 N chr17 892298 N DUP 10
SRR1766446.8638380 chr17 891857 N chr17 892298 N DUP 17
SRR1766466.10502257 chr17 891904 N chr17 892234 N DUP 15
SRR1766469.2128702 chr17 891913 N chr17 892245 N DEL 14
SRR1766479.2204105 chr17 891911 N chr17 892243 N DEL 13
SRR1766456.2639566 chr17 891911 N chr17 892169 N DEL 12
SRR1766465.506976 chr17 891911 N chr17 892169 N DEL 12
SRR1766467.2065900 chr17 891911 N chr17 892169 N DEL 12
SRR1766450.2402753 chr17 891904 N chr17 892308 N DUP 10
SRR1766459.11362980 chr17 891904 N chr17 892308 N DUP 10
SRR1766464.4980319 chr17 892044 N chr17 892301 N DUP 10
SRR1766481.1777112 chr17 891904 N chr17 892087 N DUP 10
SRR1766454.1479710 chr17 892000 N chr17 892146 N DUP 10
SRR1766472.6656346 chr17 892022 N chr17 892388 N DUP 10
SRR1766469.9795142 chr17 891889 N chr17 892037 N DEL 14
SRR1766457.1900164 chr17 891889 N chr17 892037 N DEL 10
SRR1766453.1936841 chr17 892059 N chr17 892279 N DUP 10
SRR1766471.4387627 chr17 892059 N chr17 892279 N DUP 10
SRR1766451.6151269 chr17 891904 N chr17 892234 N DUP 19
SRR1766457.1900164 chr17 891857 N chr17 892407 N DUP 12
SRR1766451.6151269 chr17 891913 N chr17 892171 N DEL 16
SRR1766453.10977745 chr17 892169 N chr17 892279 N DUP 10
SRR1766442.25512711 chr17 891911 N chr17 892169 N DEL 10
SRR1766461.1441231 chr17 891913 N chr17 892171 N DEL 14
SRR1766464.7682659 chr17 891913 N chr17 892171 N DEL 10
SRR1766470.447434 chr17 891904 N chr17 892234 N DUP 15
SRR1766471.2982393 chr17 891893 N chr17 892188 N DEL 10
SRR1766476.4130494 chr17 892169 N chr17 892279 N DUP 10
SRR1766449.2820829 chr17 891913 N chr17 892208 N DEL 17
SRR1766476.3253926 chr17 892169 N chr17 892279 N DUP 12
SRR1766448.10068846 chr17 892169 N chr17 892279 N DUP 10
SRR1766456.1177652 chr17 891857 N chr17 892407 N DUP 10
SRR1766485.7399758 chr17 891899 N chr17 892266 N DUP 12
SRR1766449.10754332 chr17 891845 N chr17 892395 N DUP 18
SRR1766475.2602459 chr17 891857 N chr17 892298 N DUP 15
SRR1766474.643074 chr17 891913 N chr17 892171 N DEL 17
SRR1766458.6587337 chr17 891893 N chr17 892188 N DEL 10
SRR1766454.8643206 chr1 1099547 N chr1 1099933 N DEL 15
SRR1766442.41952013 chr1 1099543 N chr1 1099698 N DEL 15
SRR1766481.557565 chr1 1099217 N chr1 1099827 N DEL 10
SRR1766479.1068764 chr22 11019451 N chr22 11019720 N DEL 10
SRR1766466.7557129 chr22 11019501 N chr22 11019815 N DEL 10
SRR1766486.1121972 chr10 60240259 N chr10 60240368 N DEL 13
SRR1766477.8986785 chr10 60240259 N chr10 60240368 N DEL 13
SRR1766451.10459403 chr10 60240271 N chr10 60240402 N DUP 13
SRR1766474.7729092 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766442.20425156 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766467.6718301 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766466.3883400 chr10 60240205 N chr10 60240303 N DEL 14
SRR1766482.7427773 chr10 60240205 N chr10 60240303 N DEL 13
SRR1766463.3848720 chr6 84395673 N chr6 84395751 N DUP 14
SRR1766474.8263643 chr6 84395673 N chr6 84395755 N DUP 16
SRR1766470.2023851 chr6 84395673 N chr6 84395755 N DUP 18
SRR1766445.3886393 chr6 84395676 N chr6 84395762 N DUP 16
SRR1766451.9177715 chr6 84395676 N chr6 84395762 N DUP 17
SRR1766469.151355 chr6 84395673 N chr6 84395763 N DUP 19
SRR1766483.9951045 chr9 134977404 N chr9 134977461 N DEL 14
SRR1766482.5753684 chr9 134977404 N chr9 134977461 N DEL 14
SRR1766442.27305789 chr9 134977404 N chr9 134977461 N DEL 14
SRR1766442.8032591 chr9 134977404 N chr9 134977461 N DEL 15
SRR1766467.1904545 chr9 134977404 N chr9 134977461 N DEL 15
SRR1766459.3045532 chr9 134977404 N chr9 134977461 N DEL 10
SRR1766476.4309473 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766442.38469052 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766484.3894179 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766456.4700733 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766472.3604016 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766477.10974077 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766442.43984930 chr9 134977411 N chr9 134977646 N DUP 14
SRR1766454.10726972 chr9 134977433 N chr9 134977492 N DUP 19
SRR1766450.9781022 chr9 134977469 N chr9 134977596 N DUP 12
SRR1766476.10816124 chr9 134977469 N chr9 134977596 N DUP 12
SRR1766467.4816567 chr9 134977469 N chr9 134977596 N DUP 11
SRR1766479.4540809 chr9 134977469 N chr9 134977596 N DUP 10
SRR1766456.3413997 chr9 134977405 N chr9 134977530 N DUP 13
SRR1766449.419393 chr9 134977411 N chr9 134977506 N DUP 12
SRR1766475.9121539 chr9 134977411 N chr9 134977506 N DUP 11
SRR1766461.3935249 chr9 134977463 N chr9 134977518 N DUP 12
SRR1766473.1244817 chr9 134977421 N chr9 134977492 N DUP 15
SRR1766477.11513909 chr9 134977421 N chr9 134977492 N DUP 15
SRR1766481.106377 chr9 134977523 N chr9 134977614 N DUP 10
SRR1766458.7090655 chr9 134977523 N chr9 134977614 N DUP 11
SRR1766442.9244279 chr9 134977523 N chr9 134977612 N DUP 14
SRR1766476.8526366 chr9 134977523 N chr9 134977614 N DUP 12
SRR1766471.1607677 chr9 134977523 N chr9 134977614 N DUP 12
SRR1766454.9679075 chr9 134977523 N chr9 134977614 N DUP 13
SRR1766450.6772662 chr9 134977523 N chr9 134977614 N DUP 16
SRR1766452.464242 chr9 134977411 N chr9 134977626 N DEL 12
SRR1766473.5794568 chrX 2426503 N chrX 2426597 N DUP 10
SRR1766451.6830745 chr8 58301684 N chr8 58301733 N DUP 16
SRR1766443.10652901 chr8 58301684 N chr8 58301733 N DUP 19
SRR1766479.626894 chr7 77509939 N chr7 77510115 N DUP 12
SRR1766461.10855440 chr7 77509939 N chr7 77510117 N DUP 16
SRR1766445.4718043 chr7 77509939 N chr7 77510115 N DUP 12
SRR1766476.7955973 chr7 77509939 N chr7 77510115 N DUP 12
SRR1766466.11084121 chr7 77509939 N chr7 77510115 N DUP 12
SRR1766467.1787340 chr7 77509763 N chr7 77509939 N DEL 12
SRR1766446.5200636 chr7 77509773 N chr7 77509948 N DUP 10
SRR1766467.7868723 chr20 61444434 N chr20 61444579 N DUP 15
SRR1766447.1403723 chr20 61444434 N chr20 61444579 N DUP 16
SRR1766442.37515660 chr20 61444633 N chr20 61444716 N DUP 12
SRR1766444.1083896 chr20 61444666 N chr20 61444795 N DUP 18
SRR1766456.5230040 chr12 87486322 N chr12 87486497 N DEL 14
SRR1766484.7758897 chr12 87486595 N chr12 87486699 N DUP 12
SRR1766483.1172379 chr12 87486595 N chr12 87486699 N DUP 14
SRR1766459.11229876 chr12 87486595 N chr12 87486699 N DUP 14
SRR1766462.667741 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766452.9972041 chr5 59200701 N chr5 59200790 N DUP 10
SRR1766443.7152936 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766486.4593672 chr5 59200701 N chr5 59200790 N DUP 10
SRR1766461.8382651 chr5 59200701 N chr5 59200790 N DUP 10
SRR1766480.6926333 chr5 59200701 N chr5 59200790 N DUP 15
SRR1766463.4737383 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766447.5231820 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766482.11326733 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766451.2589525 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766448.7759843 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766480.546699 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766450.1008389 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766477.6197748 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766463.6770281 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766477.9405509 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766469.9516957 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766481.9091587 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766485.5767850 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766474.9484491 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766477.9111117 chr5 59200697 N chr5 59200820 N DEL 17
SRR1766480.4686596 chr5 59200697 N chr5 59200820 N DEL 17
SRR1766466.6670269 chr5 59200697 N chr5 59200820 N DEL 16
SRR1766448.4408527 chr15 78040755 N chr15 78041014 N DEL 14
SRR1766472.1655674 chr15 78040755 N chr15 78041014 N DEL 14
SRR1766485.3376636 chr15 78040755 N chr15 78041014 N DEL 14
SRR1766455.4618863 chr15 78040778 N chr15 78041043 N DUP 10
SRR1766485.1411607 chr15 78040842 N chr15 78041040 N DEL 10
SRR1766447.1311927 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766449.8249127 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766445.9434634 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766473.2895805 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766475.8405594 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766484.353820 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766473.7372831 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766476.9797489 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766463.1748149 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766464.6431826 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766465.5629767 chr10 54332447 N chr10 54332518 N DUP 18
SRR1766474.206051 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766485.3998464 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766451.4784982 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766458.7801432 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766461.8011289 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766484.2908288 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766473.10376766 chr10 54332415 N chr10 54332481 N DUP 12
SRR1766462.7049217 chr10 54332395 N chr10 54332502 N DUP 17
SRR1766446.5320884 chr10 54332395 N chr10 54332502 N DUP 17
SRR1766476.9049963 chr10 54332415 N chr10 54332517 N DUP 12
SRR1766486.9902244 chr10 54332415 N chr10 54332481 N DUP 17
SRR1766445.2751006 chr10 54332395 N chr10 54332502 N DUP 10
SRR1766451.8621775 chr10 54332430 N chr10 54332508 N DEL 10
SRR1766470.5371781 chr10 54332420 N chr10 54332498 N DEL 10
SRR1766445.5636215 chr10 54332420 N chr10 54332498 N DEL 10
SRR1766456.961921 chr10 54332420 N chr10 54332498 N DEL 10
SRR1766452.10728406 chr10 54332425 N chr10 54332503 N DEL 10
SRR1766466.5574371 chr10 54332425 N chr10 54332503 N DEL 10
SRR1766463.5292752 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766442.24575392 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766472.4590897 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766446.1722364 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766483.3084668 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766470.7666158 chr7 29645401 N chr7 29645499 N DUP 15
SRR1766465.9718384 chr7 29645402 N chr7 29645500 N DUP 14
SRR1766451.4509251 chr7 29645400 N chr7 29645496 N DUP 15
SRR1766484.11721869 chr7 29645400 N chr7 29645496 N DUP 15
SRR1766484.8909243 chr7 29645344 N chr7 29645409 N DEL 13
SRR1766449.1479476 chr7 29645344 N chr7 29645409 N DEL 11
SRR1766484.3072567 chr6 170114198 N chr6 170114301 N DUP 13
SRR1766459.3894899 chr6 170114189 N chr6 170114322 N DUP 12
SRR1766483.4372668 chr6 170114190 N chr6 170114323 N DUP 15
SRR1766453.1733493 chr15 101764259 N chr15 101764693 N DUP 10
SRR1766455.4302704 chr15 101764319 N chr15 101764411 N DEL 10
SRR1766482.12207217 chr15 101764166 N chr15 101764347 N DUP 10
SRR1766467.7537170 chr15 101764198 N chr15 101764634 N DEL 10
SRR1766455.8309116 chr2 240813036 N chr2 240813168 N DUP 17
SRR1766450.8103163 chr2 240813025 N chr2 240813176 N DUP 17
SRR1766467.426328 chr2 240813034 N chr2 240813185 N DUP 15
SRR1766442.17802355 chr2 240812914 N chr2 240813025 N DEL 15
SRR1766445.5308104 chr2 240813034 N chr2 240813109 N DUP 12
SRR1766469.4241378 chr2 240813029 N chr2 240813104 N DUP 10
SRR1766444.3285386 chr2 240812821 N chr2 240813123 N DUP 11
SRR1766478.1226564 chr2 240813034 N chr2 240813109 N DUP 12
SRR1766442.6040113 chr2 240813025 N chr2 240813100 N DUP 17
SRR1766446.4905422 chr2 240812886 N chr2 240813035 N DEL 12
SRR1766451.1171433 chr2 240812840 N chr2 240813030 N DEL 12
SRR1766453.903357 chr2 240813025 N chr2 240813100 N DUP 10
SRR1766467.3676091 chr2 240813025 N chr2 240813100 N DUP 13
SRR1766457.3026398 chr2 240812980 N chr2 240813092 N DUP 12
SRR1766470.1657817 chr2 240813049 N chr2 240813181 N DUP 17
SRR1766470.9988440 chr2 240813034 N chr2 240813109 N DUP 11
SRR1766467.4985569 chr2 240813054 N chr2 240813110 N DUP 10
SRR1766451.5293117 chr2 240813025 N chr2 240813100 N DUP 17
SRR1766478.1226564 chr2 240813030 N chr2 240813105 N DUP 11
SRR1766466.4025446 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766479.9068596 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766454.4070858 chr1 222138464 N chr1 222138576 N DUP 12
SRR1766466.2815478 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766465.5134546 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766462.3957041 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766481.9479786 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766455.738276 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766479.10421235 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766481.403046 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766475.11536885 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766472.12031612 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766471.10008279 chr1 222138464 N chr1 222138648 N DUP 10
SRR1766474.2819192 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766447.4359764 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766453.807811 chr1 222138480 N chr1 222138594 N DEL 10
SRR1766453.4410555 chr1 222138464 N chr1 222138720 N DUP 10
SRR1766458.3284469 chr1 222138464 N chr1 222138720 N DUP 10
SRR1766461.7368103 chr1 222138549 N chr1 222138621 N DEL 11
SRR1766458.6167105 chr1 222138621 N chr1 222138716 N DUP 17
SRR1766443.8166889 chr1 222138621 N chr1 222138680 N DUP 17
SRR1766457.7801531 chr1 222138621 N chr1 222138716 N DUP 17
SRR1766463.7371081 chr1 222138621 N chr1 222138716 N DUP 17
SRR1766446.8970471 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766450.1538416 chr1 222138464 N chr1 222138720 N DUP 10
SRR1766455.2840841 chr1 222138681 N chr1 222138874 N DEL 17
SRR1766459.10233140 chr1 222138645 N chr1 222138874 N DEL 17
SRR1766468.6207798 chr1 222138645 N chr1 222138874 N DEL 17
SRR1766460.6807251 chr1 222138645 N chr1 222138874 N DEL 17
SRR1766470.1219278 chr1 222138935 N chr1 222138994 N DUP 12
SRR1766467.3963487 chr1 222138935 N chr1 222138994 N DUP 13
SRR1766485.6487619 chr1 222138935 N chr1 222138994 N DUP 13
SRR1766483.10199415 chr1 222138935 N chr1 222138994 N DUP 13
SRR1766450.6139146 chr1 222138935 N chr1 222138994 N DUP 16
SRR1766467.8566483 chr1 222138935 N chr1 222138994 N DUP 16
SRR1766481.6370041 chr1 222138977 N chr1 222139042 N DEL 19
SRR1766445.6910106 chr1 222138977 N chr1 222139042 N DEL 17
SRR1766453.6593069 chr1 222138413 N chr1 222139043 N DEL 10
SRR1766474.4024607 chr20 59956962 N chr20 59957067 N DEL 13
SRR1766468.5624000 chr16 73349761 N chr16 73349892 N DEL 14
SRR1766449.1820965 chr16 73349791 N chr16 73349847 N DEL 15
SRR1766445.8897429 chr6 39845423 N chr6 39845513 N DUP 10
SRR1766461.2539640 chr22 21307853 N chr22 21307989 N DEL 10
SRR1766478.773293 chr1 248671513 N chr1 248671565 N DEL 10
SRR1766443.3378031 chr1 248671495 N chr1 248671545 N DUP 11
SRR1766460.4100720 chr1 248671597 N chr1 248671649 N DEL 15
SRR1766444.6626282 chr1 248671550 N chr1 248671600 N DUP 10
SRR1766442.26904559 chr1 248671700 N chr1 248671752 N DEL 10
SRR1766444.2414775 chr1 248671617 N chr1 248671667 N DUP 10
SRR1766446.9745601 chr1 248671492 N chr1 248671697 N DEL 10
SRR1766475.3397961 chr1 248671690 N chr1 248671793 N DEL 15
SRR1766454.6453669 chr1 248671649 N chr1 248671854 N DEL 18
SRR1766442.46182949 chr1 248671649 N chr1 248671854 N DEL 17
SRR1766453.7832241 chr1 248671649 N chr1 248671854 N DEL 16
SRR1766452.9269382 chr1 248671649 N chr1 248671854 N DEL 15
SRR1766451.9832788 chr1 248671517 N chr1 248672181 N DEL 11
SRR1766444.6626282 chr1 248671514 N chr1 248672229 N DEL 10
SRR1766456.724119 chr17 75872137 N chr17 75872435 N DEL 14
SRR1766482.436339 chr17 75871906 N chr17 75872205 N DEL 10
SRR1766479.9599377 chr14 82607343 N chr14 82607404 N DUP 10
SRR1766452.9045460 chr14 82607295 N chr14 82607348 N DEL 17
SRR1766470.3626839 chr3 79771313 N chr3 79771366 N DEL 16
SRR1766457.2863696 chr3 79771313 N chr3 79771366 N DEL 16
SRR1766443.4299929 chr3 79771313 N chr3 79771366 N DEL 16
SRR1766442.42521545 chr3 79771313 N chr3 79771366 N DEL 16
SRR1766480.4567817 chr3 79771313 N chr3 79771366 N DEL 14
SRR1766472.3445736 chr3 79771313 N chr3 79771366 N DEL 13
SRR1766446.9308234 chr3 79771313 N chr3 79771366 N DEL 10
SRR1766447.5268777 chr3 79771313 N chr3 79771366 N DEL 10
SRR1766447.9036611 chr3 79771313 N chr3 79771366 N DEL 10
SRR1766475.410540 chr14 73372455 N chr14 73372572 N DUP 11
SRR1766454.4468928 chr3 185234642 N chr3 185234744 N DEL 10
SRR1766473.1042833 chr3 185234642 N chr3 185234744 N DEL 10
SRR1766479.10157233 chr5 113457891 N chr5 113458048 N DUP 10
SRR1766465.4316727 chrX 129915132 N chrX 129915445 N DUP 15
SRR1766484.9613249 chr22 10852268 N chr22 10852461 N DUP 10
SRR1766445.1142379 chr22 10852268 N chr22 10852461 N DUP 10
SRR1766483.5282975 chr18 47366969 N chr18 47367088 N DUP 11
SRR1766457.5688609 chr1 1109035 N chr1 1109127 N DUP 10
SRR1766442.38086200 chr1 1109035 N chr1 1109127 N DUP 16
SRR1766485.3660307 chr9 41772872 N chr9 41772993 N DEL 10
SRR1766459.8409490 chr17 82386500 N chr17 82386569 N DUP 15
SRR1766446.10385175 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766450.11060074 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766463.8032437 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766472.4152114 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766462.10319172 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766460.9634889 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766442.42094979 chr6 52014655 N chr6 52014941 N DEL 13
SRR1766484.11597001 chr6 52014655 N chr6 52014941 N DEL 13
SRR1766466.837833 chr1 22755048 N chr1 22755110 N DUP 13
SRR1766451.4577843 chr1 22754984 N chr1 22755048 N DEL 10
SRR1766484.12287193 chr4 180390409 N chr4 180390936 N DEL 11
SRR1766450.194875 chr4 180390409 N chr4 180390936 N DEL 12
SRR1766459.4419610 chr4 180390409 N chr4 180390936 N DEL 13
SRR1766471.7443098 chr4 180390409 N chr4 180390936 N DEL 12
SRR1766460.9806584 chr4 180390409 N chr4 180390936 N DEL 15
SRR1766452.9299665 chr4 180390409 N chr4 180390936 N DEL 15
SRR1766450.10652025 chr4 180390409 N chr4 180390936 N DEL 15
SRR1766479.139386 chr4 180390409 N chr4 180390936 N DEL 15
SRR1766472.3155088 chr4 180390444 N chr4 180390809 N DEL 14
SRR1766459.4403780 chr4 180390452 N chr4 180390887 N DEL 19
SRR1766451.438492 chr4 180390414 N chr4 180391137 N DUP 11
SRR1766459.5624152 chr4 180390380 N chr4 180390533 N DUP 13
SRR1766483.6671724 chr4 180390380 N chr4 180390533 N DUP 13
SRR1766453.944544 chr4 180390470 N chr4 180390925 N DEL 14
SRR1766477.1269157 chr4 180390393 N chr4 180390452 N DEL 10
SRR1766463.7852344 chr4 180390554 N chr4 180390971 N DUP 12
SRR1766453.175560 chr4 180390563 N chr4 180391010 N DEL 17
SRR1766464.5492340 chr4 180390565 N chr4 180391028 N DEL 10
SRR1766463.10119812 chr4 180390380 N chr4 180390577 N DUP 13
SRR1766463.2829584 chr4 180390531 N chr4 180390598 N DEL 19
SRR1766476.542262 chr4 180390413 N chr4 180390488 N DEL 11
SRR1766464.10665890 chr4 180390425 N chr4 180390488 N DEL 10
SRR1766447.4650057 chr4 180390505 N chr4 180391050 N DUP 16
SRR1766473.4308230 chr4 180390544 N chr4 180390617 N DUP 14
SRR1766445.2808920 chr4 180390521 N chr4 180390608 N DEL 12
SRR1766442.15525373 chr4 180390582 N chr4 180390651 N DUP 19
SRR1766463.10231352 chr4 180390544 N chr4 180390617 N DUP 14
SRR1766465.5096490 chr4 180390522 N chr4 180391031 N DUP 16
SRR1766453.8198161 chr4 180390554 N chr4 180390663 N DUP 16
SRR1766447.4244409 chr4 180390522 N chr4 180391031 N DUP 15
SRR1766462.7298785 chr4 180390410 N chr4 180390506 N DEL 15
SRR1766443.2526497 chr4 180390585 N chr4 180390654 N DUP 19
SRR1766459.5463201 chr4 180390522 N chr4 180391031 N DUP 13
SRR1766472.6517602 chr4 180390544 N chr4 180390637 N DUP 14
SRR1766463.10231352 chr4 180390401 N chr4 180390500 N DEL 10
SRR1766462.5206312 chr4 180390532 N chr4 180390597 N DUP 10
SRR1766467.9349849 chr4 180390575 N chr4 180390646 N DUP 17
SRR1766467.9349849 chr4 180390557 N chr4 180390658 N DUP 19
SRR1766443.3998687 chr4 180390598 N chr4 180391109 N DUP 11
SRR1766476.10044986 chr4 180390532 N chr4 180390597 N DUP 10
SRR1766448.6423808 chr4 180390627 N chr4 180390816 N DEL 10
SRR1766464.2668361 chr4 180390544 N chr4 180390637 N DUP 14
SRR1766456.4045381 chr4 180390530 N chr4 180391208 N DUP 19
SRR1766474.9021775 chr4 180390454 N chr4 180390669 N DUP 15
SRR1766470.8122318 chr4 180390376 N chr4 180390626 N DUP 15
SRR1766475.3706410 chr4 180390425 N chr4 180390544 N DEL 10
SRR1766461.6673320 chr4 180390576 N chr4 180390639 N DUP 16
SRR1766451.379061 chr4 180390564 N chr4 180391210 N DUP 12
SRR1766484.828261 chr4 180390474 N chr4 180390595 N DUP 16
SRR1766445.2102350 chr4 180390407 N chr4 180390498 N DEL 11
SRR1766466.5507101 chr4 180390510 N chr4 180390839 N DUP 11
SRR1766457.4507058 chr4 180390598 N chr4 180391059 N DUP 18
SRR1766446.30308 chr4 180390401 N chr4 180390534 N DEL 10
SRR1766467.10523921 chr4 180390544 N chr4 180390595 N DUP 14
SRR1766473.8686144 chr4 180390544 N chr4 180390595 N DUP 14
SRR1766453.989434 chr4 180390428 N chr4 180390569 N DEL 10
SRR1766442.37506877 chr4 180390532 N chr4 180390619 N DUP 13
SRR1766461.11144720 chr4 180390600 N chr4 180391029 N DUP 15
SRR1766483.1096213 chr4 180390569 N chr4 180391050 N DUP 17
SRR1766475.5697602 chr4 180390376 N chr4 180390626 N DUP 16
SRR1766452.2108395 chr4 180390607 N chr4 180391036 N DUP 17
SRR1766454.5424402 chr4 180390604 N chr4 180390994 N DEL 18
SRR1766476.8110657 chr4 180390544 N chr4 180390637 N DUP 15
SRR1766445.463633 chr4 180390575 N chr4 180390644 N DUP 18
SRR1766472.1079366 chr4 180390646 N chr4 180390994 N DEL 12
SRR1766458.2769907 chr4 180390544 N chr4 180390627 N DUP 15
SRR1766442.11889975 chr4 180390505 N chr4 180391050 N DUP 16
SRR1766484.11305872 chr4 180390598 N chr4 180390875 N DUP 10
SRR1766458.6553799 chr4 180390538 N chr4 180390646 N DUP 19
SRR1766466.7114130 chr4 180390522 N chr4 180390733 N DUP 14
SRR1766477.4294853 chr4 180390505 N chr4 180390738 N DUP 15
SRR1766442.2995494 chr4 180390609 N chr4 180390660 N DEL 18
SRR1766463.9271647 chr4 180390454 N chr4 180390541 N DUP 10
SRR1766446.3164411 chr4 180390618 N chr4 180390691 N DUP 14
SRR1766472.8600641 chr4 180390551 N chr4 180391066 N DUP 17
SRR1766448.5019961 chr4 180390551 N chr4 180391066 N DUP 17
SRR1766467.10246740 chr4 180390551 N chr4 180391066 N DUP 17
SRR1766478.1118388 chr4 180390628 N chr4 180390691 N DUP 14
SRR1766477.9996967 chr4 180390554 N chr4 180390745 N DUP 17
SRR1766471.5188130 chr4 180390554 N chr4 180390745 N DUP 14
SRR1766455.7549782 chr4 180390595 N chr4 180390866 N DEL 15
SRR1766481.7475507 chr4 180390893 N chr4 180390979 N DUP 16
SRR1766482.9747182 chr4 180390893 N chr4 180390979 N DUP 16
SRR1766481.6054022 chr4 180390556 N chr4 180391077 N DUP 12
SRR1766476.10967478 chr4 180390556 N chr4 180391077 N DUP 13
SRR1766453.944544 chr4 180390468 N chr4 180391067 N DUP 11
SRR1766443.6415213 chr4 180390595 N chr4 180391012 N DEL 18
SRR1766476.9582469 chr4 180390628 N chr4 180390691 N DUP 14
SRR1766483.12416279 chr4 180390973 N chr4 180391024 N DUP 16
SRR1766463.8309583 chr4 180390942 N chr4 180391027 N DUP 13
SRR1766463.9279167 chr4 180390935 N chr4 180391050 N DUP 15
SRR1766481.13197869 chr4 180390538 N chr4 180391051 N DUP 15
SRR1766470.3960076 chr4 180390546 N chr4 180391109 N DUP 13
SRR1766469.1276665 chr4 180390838 N chr4 180390980 N DEL 12
SRR1766479.8971394 chr4 180390936 N chr4 180391103 N DUP 11
SRR1766442.33295538 chr4 180390988 N chr4 180391087 N DUP 18
SRR1766454.7691693 chr4 180390574 N chr4 180391087 N DUP 10
SRR1766486.6814917 chr4 180390988 N chr4 180391087 N DUP 15
SRR1766478.2978765 chr4 180390502 N chr4 180391089 N DUP 13
SRR1766468.6005559 chr4 180390981 N chr4 180391068 N DUP 14
SRR1766469.8261919 chr4 180391005 N chr4 180391094 N DUP 17
SRR1766475.6965280 chr4 180391005 N chr4 180391094 N DUP 17
SRR1766484.2489579 chr4 180390685 N chr4 180391169 N DEL 12
SRR1766478.5627240 chr4 180390553 N chr4 180391181 N DEL 17
SRR1766442.46293936 chr4 180390413 N chr4 180391213 N DEL 10
SRR1766474.4166687 chr4 180390413 N chr4 180391213 N DEL 10
SRR1766442.33369200 chr4 180390413 N chr4 180391213 N DEL 10
SRR1766458.6553799 chr4 180390413 N chr4 180391213 N DEL 10
SRR1766454.3828767 chr4 180390387 N chr4 180391224 N DEL 15
SRR1766450.2182247 chr2 2750311 N chr2 2750440 N DUP 18
SRR1766483.3248156 chr2 2750547 N chr2 2750603 N DEL 15
SRR1766466.9420768 chr2 2750547 N chr2 2750603 N DEL 17
SRR1766453.356498 chr2 2750547 N chr2 2750603 N DEL 17
SRR1766442.22281966 chr2 2750547 N chr2 2750603 N DEL 17
SRR1766472.10192678 chr2 2750547 N chr2 2750603 N DEL 17
SRR1766463.10329068 chr17 79701428 N chr17 79701565 N DEL 19
SRR1766465.6622716 chr17 79701377 N chr17 79701898 N DEL 10
SRR1766461.2921576 chr6 162010639 N chr6 162010715 N DUP 10
SRR1766454.376527 chr6 162010639 N chr6 162010715 N DUP 10
SRR1766479.4048513 chr6 162010690 N chr6 162011085 N DUP 11
SRR1766448.3475578 chr6 162010638 N chr6 162010721 N DUP 19
SRR1766464.10151878 chr6 162010742 N chr6 162010859 N DUP 15
SRR1766472.2579692 chr6 162010726 N chr6 162010863 N DUP 16
SRR1766461.5979337 chr6 162010736 N chr6 162011095 N DUP 11
SRR1766459.2315868 chr6 162010729 N chr6 162010806 N DUP 17
SRR1766458.6783959 chr6 162010730 N chr6 162010929 N DUP 16
SRR1766442.24017496 chr6 162011193 N chr6 162011641 N DUP 17
SRR1766452.15055 chr6 162011200 N chr6 162011285 N DEL 14
SRR1766476.4651601 chr21 44592020 N chr21 44592376 N DUP 10
SRR1766483.8148887 chr21 44592020 N chr21 44592376 N DUP 10
SRR1766472.9101274 chr21 44592020 N chr21 44592376 N DUP 10
SRR1766483.5298277 chr21 44592020 N chr21 44592376 N DUP 10
SRR1766450.985912 chr21 44592023 N chr21 44592379 N DUP 10
SRR1766473.8103408 chr10 62370442 N chr10 62371227 N DEL 18
SRR1766474.9835975 chr10 62370456 N chr10 62370520 N DEL 14
SRR1766483.1161636 chr10 62370456 N chr10 62370520 N DEL 14
SRR1766442.10435810 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766482.4763274 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766442.44983845 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766472.6901547 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766481.11281261 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766479.5205598 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766451.6475581 chr10 62370459 N chr10 62371349 N DUP 13
SRR1766454.5464023 chr10 62370472 N chr10 62370556 N DUP 12
SRR1766472.7780208 chr10 62370472 N chr10 62370556 N DUP 12
SRR1766469.9363987 chr10 62370439 N chr10 62370606 N DUP 10
SRR1766468.4165849 chr10 62370628 N chr10 62370685 N DUP 16
SRR1766486.2026388 chr10 62370607 N chr10 62371260 N DUP 18
SRR1766483.7509108 chr10 62370489 N chr10 62370689 N DEL 14
SRR1766463.2283060 chr10 62370489 N chr10 62370689 N DEL 14
SRR1766450.4901618 chr10 62370489 N chr10 62370689 N DEL 13
SRR1766467.11907405 chr10 62370791 N chr10 62370869 N DEL 11
SRR1766460.6498764 chr10 62370791 N chr10 62370869 N DEL 12
SRR1766449.408250 chr10 62370791 N chr10 62370869 N DEL 12
SRR1766483.3007261 chr10 62370707 N chr10 62370801 N DUP 13
SRR1766446.8689418 chr10 62370707 N chr10 62370801 N DUP 13
SRR1766475.3600823 chr10 62370707 N chr10 62370801 N DUP 13
SRR1766460.3236897 chr10 62370997 N chr10 62371319 N DUP 14
SRR1766477.7288064 chr10 62370997 N chr10 62371319 N DUP 14
SRR1766478.9704075 chr10 62370998 N chr10 62371320 N DUP 13
SRR1766474.1030344 chr10 62371134 N chr10 62371189 N DUP 17
SRR1766472.10783213 chr10 62371208 N chr10 62371297 N DUP 17
SRR1766442.38681972 chr10 62371208 N chr10 62371297 N DUP 16
SRR1766458.2012467 chr10 62370572 N chr10 62371128 N DEL 17
SRR1766460.4981163 chr10 62370544 N chr10 62371226 N DEL 11
SRR1766447.2680118 chr10 62370544 N chr10 62371226 N DEL 11
SRR1766459.5340769 chr10 62371035 N chr10 62371289 N DUP 11
SRR1766449.9354824 chr10 62370574 N chr10 62371227 N DEL 15
SRR1766463.9309583 chr10 62370641 N chr10 62371350 N DUP 10
SRR1766472.1990295 chr10 62370641 N chr10 62371350 N DUP 10
SRR1766442.23639227 chr10 62370661 N chr10 62371350 N DUP 12
SRR1766459.7640060 chr10 62370661 N chr10 62371350 N DUP 13
SRR1766468.7101019 chr10 62370661 N chr10 62371350 N DUP 15
SRR1766447.3273557 chr10 62370661 N chr10 62371350 N DUP 16
SRR1766470.4571153 chr10 62370661 N chr10 62371350 N DUP 18
SRR1766475.6643257 chr10 62370463 N chr10 62371362 N DUP 14
SRR1766442.16091078 chr10 62370463 N chr10 62371362 N DUP 16
SRR1766472.100128 chr10 62371441 N chr10 62371531 N DUP 17
SRR1766449.1569407 chr10 62371147 N chr10 62371401 N DEL 11
SRR1766472.2210632 chr10 62371147 N chr10 62371401 N DEL 12
SRR1766442.35009943 chr10 62371342 N chr10 62371419 N DEL 17
SRR1766483.8121208 chr10 62370450 N chr10 62371423 N DEL 11
SRR1766470.4571153 chr10 62371362 N chr10 62371499 N DEL 14
SRR1766443.3644545 chr10 62371362 N chr10 62371499 N DEL 11
SRR1766472.4502727 chr10 62370389 N chr10 62371471 N DEL 12
SRR1766485.6747037 chr10 62371362 N chr10 62371499 N DEL 19
SRR1766446.2942575 chr10 62371362 N chr10 62371499 N DEL 19
SRR1766456.5460621 chr10 62370536 N chr10 62371499 N DEL 16
SRR1766446.9787988 chr10 62371365 N chr10 62371520 N DEL 19
SRR1766463.9309583 chr10 62371365 N chr10 62371520 N DEL 19
SRR1766450.8728826 chr10 62371343 N chr10 62371520 N DEL 13
SRR1766447.3718226 chr10 62370457 N chr10 62371521 N DEL 12
SRR1766476.10094059 chr10 62370458 N chr10 62371522 N DEL 12
SRR1766462.6477231 chr10 62370450 N chr10 62371523 N DEL 11
SRR1766478.3632890 chr9 89254390 N chr9 89254628 N DUP 16
SRR1766471.1406341 chr9 89254362 N chr9 89254418 N DUP 10
SRR1766471.11312798 chr9 89254135 N chr9 89254628 N DUP 12
SRR1766444.3368329 chr9 89254391 N chr9 89254640 N DEL 12
SRR1766464.8671432 chr9 89254332 N chr9 89254813 N DEL 10
SRR1766473.8416303 chr9 86463042 N chr9 86463123 N DUP 11
SRR1766465.543609 chr9 86463063 N chr9 86463130 N DEL 17
SRR1766474.722261 chr9 86463063 N chr9 86463130 N DEL 17
SRR1766442.30482406 chr9 86463063 N chr9 86463130 N DEL 16
SRR1766479.6879434 chr9 86463065 N chr9 86463132 N DEL 11
SRR1766459.9487662 chr9 86463062 N chr9 86463133 N DEL 11
SRR1766477.9032097 chr13 83380677 N chr13 83380782 N DEL 11
SRR1766481.12524624 chr13 83380656 N chr13 83380865 N DEL 10
SRR1766460.10782732 chr21 41806374 N chr21 41806690 N DEL 11
SRR1766442.4372818 chr21 41806210 N chr21 41806290 N DUP 10
SRR1766482.13240996 chr21 41806383 N chr21 41806454 N DEL 17
SRR1766481.8927194 chr21 41806151 N chr21 41806327 N DUP 17
SRR1766469.9926387 chr21 41806325 N chr21 41806417 N DEL 16
SRR1766473.8889776 chr21 41806489 N chr21 41806547 N DEL 18
SRR1766445.566274 chr21 41806307 N chr21 41806426 N DEL 16
SRR1766476.3703027 chr21 41806186 N chr21 41806242 N DUP 17
SRR1766476.7958269 chr21 41806210 N chr21 41806546 N DUP 16
SRR1766444.611543 chr21 41806183 N chr21 41806238 N DEL 12
SRR1766484.2166193 chr21 41806323 N chr21 41806639 N DEL 18
SRR1766452.9152131 chr21 41806263 N chr21 41806334 N DUP 14
SRR1766445.1901079 chr21 41806288 N chr21 41806362 N DUP 19
SRR1766442.44317868 chr21 41806255 N chr21 41806727 N DUP 12
SRR1766442.31815950 chr21 41806169 N chr21 41806331 N DUP 14
SRR1766474.10598312 chr21 41806169 N chr21 41806239 N DEL 11
SRR1766446.2582196 chr21 41806135 N chr21 41806253 N DEL 10
SRR1766479.4774370 chr21 41806214 N chr21 41806282 N DUP 10
SRR1766470.8640975 chr21 41806195 N chr21 41806585 N DUP 13
SRR1766461.10308705 chr21 41806169 N chr21 41806331 N DUP 14
SRR1766446.8352937 chr21 41806246 N chr21 41806302 N DUP 13
SRR1766474.6163715 chr21 41806182 N chr21 41806343 N DUP 10
SRR1766480.3595308 chr21 41806222 N chr21 41806443 N DEL 16
SRR1766456.5892728 chr21 41806210 N chr21 41806495 N DUP 10
SRR1766463.9678769 chr21 41806210 N chr21 41806350 N DUP 12
SRR1766462.507819 chr21 41806216 N chr21 41806329 N DUP 13
SRR1766460.5737883 chr21 41806331 N chr21 41806536 N DEL 19
SRR1766451.6119418 chr21 41806207 N chr21 41806323 N DUP 19
SRR1766479.4774370 chr21 41806360 N chr21 41806753 N DEL 10
SRR1766442.19177731 chr21 41806140 N chr21 41806544 N DEL 12
SRR1766442.35918755 chr21 41806152 N chr21 41806306 N DEL 12
SRR1766461.6400848 chr21 41806239 N chr21 41806694 N DUP 10
SRR1766486.3566662 chr21 41806135 N chr21 41806253 N DEL 12
SRR1766455.5441746 chr21 41806195 N chr21 41806368 N DUP 17
SRR1766454.9188359 chr21 41806337 N chr21 41806417 N DEL 19
SRR1766467.2469423 chr21 41806222 N chr21 41806775 N DUP 15
SRR1766471.7782337 chr21 41806216 N chr21 41806329 N DUP 13
SRR1766452.5411341 chr21 41806228 N chr21 41806320 N DUP 15
SRR1766467.6093453 chr21 41806462 N chr21 41806581 N DUP 12
SRR1766452.4513262 chr21 41806195 N chr21 41806293 N DUP 14
SRR1766483.6090902 chr21 41806284 N chr21 41806764 N DEL 18
SRR1766447.7925912 chr21 41806198 N chr21 41806683 N DUP 10
SRR1766455.504532 chr21 41806201 N chr21 41806365 N DUP 12
SRR1766449.1067258 chr21 41806161 N chr21 41806228 N DEL 12
SRR1766455.5792477 chr21 41806243 N chr21 41806308 N DUP 10
SRR1766447.2395898 chr21 41806194 N chr21 41806752 N DEL 14
SRR1766485.6322990 chr21 41806240 N chr21 41806380 N DUP 12
SRR1766481.4157761 chr21 41806162 N chr21 41806380 N DUP 10
SRR1766470.4625374 chr21 41806196 N chr21 41806720 N DUP 10
SRR1766456.3360709 chr21 41806237 N chr21 41806323 N DUP 12
SRR1766462.6370980 chr21 41806181 N chr21 41806303 N DUP 12
SRR1766479.12294387 chr21 41806150 N chr21 41806772 N DUP 13
SRR1766474.5784086 chr21 41806254 N chr21 41806448 N DEL 12
SRR1766442.39351101 chr21 41806222 N chr21 41806392 N DUP 11
SRR1766442.3101599 chr21 41806209 N chr21 41806593 N DUP 13
SRR1766473.2361154 chr21 41806195 N chr21 41806329 N DUP 18
SRR1766448.5043384 chr21 41806351 N chr21 41806521 N DEL 17
SRR1766483.2245272 chr21 41806143 N chr21 41806228 N DEL 16
SRR1766470.7074814 chr21 41806136 N chr21 41806336 N DUP 17
SRR1766442.12570152 chr21 41806241 N chr21 41806757 N DEL 13
SRR1766464.5726126 chr21 41806291 N chr21 41806683 N DUP 13
SRR1766457.9369004 chr21 41806490 N chr21 41806564 N DUP 17
SRR1766460.650262 chr21 41806213 N chr21 41806719 N DUP 13
SRR1766447.1323725 chr21 41806182 N chr21 41806343 N DUP 13
SRR1766448.9185457 chr21 41806198 N chr21 41806359 N DUP 14
SRR1766442.43917223 chr21 41806306 N chr21 41806829 N DUP 16
SRR1766466.6208572 chr21 41806155 N chr21 41806235 N DUP 12
SRR1766454.8334503 chr21 41806246 N chr21 41806634 N DEL 11
SRR1766469.7286902 chr21 41806159 N chr21 41806227 N DUP 12
SRR1766443.3255838 chr21 41806418 N chr21 41806769 N DUP 11
SRR1766473.11579232 chr21 41806182 N chr21 41806667 N DUP 10
SRR1766459.2526939 chr21 41806258 N chr21 41806323 N DUP 12
SRR1766470.8640975 chr21 41806220 N chr21 41806693 N DUP 18
SRR1766452.10527393 chr21 41806140 N chr21 41806544 N DEL 12
SRR1766442.44763926 chr21 41806246 N chr21 41806561 N DUP 10
SRR1766451.1906347 chr21 41806354 N chr21 41806524 N DEL 13
SRR1766449.5210184 chr21 41806182 N chr21 41806283 N DUP 16
SRR1766463.8505495 chr21 41806186 N chr21 41806305 N DUP 10
SRR1766466.8986444 chr21 41806379 N chr21 41806644 N DEL 13
SRR1766454.7733584 chr21 41689406 N chr21 41689463 N DEL 12
SRR1766447.4972719 chr21 41689406 N chr21 41689463 N DEL 17
SRR1766461.2009814 chr21 41689406 N chr21 41689463 N DEL 19
SRR1766474.10444562 chr21 41689406 N chr21 41689463 N DEL 15
SRR1766451.10269866 chr2 237213089 N chr2 237213271 N DEL 15
SRR1766462.2859043 chr2 237213089 N chr2 237213271 N DEL 10
SRR1766483.5364740 chr12 129136984 N chr12 129137040 N DUP 15
SRR1766486.5897967 chr12 129136944 N chr12 129137034 N DEL 14
SRR1766466.8294429 chr12 129137128 N chr12 129137346 N DEL 14
SRR1766462.8529724 chr12 129137305 N chr12 129137373 N DUP 13
SRR1766459.9443173 chr9 29018197 N chr9 29018263 N DUP 13
SRR1766450.766250 chr16 69478630 N chr16 69478679 N DUP 10
SRR1766449.8723641 chr1 143252837 N chr1 143252956 N DUP 13
SRR1766452.10088354 chr1 143252802 N chr1 143252855 N DEL 10
SRR1766482.7535552 chr1 48227437 N chr1 48227719 N DEL 12
SRR1766468.4008914 chr1 48227352 N chr1 48227748 N DUP 10
SRR1766484.10413642 chr1 48227352 N chr1 48227748 N DUP 10
SRR1766458.7365467 chr1 48227439 N chr1 48227670 N DEL 12
SRR1766442.27452924 chr1 48227439 N chr1 48227603 N DEL 14
SRR1766472.9722936 chr1 48227439 N chr1 48227603 N DEL 11
SRR1766457.8538438 chr1 48227452 N chr1 48227616 N DEL 10
SRR1766458.4516773 chr9 43348090 N chr9 43348259 N DUP 10
SRR1766449.5439652 chr13 64512251 N chr13 64512319 N DEL 10
SRR1766452.6196879 chr13 64512282 N chr13 64512348 N DUP 10
SRR1766450.1640922 chr5 43031960 N chr5 43032079 N DEL 14
SRR1766445.2880406 chr5 43031941 N chr5 43032262 N DUP 10
SRR1766485.9416488 chr5 43032123 N chr5 43032195 N DEL 19
SRR1766473.4245758 chr5 43031941 N chr5 43032262 N DUP 15
SRR1766448.2870126 chr5 43031941 N chr5 43032262 N DUP 16
SRR1766473.9068340 chr5 43031941 N chr5 43032262 N DUP 16
SRR1766478.10334282 chr5 43032078 N chr5 43032199 N DUP 19
SRR1766486.8988579 chr5 43032181 N chr5 43032262 N DUP 18
SRR1766453.6605225 chr5 43032181 N chr5 43032262 N DUP 18
SRR1766481.6751386 chr5 43032078 N chr5 43032199 N DUP 16
SRR1766442.4235579 chr5 43031926 N chr5 43032389 N DEL 10
SRR1766457.3913274 chr5 43031900 N chr5 43032391 N DEL 10
SRR1766450.1640922 chr5 43032367 N chr5 43032450 N DEL 16
SRR1766446.8876971 chr5 43032454 N chr5 43032516 N DUP 11
SRR1766443.4607614 chr22 18369679 N chr22 18370310 N DEL 15
SRR1766453.6845333 chr22 18369763 N chr22 18370392 N DUP 13
SRR1766477.10486013 chr22 18369763 N chr22 18370392 N DUP 15
SRR1766480.4704091 chr22 18369829 N chr22 18370460 N DEL 10
SRR1766476.3471834 chr22 18369763 N chr22 18370392 N DUP 10
SRR1766454.430473 chr22 18369829 N chr22 18370460 N DEL 10
SRR1766451.10079258 chr18 57510089 N chr18 57510405 N DEL 11
SRR1766457.3096592 chr18 57510089 N chr18 57510405 N DEL 11
SRR1766470.3025904 chr18 57510089 N chr18 57510405 N DEL 15
SRR1766449.10607714 chr18 57510107 N chr18 57510423 N DEL 19
SRR1766481.6960857 chr18 57510313 N chr18 57510944 N DEL 10
SRR1766459.2202818 chr4 1828666 N chr4 1828920 N DEL 10
SRR1766480.1877353 chr4 1828648 N chr4 1828701 N DEL 17
SRR1766458.6712066 chr4 1828648 N chr4 1828701 N DEL 14
SRR1766460.6051148 chr4 1828648 N chr4 1828701 N DEL 12
SRR1766467.3652921 chr4 1828920 N chr4 1829377 N DUP 10
SRR1766475.2742768 chr4 1828933 N chr4 1829470 N DEL 15
SRR1766452.9664530 chr15 27313378 N chr15 27313443 N DUP 10
SRR1766447.6576208 chr15 27313377 N chr15 27313428 N DUP 10
SRR1766482.5136050 chr18 7984721 N chr18 7984823 N DUP 10
SRR1766449.3861167 chr1 189818374 N chr1 189818441 N DEL 14
SRR1766455.6062088 chr1 189818374 N chr1 189818441 N DEL 15
SRR1766457.7087631 chr1 189818463 N chr1 189818544 N DEL 19
SRR1766481.905479 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766469.7515319 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766445.2964457 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766485.5643203 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766451.8874075 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766472.626444 chr1 189818465 N chr1 189818546 N DEL 13
SRR1766454.10039188 chr1 189818466 N chr1 189818547 N DEL 12
SRR1766442.35552044 chr1 189818615 N chr1 189818692 N DUP 11
SRR1766447.10476117 chr1 189818615 N chr1 189818692 N DUP 13
SRR1766485.12049722 chr1 189818615 N chr1 189818692 N DUP 12
SRR1766470.4120270 chr7 156439918 N chr7 156440012 N DUP 13
SRR1766455.9511091 chr7 156439918 N chr7 156440012 N DUP 14
SRR1766484.11084322 chr7 156439918 N chr7 156440012 N DUP 16
SRR1766475.7520862 chr15 101763980 N chr15 101764167 N DUP 10
SRR1766448.5979964 chr15 101763979 N chr15 101764168 N DEL 10
SRR1766455.4302704 chr15 101764319 N chr15 101764411 N DEL 10
SRR1766460.123773 chr15 101764013 N chr15 101764114 N DEL 10
SRR1766465.10950306 chr15 101764342 N chr15 101764434 N DEL 15
SRR1766467.7537170 chr15 101764319 N chr15 101764411 N DEL 10
SRR1766457.3751975 chr1 248840752 N chr1 248841239 N DEL 10
SRR1766453.1492532 chr1 248840759 N chr1 248840814 N DEL 10
SRR1766452.10515502 chr1 248840768 N chr1 248841039 N DEL 10
SRR1766460.8491756 chr1 248840931 N chr1 248841040 N DEL 15
SRR1766457.3751975 chr1 248841158 N chr1 248841211 N DUP 15
SRR1766448.6656103 chr20 46491826 N chr20 46492391 N DEL 10
SRR1766475.4687221 chr20 46491704 N chr20 46492269 N DEL 14
SRR1766482.5618929 chr20 46491924 N chr20 46492489 N DEL 10
SRR1766444.1779596 chr9 96026767 N chr9 96027098 N DEL 14
SRR1766464.7057425 chr9 96026835 N chr9 96026914 N DEL 10
SRR1766446.7607364 chr16 16650860 N chr16 16650921 N DEL 11
SRR1766458.1908230 chr15 50635468 N chr15 50635823 N DUP 12
SRR1766456.4605365 chr5 3856913 N chr5 3856964 N DEL 19
SRR1766462.1133999 chr5 3856913 N chr5 3856964 N DEL 16
SRR1766450.8934125 chr5 3856917 N chr5 3856968 N DEL 11
SRR1766445.9705740 chr5 3856915 N chr5 3856966 N DEL 13
SRR1766450.340076 chr5 3856914 N chr5 3856965 N DEL 14
SRR1766463.388858 chr5 3856914 N chr5 3856965 N DEL 14
SRR1766484.5640815 chr10 49965668 N chr10 49966225 N DEL 15
SRR1766470.955295 chr10 49965668 N chr10 49966225 N DEL 15
SRR1766451.9536241 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766457.5140021 chr5 10347422 N chr5 10347479 N DUP 10
SRR1766479.4915557 chr5 10347121 N chr5 10347406 N DEL 14
SRR1766455.4745641 chr5 10347459 N chr5 10347518 N DEL 10
SRR1766457.2314894 chr5 10346474 N chr5 10346553 N DEL 19
SRR1766454.598117 chr5 10347096 N chr5 10347406 N DEL 16
SRR1766445.6967072 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766486.10573528 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766442.5346800 chr5 10347096 N chr5 10347406 N DEL 16
SRR1766486.5371104 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766448.4911493 chr5 10347459 N chr5 10347518 N DEL 10
SRR1766475.3765078 chr5 10347459 N chr5 10347518 N DEL 10
SRR1766462.85102 chr5 10347121 N chr5 10347406 N DEL 14
SRR1766472.603517 chr5 10347422 N chr5 10347479 N DUP 19
SRR1766471.467521 chr5 10347117 N chr5 10347398 N DEL 14
SRR1766444.4825970 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766453.3510036 chr5 10347462 N chr5 10347521 N DEL 10
SRR1766442.27003599 chr5 10347422 N chr5 10347479 N DUP 17
SRR1766464.6603080 chr5 10347121 N chr5 10347406 N DEL 11
SRR1766442.1088889 chr5 10346474 N chr5 10346553 N DEL 18
SRR1766465.11248369 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766461.8476723 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766473.9018190 chr5 10347121 N chr5 10347406 N DEL 12
SRR1766464.6603080 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766450.2372217 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766485.11054307 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766467.6090314 chr5 10347096 N chr5 10347406 N DEL 16
SRR1766466.178559 chr5 10347459 N chr5 10347518 N DEL 10
SRR1766470.5490836 chr5 10347459 N chr5 10347518 N DEL 15
SRR1766445.4449075 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766450.7122101 chr5 10347096 N chr5 10347406 N DEL 16
SRR1766473.7110824 chr17 32227782 N chr17 32227895 N DUP 14
SRR1766457.321800 chr13 62019547 N chr13 62019606 N DEL 12
SRR1766460.7246157 chr13 62019772 N chr13 62019847 N DUP 13
SRR1766482.12705189 chr13 62019790 N chr13 62019849 N DUP 11
SRR1766457.5752772 chr14 56355292 N chr14 56355345 N DUP 12
SRR1766464.7165385 chr14 56355301 N chr14 56355402 N DUP 15
SRR1766449.830077 chr14 56355301 N chr14 56355402 N DUP 14
SRR1766442.37521161 chr14 56355301 N chr14 56355402 N DUP 15
SRR1766476.7815557 chr14 56355337 N chr14 56355420 N DUP 14
SRR1766473.10082444 chr14 56355337 N chr14 56355420 N DUP 14
SRR1766445.417605 chr14 56355337 N chr14 56355420 N DUP 19
SRR1766452.6695738 chr14 56355377 N chr14 56355452 N DEL 15
SRR1766471.10971266 chr14 56355377 N chr14 56355452 N DEL 15
SRR1766468.5157910 chr14 56355377 N chr14 56355452 N DEL 15
SRR1766442.27903440 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766459.917116 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766459.5558079 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766442.18099783 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766454.123169 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766460.9076839 chr14 56355331 N chr14 56355452 N DEL 15
SRR1766471.7382822 chr14 56355331 N chr14 56355452 N DEL 19
SRR1766442.12914548 chr14 56355313 N chr14 56355452 N DEL 10
SRR1766452.1701095 chr14 56355313 N chr14 56355452 N DEL 10
SRR1766448.8583577 chr14 56355315 N chr14 56355454 N DEL 10
SRR1766451.3735200 chr14 56355315 N chr14 56355454 N DEL 10
SRR1766442.31185038 chr14 56355316 N chr14 56355455 N DEL 10
SRR1766455.7262819 chr3 106073719 N chr3 106074033 N DEL 10
SRR1766442.3069708 chr3 106073938 N chr3 106074161 N DEL 10
SRR1766452.326692 chr3 106073938 N chr3 106074161 N DEL 10
SRR1766449.6523629 chr3 106073690 N chr3 106074400 N DUP 10
SRR1766448.8153443 chr3 106073691 N chr3 106074401 N DUP 13
SRR1766480.6954657 chr10 106718904 N chr10 106718971 N DEL 15
SRR1766443.6792589 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766470.149485 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766476.786500 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766468.1825976 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766442.8411782 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766479.7063926 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766479.2115776 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766448.10918086 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766458.7373508 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766483.6157318 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766482.6638258 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766469.6912644 chr10 106719000 N chr10 106719133 N DEL 15
SRR1766454.338703 chr10 106719000 N chr10 106719133 N DEL 15
SRR1766483.4855414 chr10 106719000 N chr10 106719133 N DEL 15
SRR1766452.6467156 chr10 106719000 N chr10 106719133 N DEL 15
SRR1766470.11190758 chr8 29667216 N chr8 29667317 N DUP 13
SRR1766461.4456442 chr8 29666962 N chr8 29667289 N DEL 11
SRR1766451.5456172 chr6 158705646 N chr6 158705803 N DUP 11
SRR1766486.3590123 chr3 5135493 N chr3 5135670 N DUP 11
SRR1766462.6112610 chrX 33010119 N chrX 33010180 N DEL 18
SRR1766442.39320619 chrX 33010119 N chrX 33010180 N DEL 18
SRR1766471.1964679 chrX 33010120 N chrX 33010181 N DEL 13
SRR1766471.6413838 chrX 33010120 N chrX 33010181 N DEL 13
SRR1766455.1942686 chrX 33010095 N chrX 33010198 N DEL 10
SRR1766453.997981 chrX 123846064 N chrX 123846373 N DEL 10
SRR1766481.5939938 chr7 56367950 N chr7 56368096 N DEL 10
SRR1766483.533353 chr7 56367860 N chr7 56368088 N DEL 11
SRR1766472.5122703 chr7 157057325 N chr7 157057548 N DUP 10
SRR1766461.11082585 chr3 128955025 N chr3 128955252 N DEL 10
SRR1766464.3991584 chr3 128955025 N chr3 128955252 N DEL 10
SRR1766457.9455848 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766442.23936417 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766463.988270 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766462.8210323 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766452.6744293 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766455.8565815 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766448.10239597 chr12 12944892 N chr12 12944950 N DEL 10
SRR1766442.33013779 chr12 12944892 N chr12 12944950 N DEL 15
SRR1766479.11636452 chr12 12944896 N chr12 12944950 N DEL 12
SRR1766474.6293010 chr12 12944896 N chr12 12944950 N DEL 13
SRR1766486.5234875 chr10 15149213 N chr10 15149439 N DUP 10
SRR1766442.17362096 chr10 15149213 N chr10 15149439 N DUP 10
SRR1766442.27007108 chr10 15149353 N chr10 15149410 N DEL 11
SRR1766462.6108573 chr10 15149414 N chr10 15149532 N DUP 14
SRR1766483.3418252 chr10 15149320 N chr10 15149584 N DUP 11
SRR1766459.3240647 chr10 15149414 N chr10 15149532 N DUP 14
SRR1766484.9770339 chr10 15149414 N chr10 15149532 N DUP 18
SRR1766465.5263945 chr10 15149414 N chr10 15149532 N DUP 19
SRR1766480.425796 chr10 15149593 N chr10 15149658 N DUP 15
SRR1766460.1628626 chr10 15149531 N chr10 15149592 N DEL 19
SRR1766447.6190164 chr10 15149464 N chr10 15149693 N DUP 17
SRR1766478.1232114 chr10 15149597 N chr10 15149698 N DUP 13
SRR1766460.8561626 chr10 15149531 N chr10 15149598 N DEL 15
SRR1766450.9178643 chr10 15149531 N chr10 15149598 N DEL 16
SRR1766449.5700154 chr10 15149622 N chr10 15149690 N DUP 12
SRR1766486.5771749 chr10 15149654 N chr10 15149716 N DUP 12
SRR1766445.8698855 chr10 15149345 N chr10 15149735 N DUP 14
SRR1766470.1082725 chr10 15149498 N chr10 15149628 N DEL 19
SRR1766472.3522019 chr10 15149655 N chr10 15149726 N DUP 14
SRR1766463.2112154 chr10 15149597 N chr10 15149698 N DUP 12
SRR1766480.3315942 chr10 15149501 N chr10 15149649 N DEL 12
SRR1766475.4714776 chr10 15149679 N chr10 15149738 N DUP 10
SRR1766486.1050257 chr10 15149601 N chr10 15149699 N DUP 17
SRR1766463.5798224 chr10 15149222 N chr10 15149750 N DUP 11
SRR1766458.2349347 chr10 15149662 N chr10 15149742 N DUP 10
SRR1766450.3578925 chr10 15149630 N chr10 15149712 N DEL 10
SRR1766470.7172163 chr14 104720558 N chr14 104720696 N DEL 16
SRR1766461.7718003 chr14 104720523 N chr14 104720696 N DEL 13
SRR1766470.7353141 chr14 104720523 N chr14 104720696 N DEL 10
SRR1766484.4619882 chr14 104720491 N chr14 104721208 N DUP 13
SRR1766459.10691782 chr14 104720491 N chr14 104721208 N DUP 13
SRR1766484.11737318 chr14 104720561 N chr14 104721208 N DUP 13
SRR1766448.1320047 chr14 104720601 N chr14 104721286 N DUP 10
SRR1766442.41069344 chr14 104720516 N chr14 104720905 N DEL 13
SRR1766445.141934 chr1 2142471 N chr1 2142557 N DEL 15
SRR1766469.8249993 chr1 2142471 N chr1 2142557 N DEL 15
SRR1766480.86281 chr1 2142075 N chr1 2142581 N DEL 16
SRR1766484.7670346 chr1 2142471 N chr1 2142557 N DEL 12
SRR1766453.7730850 chr1 2142471 N chr1 2142557 N DEL 14
SRR1766459.10597847 chr1 2142075 N chr1 2142581 N DEL 11
SRR1766469.5569084 chr10 10462637 N chr10 10462767 N DEL 13
SRR1766470.6498967 chr10 10462637 N chr10 10462768 N DEL 12
SRR1766454.10663833 chr2 83914609 N chr2 83914757 N DUP 10
SRR1766472.11313346 chr2 83914513 N chr2 83914756 N DUP 14
SRR1766450.4542906 chr2 83914513 N chr2 83914756 N DUP 18
SRR1766482.4114782 chr8 140120705 N chr8 140120870 N DEL 12
SRR1766459.805884 chr4 713574 N chr4 713627 N DEL 15
SRR1766460.2709101 chr9 136307873 N chr9 136308959 N DEL 10
SRR1766468.2447764 chr9 136307506 N chr9 136307914 N DEL 10
SRR1766453.10487929 chr9 136308044 N chr9 136308226 N DEL 14
SRR1766469.8541234 chr9 136308199 N chr9 136308393 N DEL 10
SRR1766484.9000563 chr9 136307980 N chr9 136308161 N DUP 12
SRR1766463.10099757 chr9 136308044 N chr9 136308226 N DEL 17
SRR1766448.6450734 chr9 136307490 N chr9 136308435 N DUP 10
SRR1766460.472459 chr9 136307927 N chr9 136308505 N DEL 12
SRR1766482.11133851 chr9 136308509 N chr9 136308579 N DUP 12
SRR1766479.9441339 chr9 136307505 N chr9 136308536 N DEL 13
SRR1766453.9354321 chr9 136308547 N chr9 136309178 N DUP 15
SRR1766470.2536131 chr9 136308307 N chr9 136308783 N DEL 10
SRR1766450.4962109 chr2 152923103 N chr2 152923271 N DUP 12
SRR1766452.8931481 chrX 71740761 N chrX 71741098 N DEL 11
SRR1766474.1176446 chrX 71740802 N chrX 71741152 N DEL 12
SRR1766474.6727292 chrX 71741215 N chrX 71741272 N DEL 11
SRR1766451.3763295 chr19 20149956 N chr19 20150084 N DEL 10
SRR1766474.10888272 chr1 86111253 N chr1 86111373 N DEL 10
SRR1766450.8148628 chr1 86111297 N chr1 86111415 N DUP 10
SRR1766444.4894844 chr6 140064306 N chr6 140064407 N DEL 14
SRR1766449.9087558 chr9 107729048 N chr9 107729364 N DEL 10
SRR1766461.9693040 chr9 107729083 N chr9 107729399 N DEL 10
SRR1766450.6158500 chr19 14002209 N chr19 14002559 N DEL 16
SRR1766472.8993461 chr20 22762322 N chr20 22762437 N DEL 17
SRR1766477.4925378 chr10 100525781 N chr10 100525866 N DUP 18
SRR1766448.6033794 chrY 56832640 N chrY 56832691 N DEL 13
SRR1766442.38311926 chrY 56832624 N chrY 56832703 N DUP 11
SRR1766479.10093370 chrY 56832521 N chrY 56832689 N DEL 12
SRR1766442.31466519 chrY 56832624 N chrY 56832703 N DUP 13
SRR1766475.8007632 chrY 56832533 N chrY 56832646 N DEL 15
SRR1766466.2012533 chrY 56832479 N chrY 56832667 N DEL 10
SRR1766463.5068019 chrY 56832638 N chrY 56832694 N DEL 10
SRR1766475.2164559 chrY 56832624 N chrY 56832703 N DUP 11
SRR1766458.8372337 chrY 56832501 N chrY 56832672 N DUP 10
SRR1766462.9955769 chrY 56832526 N chrY 56832694 N DEL 15
SRR1766486.8525340 chrY 56832502 N chrY 56832658 N DUP 18
SRR1766463.6734647 chrY 56832526 N chrY 56832674 N DEL 15
SRR1766445.10308449 chrY 56832502 N chrY 56832688 N DUP 18
SRR1766483.9136165 chrY 56832521 N chrY 56832689 N DEL 10
SRR1766479.10303115 chrY 56832521 N chrY 56832689 N DEL 15
SRR1766484.11567279 chrY 56832536 N chrY 56832694 N DEL 10
SRR1766478.3691734 chrY 56832638 N chrY 56832694 N DEL 10
SRR1766442.45774751 chrY 56832497 N chrY 56832645 N DEL 10
SRR1766486.1471825 chrY 56832642 N chrY 56832693 N DEL 11
SRR1766466.7808909 chr4 117720751 N chr4 117720812 N DEL 10
SRR1766479.2587893 chr20 7435649 N chr20 7435727 N DUP 10
SRR1766483.4645820 chr20 7435646 N chr20 7435724 N DUP 10
SRR1766452.9837535 chr20 7435649 N chr20 7435727 N DUP 10
SRR1766457.9327095 chr20 7435649 N chr20 7435727 N DUP 10
SRR1766460.1446938 chr20 7435649 N chr20 7435727 N DUP 10
SRR1766470.1923036 chr20 7435646 N chr20 7435724 N DUP 11
SRR1766484.4910515 chr20 7435646 N chr20 7435724 N DUP 11
SRR1766483.10479412 chr20 7435649 N chr20 7435727 N DUP 14
SRR1766476.980463 chr20 7435646 N chr20 7435724 N DUP 15
SRR1766473.5591225 chr20 7435649 N chr20 7435727 N DUP 15
SRR1766450.3199741 chr20 7435564 N chr20 7435649 N DEL 11
SRR1766451.6086716 chr20 7435716 N chr20 7435799 N DUP 11
SRR1766464.10206603 chr20 7435716 N chr20 7435799 N DUP 14
SRR1766470.4212007 chr20 7435716 N chr20 7435799 N DUP 13
SRR1766456.5998792 chr20 7435716 N chr20 7435799 N DUP 14
SRR1766443.4427402 chr20 7435716 N chr20 7435799 N DUP 16
SRR1766467.9584497 chr20 7435666 N chr20 7435787 N DUP 11
SRR1766442.7553470 chr20 7435565 N chr20 7435691 N DEL 11
SRR1766472.4935429 chr20 7435564 N chr20 7435690 N DEL 12
SRR1766456.4351115 chr18 2503138 N chr18 2503241 N DUP 13
SRR1766465.2727385 chr18 2503137 N chr18 2503240 N DUP 14
SRR1766462.936562 chr18 2503140 N chr18 2503243 N DUP 11
SRR1766471.11903613 chr18 2503139 N chr18 2503242 N DUP 12
SRR1766479.8949503 chr3 129818550 N chr3 129818726 N DEL 10
SRR1766460.8110663 chr3 129818550 N chr3 129818726 N DEL 10
SRR1766455.1902287 chr3 129818550 N chr3 129818726 N DEL 14
SRR1766459.7798327 chr10 97528266 N chr10 97528713 N DUP 10
SRR1766474.9418331 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766478.10634670 chr10 97528269 N chr10 97528542 N DUP 12
SRR1766485.4316907 chr10 97528285 N chr10 97528462 N DEL 12
SRR1766482.8103838 chr10 97528318 N chr10 97528494 N DEL 10
SRR1766478.3385295 chr10 97528742 N chr10 97528891 N DEL 10
SRR1766471.10122187 chr10 97528266 N chr10 97528713 N DUP 10
SRR1766459.7798327 chr10 97528266 N chr10 97528713 N DUP 10
SRR1766447.6587341 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766466.4707542 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766442.21617368 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766446.5274089 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766453.7178381 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766459.544123 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766452.2676140 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766442.35961471 chr10 97528298 N chr10 97528747 N DEL 10
SRR1766454.2360020 chr10 97528776 N chr10 97528827 N DEL 11
SRR1766473.4108898 chr10 97528489 N chr10 97528861 N DEL 10
SRR1766450.2325619 chr10 97528330 N chr10 97529050 N DUP 11
SRR1766472.4878735 chr10 97528405 N chr10 97529250 N DUP 10
SRR1766470.10294740 chr3 184414636 N chr3 184414785 N DEL 12
SRR1766449.5866435 chr3 184414761 N chr3 184414915 N DEL 10
SRR1766472.4608855 chr3 184414961 N chr3 184415050 N DEL 13
SRR1766442.7352387 chr12 40773785 N chr12 40773846 N DEL 10
SRR1766472.7203057 chr12 40773785 N chr12 40773846 N DEL 14
SRR1766473.2772632 chr12 40773787 N chr12 40773848 N DEL 13
SRR1766452.5319159 chrX 532911 N chrX 533084 N DUP 10
SRR1766479.3812222 chrX 532911 N chrX 533084 N DUP 10
SRR1766459.8470207 chrX 532911 N chrX 533084 N DUP 10
SRR1766461.7756351 chrX 532911 N chrX 533084 N DUP 10
SRR1766461.7307005 chrX 532911 N chrX 533084 N DUP 10
SRR1766472.9522075 chrX 532910 N chrX 533083 N DUP 10
SRR1766455.2629016 chrX 532736 N chrX 532905 N DEL 18
SRR1766446.1965177 chrX 532736 N chrX 532905 N DEL 17
SRR1766458.1053295 chrX 532498 N chrX 532846 N DEL 13
SRR1766450.6752566 chrX 532358 N chrX 532698 N DUP 12
SRR1766484.10044483 chrX 532358 N chrX 532698 N DUP 12
SRR1766483.6348287 chrX 532358 N chrX 532698 N DUP 14
SRR1766470.10694971 chrX 532814 N chrX 532984 N DUP 11
SRR1766475.3914026 chrX 532334 N chrX 532836 N DUP 16
SRR1766471.7625282 chrX 532334 N chrX 532836 N DUP 16
SRR1766451.5814113 chrX 532334 N chrX 532836 N DUP 11
SRR1766455.1843895 chrX 532334 N chrX 532495 N DUP 10
SRR1766466.741586 chrX 532402 N chrX 533084 N DUP 15
SRR1766479.12130205 chrX 532334 N chrX 532489 N DUP 10
SRR1766482.3287684 chrX 532688 N chrX 532857 N DEL 10
SRR1766442.42037449 chrX 532402 N chrX 533084 N DUP 15
SRR1766451.2837471 chrX 532338 N chrX 532487 N DUP 10
SRR1766462.325216 chrX 532770 N chrX 532937 N DUP 10
SRR1766479.7259905 chrX 532910 N chrX 533083 N DUP 15
SRR1766485.8417833 chrX 532880 N chrX 533053 N DUP 15
SRR1766448.8150322 chrX 532911 N chrX 533084 N DUP 11
SRR1766483.8662027 chrX 532911 N chrX 533084 N DUP 10
SRR1766447.4543671 chrX 532911 N chrX 533084 N DUP 10
SRR1766481.6379179 chrX 532905 N chrX 533078 N DUP 15
SRR1766483.2085544 chrX 532905 N chrX 533078 N DUP 10
SRR1766442.45090361 chrX 532911 N chrX 533084 N DUP 15
SRR1766486.1970114 chrX 532911 N chrX 533084 N DUP 15
SRR1766463.5423529 chrX 532910 N chrX 533083 N DUP 15
SRR1766459.5797587 chrX 532911 N chrX 533084 N DUP 10
SRR1766452.2924394 chrX 532911 N chrX 533084 N DUP 10
SRR1766449.8737437 chrX 532477 N chrX 532816 N DEL 11
SRR1766455.7942497 chrX 532477 N chrX 532816 N DEL 11
SRR1766459.5079220 chrX 532477 N chrX 532816 N DEL 13
SRR1766484.10425771 chrX 532477 N chrX 532816 N DEL 18
SRR1766442.45639657 chrX 532911 N chrX 533084 N DUP 10
SRR1766460.2188702 chrX 532477 N chrX 532816 N DEL 18
SRR1766461.6522231 chrX 532911 N chrX 533084 N DUP 10
SRR1766470.6796442 chrX 532477 N chrX 532816 N DEL 18
SRR1766448.4524579 chrX 532814 N chrX 532987 N DUP 15
SRR1766454.3179782 chrX 532814 N chrX 532987 N DUP 15
SRR1766442.41208733 chrX 532813 N chrX 532988 N DEL 11
SRR1766471.4497294 chr7 4125056 N chr7 4125301 N DEL 14
SRR1766486.10138534 chr7 4125175 N chr7 4125538 N DEL 10
SRR1766476.11171341 chr7 4125034 N chr7 4125265 N DUP 10
SRR1766484.573583 chr7 4125023 N chr7 4125157 N DEL 10
SRR1766485.6945862 chr7 4125059 N chr7 4125493 N DEL 15
SRR1766460.2223474 chr7 4125055 N chr7 4125497 N DEL 11
SRR1766453.10211856 chr11 39227973 N chr11 39228088 N DEL 16
SRR1766469.10040682 chr11 39227973 N chr11 39228088 N DEL 17
SRR1766466.7695446 chr22 10851006 N chr22 10851403 N DEL 11
SRR1766457.8596287 chr22 10851006 N chr22 10851403 N DEL 11
SRR1766448.8537627 chr5 95927538 N chr5 95927687 N DEL 11
SRR1766482.5734359 chr5 95927538 N chr5 95927687 N DEL 12
SRR1766453.4684209 chr5 95927538 N chr5 95927687 N DEL 13
SRR1766473.2657398 chr5 95927538 N chr5 95927687 N DEL 14
SRR1766448.1948502 chr5 95927538 N chr5 95927687 N DEL 18
SRR1766456.4332329 chr5 95927538 N chr5 95927687 N DEL 18
SRR1766484.7202850 chr5 95927538 N chr5 95927687 N DEL 18
SRR1766453.9194829 chr5 95927538 N chr5 95927687 N DEL 18
SRR1766464.10687207 chr5 95927575 N chr5 95927626 N DEL 10
SRR1766450.3401078 chr5 95927602 N chr5 95927673 N DUP 14
SRR1766485.6700458 chr5 95927602 N chr5 95927673 N DUP 14
SRR1766450.907134 chr5 95927575 N chr5 95927626 N DEL 13
SRR1766479.10926599 chr5 95927575 N chr5 95927626 N DEL 13
SRR1766472.390523 chr5 95927538 N chr5 95927687 N DEL 17
SRR1766462.1362974 chr5 95927538 N chr5 95927687 N DEL 16
SRR1766448.8537627 chr5 95927723 N chr5 95927856 N DEL 14
SRR1766442.17561281 chr5 95927723 N chr5 95927856 N DEL 14
SRR1766442.42413776 chr5 95927723 N chr5 95927856 N DEL 14
SRR1766453.9194829 chr5 95927723 N chr5 95927856 N DEL 14
SRR1766474.3141017 chr5 95927599 N chr5 95927856 N DEL 14
SRR1766447.2933504 chr5 95927599 N chr5 95927856 N DEL 13
SRR1766449.4709640 chr5 95927599 N chr5 95927856 N DEL 10
SRR1766485.1385375 chr5 95927599 N chr5 95927886 N DEL 10
SRR1766442.39842660 chr5 95927599 N chr5 95927886 N DEL 13
SRR1766482.8962914 chr5 95927599 N chr5 95927886 N DEL 15
SRR1766457.1080109 chr5 95927854 N chr5 95927941 N DUP 15
SRR1766451.6600763 chr5 95927573 N chr5 95927886 N DEL 10
SRR1766442.10168482 chr13 27998912 N chr13 27999042 N DUP 14
SRR1766452.1060388 chr13 27998964 N chr13 27999037 N DUP 19
SRR1766464.3101435 chr13 27999088 N chr13 27999286 N DEL 11
SRR1766476.1476588 chr13 27998960 N chr13 27999064 N DUP 15
SRR1766486.2975113 chr13 27998960 N chr13 27999064 N DUP 18
SRR1766473.217054 chr13 27999047 N chr13 27999112 N DUP 14
SRR1766455.5249921 chr13 27999047 N chr13 27999112 N DUP 14
SRR1766445.7825528 chr13 27998984 N chr13 27999042 N DEL 14
SRR1766453.780664 chr13 27998960 N chr13 27999064 N DUP 19
SRR1766465.3351649 chr13 27999042 N chr13 27999107 N DUP 18
SRR1766453.2406926 chr13 27998967 N chr13 27999171 N DUP 17
SRR1766454.4206526 chr13 27998983 N chr13 27999041 N DEL 16
SRR1766485.427727 chr13 27998960 N chr13 27999174 N DUP 15
SRR1766462.2537060 chr13 27998964 N chr13 27999258 N DUP 19
SRR1766486.6316215 chr13 27998961 N chr13 27999127 N DUP 18
SRR1766445.1502972 chr13 27999109 N chr13 27999172 N DEL 16
SRR1766475.9643434 chr13 27999109 N chr13 27999172 N DEL 15
SRR1766482.8602446 chr13 27999093 N chr13 27999246 N DEL 15
SRR1766482.9737075 chr13 27999112 N chr13 27999286 N DEL 13
SRR1766448.6395271 chr13 27999093 N chr13 27999246 N DEL 16
SRR1766472.9208603 chr13 27999093 N chr13 27999246 N DEL 16
SRR1766442.33258567 chr13 27999305 N chr13 27999364 N DUP 13
SRR1766468.3392298 chr13 27999305 N chr13 27999364 N DUP 15
SRR1766465.3351649 chr13 27999292 N chr13 27999369 N DEL 14
SRR1766449.2341929 chr8 141107329 N chr8 141108064 N DEL 10
SRR1766466.3563887 chr8 141107366 N chr8 141107613 N DEL 10
SRR1766479.4036519 chr8 141107540 N chr8 141107949 N DEL 19
SRR1766479.503744 chr8 141107528 N chr8 141107801 N DUP 10
SRR1766462.4683611 chr8 141107467 N chr8 141107602 N DEL 10
SRR1766485.300084 chr8 141107639 N chr8 141107774 N DUP 17
SRR1766480.3151908 chr8 141107639 N chr8 141107828 N DUP 15
SRR1766453.9259003 chr8 141107639 N chr8 141107774 N DUP 17
SRR1766463.2999767 chr8 141107637 N chr8 141107774 N DEL 10
SRR1766465.2183344 chr14 94803992 N chr14 94804114 N DUP 12
SRR1766443.11202283 chr2 41747326 N chr2 41747782 N DEL 12
SRR1766473.7426786 chr2 41747326 N chr2 41747782 N DEL 17
SRR1766465.9079019 chr2 41747529 N chr2 41747708 N DEL 10
SRR1766468.1525396 chr2 41747930 N chr2 41748257 N DEL 10
SRR1766453.5686119 chr17 79555643 N chr17 79555708 N DUP 10
SRR1766468.1056974 chr17 79555761 N chr17 79555844 N DUP 10
SRR1766483.10739498 chr17 79555628 N chr17 79555761 N DEL 15
SRR1766442.40057164 chr17 79555688 N chr17 79555836 N DEL 15
SRR1766442.23473056 chr17 79555848 N chr17 79555939 N DEL 11
SRR1766478.6765001 chr22 44813507 N chr22 44813579 N DEL 18
SRR1766466.518549 chr22 44813507 N chr22 44813579 N DEL 18
SRR1766442.2530365 chr22 44813507 N chr22 44813579 N DEL 18
SRR1766443.1886040 chr22 44813507 N chr22 44813579 N DEL 18
SRR1766453.4508940 chr22 44813408 N chr22 44813579 N DEL 16
SRR1766451.2645951 chr22 44813408 N chr22 44813579 N DEL 15
SRR1766474.3387641 chr5 105934197 N chr5 105934254 N DEL 14
SRR1766479.1327134 chr5 105934197 N chr5 105934254 N DEL 14
SRR1766451.784357 chr5 105934197 N chr5 105934254 N DEL 13
SRR1766451.8174136 chr5 105934201 N chr5 105934254 N DEL 14
SRR1766471.10894678 chr22 16311144 N chr22 16311220 N DEL 10
SRR1766450.9270371 chr22 16311144 N chr22 16311220 N DEL 12
SRR1766442.13274391 chr22 16311116 N chr22 16311216 N DUP 13
SRR1766442.38890689 chr22 16311028 N chr22 16311130 N DEL 10
SRR1766456.557089 chr5 76812328 N chr5 76812562 N DEL 12
SRR1766480.7537691 chr14 103896736 N chr14 103896870 N DEL 12
SRR1766455.7545021 chr14 103896736 N chr14 103896870 N DEL 14
SRR1766456.3212529 chr14 103896736 N chr14 103896870 N DEL 14
SRR1766463.9267279 chr14 103896736 N chr14 103896870 N DEL 14
SRR1766475.8483473 chr14 103896777 N chr14 103896877 N DUP 10
SRR1766477.11111545 chr17 32027468 N chr17 32027703 N DEL 12
SRR1766449.10273736 chr17 32027499 N chr17 32027692 N DUP 16
SRR1766479.11758575 chr17 32027516 N chr17 32027665 N DEL 10
SRR1766458.5217232 chr1 27086744 N chr1 27087193 N DUP 11
SRR1766446.5051086 chr1 27086975 N chr1 27087122 N DEL 10
SRR1766481.2658246 chr10 127017056 N chr10 127017195 N DEL 13
SRR1766458.7463648 chr10 127017024 N chr10 127017217 N DUP 10
SRR1766480.4291630 chr10 127017135 N chr10 127017350 N DEL 12
SRR1766465.5244032 chr13 21187006 N chr13 21187161 N DUP 10
SRR1766464.6347688 chr13 21186961 N chr13 21187116 N DUP 13
SRR1766481.5743445 chrX 532910 N chrX 533083 N DUP 15
SRR1766479.7259905 chrX 532910 N chrX 533083 N DUP 15
SRR1766485.8417833 chrX 532880 N chrX 533053 N DUP 15
SRR1766448.8150322 chrX 532911 N chrX 533084 N DUP 14
SRR1766483.8662027 chrX 532911 N chrX 533084 N DUP 12
SRR1766455.8427191 chrX 532910 N chrX 533083 N DUP 10
SRR1766465.10786183 chrX 532905 N chrX 533078 N DUP 15
SRR1766447.4543671 chrX 532911 N chrX 533084 N DUP 10
SRR1766449.5255823 chrX 532905 N chrX 533078 N DUP 15
SRR1766481.6379179 chrX 532905 N chrX 533078 N DUP 15
SRR1766483.2085544 chrX 532905 N chrX 533078 N DUP 10
SRR1766442.45090361 chrX 532911 N chrX 533084 N DUP 15
SRR1766486.1970114 chrX 532911 N chrX 533084 N DUP 15
SRR1766463.5423529 chrX 532910 N chrX 533083 N DUP 15
SRR1766459.5797587 chrX 532911 N chrX 533084 N DUP 10
SRR1766452.2924394 chrX 532911 N chrX 533084 N DUP 10
SRR1766449.8737437 chrX 532832 N chrX 533002 N DUP 11
SRR1766455.7942497 chrX 532832 N chrX 533002 N DUP 11
SRR1766459.5079220 chrX 532832 N chrX 533002 N DUP 13
SRR1766484.10425771 chrX 532832 N chrX 533002 N DUP 18
SRR1766442.45639657 chrX 532911 N chrX 533084 N DUP 10
SRR1766460.2188702 chrX 532832 N chrX 533002 N DUP 18
SRR1766461.6522231 chrX 532911 N chrX 533084 N DUP 10
SRR1766470.6796442 chrX 532911 N chrX 533084 N DUP 10
SRR1766448.4524579 chrX 532832 N chrX 533005 N DUP 15
SRR1766454.3179782 chrX 532832 N chrX 533005 N DUP 15
SRR1766475.10489133 chr2 605329 N chr2 605558 N DUP 10
SRR1766476.6345955 chrX 140724592 N chrX 140724650 N DUP 17
SRR1766451.2489842 chrX 140724592 N chrX 140724656 N DUP 15
SRR1766454.3443467 chr10 132335439 N chr10 132335536 N DEL 10
SRR1766475.2115389 chr10 132335405 N chr10 132335596 N DUP 10
SRR1766447.9716661 chr6 31068343 N chr6 31068407 N DEL 14
SRR1766444.2088856 chr5 154652435 N chr5 154652756 N DEL 17
SRR1766465.9233155 chr6 112528600 N chr6 112528834 N DEL 10
SRR1766475.935907 chr16 46382002 N chr16 46382196 N DUP 11
SRR1766450.5351797 chr16 46382002 N chr16 46382222 N DUP 11
SRR1766445.10481479 chr16 46382002 N chr16 46382222 N DUP 12
SRR1766469.7048807 chr16 46382002 N chr16 46382222 N DUP 13
SRR1766463.2338987 chr16 46382130 N chr16 46382207 N DUP 14
SRR1766460.2705199 chr22 32564795 N chr22 32565128 N DEL 14
SRR1766482.7946696 chr22 32564795 N chr22 32565104 N DEL 15
SRR1766483.1025822 chr22 32564725 N chr22 32565032 N DUP 10
SRR1766451.9147954 chr22 32565043 N chr22 32565140 N DEL 18
SRR1766448.9008747 chr22 32564843 N chr22 32565054 N DUP 10
SRR1766442.22811814 chr22 32565026 N chr22 32565193 N DUP 15
SRR1766447.6659521 chr22 32565178 N chr22 32565299 N DEL 10
SRR1766443.3463904 chr22 32565178 N chr22 32565299 N DEL 10
SRR1766463.3201162 chr22 32564840 N chr22 32565195 N DUP 10
SRR1766462.6431756 chr22 32565188 N chr22 32565261 N DEL 10
SRR1766477.1060338 chr22 32564829 N chr22 32565234 N DEL 15
SRR1766442.20815922 chr22 32564750 N chr22 32565299 N DEL 10
SRR1766442.35126576 chr22 32565019 N chr22 32565332 N DEL 10
SRR1766477.11109204 chr5 120331265 N chr5 120331571 N DEL 10
SRR1766447.5881935 chr5 120331263 N chr5 120331571 N DEL 17
SRR1766448.8231890 chr5 120331265 N chr5 120331571 N DEL 13
SRR1766466.8467543 chr5 120331265 N chr5 120331571 N DEL 14
SRR1766446.1600829 chr5 120331266 N chr5 120331571 N DEL 15
SRR1766468.3080200 chr5 120331267 N chr5 120331571 N DEL 15
SRR1766483.7684297 chr22 31018598 N chr22 31018647 N DUP 10
SRR1766478.10808845 chr22 31018615 N chr22 31018770 N DUP 10
SRR1766450.6266288 chr8 144513900 N chr8 144513984 N DEL 10
SRR1766466.632635 chr8 144513900 N chr8 144513984 N DEL 11
SRR1766471.2806676 chr8 144513878 N chr8 144513960 N DUP 10
SRR1766455.3617250 chr4 20084508 N chr4 20084587 N DEL 10
SRR1766465.7761975 chr20 29231754 N chr20 29232439 N DEL 15
SRR1766447.4460022 chr21 46691879 N chr21 46692345 N DEL 15
SRR1766452.5364863 chr21 46691862 N chr21 46692069 N DUP 11
SRR1766462.5033484 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766442.27976247 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766442.47148570 chr21 46691947 N chr21 46692039 N DUP 11
SRR1766448.2550757 chr21 46692125 N chr21 46692589 N DEL 10
SRR1766454.3167232 chr21 46691995 N chr21 46692090 N DEL 15
SRR1766442.22852177 chr21 46692125 N chr21 46692589 N DEL 10
SRR1766458.5689457 chr21 46692159 N chr21 46692530 N DEL 13
SRR1766460.7883951 chr21 46692115 N chr21 46692207 N DUP 10
SRR1766483.1149532 chr21 46692159 N chr21 46692623 N DEL 10
SRR1766454.3140822 chr21 46692219 N chr21 46692590 N DEL 10
SRR1766454.1534689 chr21 46691940 N chr21 46692404 N DUP 10
SRR1766442.26888038 chr21 46692228 N chr21 46692506 N DEL 10
SRR1766451.2021055 chr21 46692228 N chr21 46692506 N DEL 10
SRR1766453.9792203 chr21 46691924 N chr21 46692204 N DEL 10
SRR1766482.6705002 chr21 46692219 N chr21 46692590 N DEL 15
SRR1766450.990571 chr21 46692228 N chr21 46692506 N DEL 10
SRR1766445.7257402 chr21 46692222 N chr21 46692684 N DUP 12
SRR1766474.9280975 chr21 46692039 N chr21 46692226 N DEL 15
SRR1766455.6462125 chr21 46691947 N chr21 46692132 N DUP 10
SRR1766442.6529872 chr21 46692321 N chr21 46692506 N DEL 10
SRR1766482.3990530 chr21 46692345 N chr21 46692530 N DEL 10
SRR1766445.8958413 chr21 46692033 N chr21 46692220 N DEL 10
SRR1766442.4205767 chr21 46692478 N chr21 46692665 N DEL 11
SRR1766450.3549229 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766476.8716028 chr21 46692345 N chr21 46692530 N DEL 11
SRR1766446.10311746 chr21 46692025 N chr21 46692489 N DEL 11
SRR1766457.2652553 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766442.3612491 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766445.9763279 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766458.7058430 chr21 46692318 N chr21 46692503 N DEL 15
SRR1766446.5267120 chr21 46692388 N chr21 46692573 N DEL 11
SRR1766473.3935525 chr21 46692579 N chr21 46692671 N DUP 12
SRR1766446.6766721 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766464.9797292 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766449.8392860 chr21 46692503 N chr21 46692595 N DUP 12
SRR1766460.10115496 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766466.10355654 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766481.7896101 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766458.5689457 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766454.3140822 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766461.5546154 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766452.2603472 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766470.4827682 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766464.6243082 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766471.1047566 chr21 46691941 N chr21 46692589 N DUP 10
SRR1766442.45738844 chr21 46692579 N chr21 46692671 N DUP 11
SRR1766442.8213125 chr21 46692579 N chr21 46692671 N DUP 15
SRR1766460.11257622 chr7 107679963 N chr7 107680055 N DEL 11
SRR1766466.5498767 chr6 16616704 N chr6 16616761 N DEL 11
SRR1766485.11596683 chr16 28442261 N chr16 28442472 N DEL 14
SRR1766475.7129747 chr2 4449607 N chr2 4449787 N DUP 14
SRR1766467.10393611 chr14 70477693 N chr14 70477774 N DUP 11
SRR1766463.6801109 chr20 61173334 N chr20 61173415 N DEL 10
SRR1766455.7617254 chr20 61173354 N chr20 61173415 N DEL 11
SRR1766457.6255076 chr8 67831217 N chr8 67831268 N DEL 17
SRR1766482.12785928 chr2 108765372 N chr2 108765560 N DUP 10
SRR1766468.3654191 chr2 108765585 N chr2 108765940 N DEL 15
SRR1766446.8711744 chr4 9981273 N chr4 9981489 N DEL 13
SRR1766463.689315 chr4 9981324 N chr4 9981419 N DUP 12
SRR1766442.35794695 chr4 9981324 N chr4 9981419 N DUP 15
SRR1766442.40441387 chr4 9981324 N chr4 9981419 N DUP 10
SRR1766463.7436736 chr4 9981355 N chr4 9981441 N DUP 10
SRR1766474.1433164 chr2 234899245 N chr2 234899296 N DEL 12
SRR1766475.6598973 chr2 234899245 N chr2 234899296 N DEL 13
SRR1766460.4989477 chr7 71592662 N chr7 71592716 N DEL 12
SRR1766450.6179352 chr2 239017444 N chr2 239018267 N DEL 10
SRR1766464.6106891 chr2 239017750 N chr2 239018267 N DEL 10
SRR1766444.6678286 chr2 239017965 N chr2 239018508 N DUP 12
SRR1766470.1261992 chr2 239018195 N chr2 239018298 N DEL 10
SRR1766462.521502 chr9 37918523 N chr9 37918584 N DEL 17
SRR1766480.6460053 chr9 37918523 N chr9 37918584 N DEL 17
SRR1766484.1566948 chr19 39153429 N chr19 39153611 N DUP 10
SRR1766468.3243441 chr19 39153429 N chr19 39153611 N DUP 15
SRR1766472.614869 chr19 39153429 N chr19 39153611 N DUP 15
SRR1766454.1822591 chr12 86502963 N chr12 86503678 N DEL 11
SRR1766451.747059 chr12 86502963 N chr12 86503678 N DEL 16
SRR1766452.10672015 chr12 86502936 N chr12 86503678 N DEL 16
SRR1766479.8499000 chr12 86502936 N chr12 86503678 N DEL 16
SRR1766483.12476605 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766458.1954919 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766475.8305492 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766470.2589770 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766476.3414480 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766486.5654796 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766443.2252384 chr12 86503218 N chr12 86503477 N DUP 10
SRR1766452.4805788 chr12 86503218 N chr12 86503623 N DUP 12
SRR1766447.4420733 chr12 86503218 N chr12 86503623 N DUP 12
SRR1766448.4502342 chr12 86503218 N chr12 86503623 N DUP 11
SRR1766483.7132869 chr12 86503218 N chr12 86503623 N DUP 11
SRR1766480.7626066 chr12 86503218 N chr12 86503623 N DUP 10
SRR1766465.4167578 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766470.8861870 chr12 86503583 N chr12 86503796 N DEL 14
SRR1766482.238544 chr12 86503583 N chr12 86503796 N DEL 12
SRR1766446.3770000 chr12 86503583 N chr12 86503796 N DEL 12
SRR1766464.689097 chr12 86503218 N chr12 86503623 N DUP 14
SRR1766450.8208644 chr12 86503015 N chr12 86503757 N DEL 13
SRR1766460.9088046 chr12 86503040 N chr12 86503784 N DEL 11
SRR1766476.1227802 chr12 86503452 N chr12 86503753 N DUP 11
SRR1766454.7315669 chr12 86503146 N chr12 86503480 N DEL 14
SRR1766445.10648095 chr12 86503015 N chr12 86503478 N DEL 16
SRR1766463.3142576 chr12 86503015 N chr12 86503478 N DEL 10
SRR1766472.11196187 chr12 86503583 N chr12 86503796 N DEL 11
SRR1766448.5492515 chr12 86503583 N chr12 86503796 N DEL 13
SRR1766450.5038210 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766469.3903658 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766479.5023210 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766452.5596729 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766445.3268784 chr12 86503040 N chr12 86503784 N DEL 12
SRR1766457.2510486 chr12 86503218 N chr12 86503623 N DUP 14
SRR1766447.10962633 chr12 86503173 N chr12 86503937 N DEL 17
SRR1766448.4914540 chr12 86503173 N chr12 86503937 N DEL 17
SRR1766475.8163142 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766442.36290555 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766475.5221749 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766479.8525665 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766480.7626066 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766458.6030704 chr12 86503000 N chr12 86503937 N DEL 19
SRR1766453.1978957 chr12 86502842 N chr12 86503937 N DEL 17
SRR1766473.6012036 chr12 86502842 N chr12 86503937 N DEL 17
SRR1766442.32326032 chr12 86502799 N chr12 86503940 N DEL 12
SRR1766474.10867554 chr12 86503002 N chr12 86503939 N DEL 13
SRR1766465.5883884 chr12 86502799 N chr12 86503940 N DEL 12
SRR1766443.1518904 chr5 1422508 N chr5 1422621 N DEL 14
SRR1766451.6565019 chr5 1422521 N chr5 1422598 N DEL 10
SRR1766453.4421351 chr5 1422521 N chr5 1422598 N DEL 10
SRR1766460.10481947 chr5 1422521 N chr5 1422598 N DEL 15
SRR1766446.7632159 chr5 1422521 N chr5 1422598 N DEL 10
SRR1766462.7793342 chr5 1422521 N chr5 1422598 N DEL 10
SRR1766467.4156380 chr5 1422929 N chr5 1423232 N DEL 14
SRR1766456.3987549 chr5 1422962 N chr5 1423037 N DEL 15
SRR1766452.8274267 chr5 1422659 N chr5 1423366 N DEL 15
SRR1766446.8387355 chr5 1422721 N chr5 1422904 N DEL 15
SRR1766459.11405611 chr5 1422743 N chr5 1422926 N DEL 10
SRR1766483.9581925 chr5 1422645 N chr5 1422904 N DEL 14
SRR1766451.6565019 chr5 1422598 N chr5 1422893 N DUP 17
SRR1766461.6318056 chr5 1422704 N chr5 1423187 N DEL 10
SRR1766450.2401568 chr5 1422710 N chr5 1423115 N DUP 13
SRR1766468.1017296 chr5 1422659 N chr5 1423366 N DEL 11
SRR1766467.7203391 chr5 1422686 N chr5 1422907 N DEL 18
SRR1766461.559133 chr5 1422993 N chr5 1423180 N DEL 18
SRR1766480.6248292 chr5 1422949 N chr5 1423250 N DEL 16
SRR1766458.4364186 chr5 1422887 N chr5 1423262 N DEL 10
SRR1766448.4973613 chr5 1422598 N chr5 1423345 N DEL 10
SRR1766481.8306630 chr5 1422881 N chr5 1423330 N DEL 10
SRR1766457.5667459 chr5 1422960 N chr5 1423345 N DEL 13
SRR1766473.8570077 chr5 1422960 N chr5 1423421 N DEL 17
SRR1766442.38880851 chr5 1422960 N chr5 1423421 N DEL 15
SRR1766485.2364021 chr7 79625289 N chr7 79625731 N DEL 19
SRR1766460.5126526 chr7 79625289 N chr7 79625731 N DEL 15
SRR1766480.2526661 chr7 79625289 N chr7 79625731 N DEL 13
SRR1766473.11175073 chr7 79625387 N chr7 79625546 N DUP 13
SRR1766442.12609679 chr7 79625272 N chr7 79625565 N DUP 13
SRR1766476.3754791 chr7 79625437 N chr7 79625575 N DEL 13
SRR1766443.6920293 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766457.7808506 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766474.7472757 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766463.5958978 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766474.259067 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766448.9678324 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766477.11399962 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766460.10637313 chr7 79625262 N chr7 79625577 N DEL 13
SRR1766457.3942266 chr7 79625263 N chr7 79625578 N DEL 12
SRR1766455.769442 chr7 79625404 N chr7 79625731 N DEL 17
SRR1766458.3622690 chr7 79625404 N chr7 79625731 N DEL 17
SRR1766485.3527106 chr7 79625267 N chr7 79625733 N DEL 13
SRR1766478.1821811 chr7 79625266 N chr7 79625732 N DEL 14
SRR1766476.8620447 chr2 195568522 N chr2 195568699 N DUP 13
SRR1766444.965161 chr2 195568522 N chr2 195568699 N DUP 11
SRR1766472.55170 chr9 65463290 N chr9 65463409 N DUP 10
SRR1766465.5267955 chr9 65463526 N chr9 65463585 N DUP 11
SRR1766486.191736 chr9 65463576 N chr9 65463822 N DEL 14
SRR1766450.29170 chr9 65463959 N chr9 65464078 N DEL 15
SRR1766445.4150389 chr9 65463966 N chr9 65464085 N DEL 11
SRR1766449.975507 chr9 65463462 N chr9 65463983 N DUP 10
SRR1766448.6874688 chr9 65464163 N chr9 65464342 N DEL 12
SRR1766469.2135139 chr9 65463591 N chr9 65464146 N DEL 10
SRR1766462.5534147 chr9 65463999 N chr9 65464232 N DUP 10
SRR1766461.7998064 chr9 65463964 N chr9 65464199 N DEL 10
SRR1766474.5992460 chr18 5307846 N chr18 5307991 N DUP 10
SRR1766482.12475002 chr18 5307846 N chr18 5307991 N DUP 10
SRR1766467.19534 chr18 5307846 N chr18 5307991 N DUP 10
SRR1766467.5165606 chr18 5307846 N chr18 5307991 N DUP 10
SRR1766468.6569986 chr18 5307864 N chr18 5307991 N DUP 13
SRR1766459.7245454 chr18 5307844 N chr18 5307899 N DEL 10
SRR1766457.7471719 chr18 5307846 N chr18 5307901 N DEL 10
SRR1766464.7261643 chr18 5307848 N chr18 5307903 N DEL 10
SRR1766442.7950695 chr7 153099455 N chr7 153099592 N DUP 14
SRR1766458.4748583 chr7 153099506 N chr7 153099610 N DUP 12
SRR1766477.10462747 chr7 153099506 N chr7 153099610 N DUP 19
SRR1766471.259 chr7 153099510 N chr7 153099581 N DEL 17
SRR1766473.4535927 chr7 153099510 N chr7 153099581 N DEL 17
SRR1766455.8674197 chr7 153099510 N chr7 153099581 N DEL 16
SRR1766465.7834250 chr7 153099477 N chr7 153099581 N DEL 10
SRR1766460.2375924 chr7 153099477 N chr7 153099581 N DEL 10
SRR1766460.1390015 chr12 130843991 N chr12 130844094 N DEL 14
SRR1766486.3970704 chr18 72700595 N chr18 72700674 N DEL 17
SRR1766474.2729783 chr18 72700593 N chr18 72700644 N DUP 13
SRR1766486.3837591 chr18 72700593 N chr18 72700644 N DUP 10
SRR1766486.8019183 chr18 72700585 N chr18 72700676 N DUP 17
SRR1766450.7661405 chr18 72700585 N chr18 72700676 N DUP 17
SRR1766475.3957081 chr18 72700595 N chr18 72700646 N DUP 10
SRR1766444.4425999 chr18 72700607 N chr18 72700728 N DUP 11
SRR1766458.6652782 chr18 72700607 N chr18 72700728 N DUP 14
SRR1766449.10167784 chr18 72700607 N chr18 72700728 N DUP 14
SRR1766452.3049058 chr18 72700607 N chr18 72700728 N DUP 14
SRR1766455.8822209 chr18 72700607 N chr18 72700728 N DUP 14
SRR1766482.6669758 chr18 72700714 N chr18 72700779 N DEL 17
SRR1766486.11203849 chr18 72700660 N chr18 72700717 N DEL 12
SRR1766458.8526070 chr18 72700723 N chr18 72700812 N DUP 11
SRR1766452.9140727 chr18 72700723 N chr18 72700802 N DUP 18
SRR1766447.1653752 chr18 72700586 N chr18 72700689 N DEL 16
SRR1766455.4383246 chr18 72700586 N chr18 72700689 N DEL 15
SRR1766456.2661636 chr18 72700679 N chr18 72700800 N DUP 14
SRR1766455.451742 chr18 72700717 N chr18 72700808 N DUP 16
SRR1766452.7514105 chr18 72700609 N chr18 72700806 N DUP 10
SRR1766477.8502443 chr18 72700688 N chr18 72700759 N DUP 16
SRR1766442.12898108 chr18 72700569 N chr18 72700820 N DUP 10
SRR1766448.1798010 chr18 72700638 N chr18 72700839 N DUP 15
SRR1766480.7812158 chr18 72700739 N chr18 72700846 N DUP 19
SRR1766460.4303843 chr18 72700713 N chr18 72700768 N DUP 18
SRR1766442.44724368 chr18 72700791 N chr18 72700854 N DEL 14
SRR1766455.9733843 chr18 72700791 N chr18 72700854 N DEL 15
SRR1766466.1964496 chr18 72700724 N chr18 72700779 N DEL 10
SRR1766463.2524836 chr18 72700698 N chr18 72700785 N DEL 11
SRR1766486.8019183 chr18 72700698 N chr18 72700785 N DEL 11
SRR1766474.2729783 chr18 72700648 N chr18 72700837 N DEL 16
SRR1766442.25737276 chr18 72700752 N chr18 72700851 N DEL 14
SRR1766481.3362828 chr18 72700752 N chr18 72700851 N DEL 14
SRR1766450.3832692 chr4 113340843 N chr4 113340998 N DEL 12
SRR1766468.5266684 chr4 113340858 N chr4 113340998 N DEL 10
SRR1766442.31217042 chr18 56600456 N chr18 56600729 N DEL 12
SRR1766466.8081937 chr18 56600477 N chr18 56600750 N DEL 10
SRR1766482.3069028 chr18 56600477 N chr18 56600682 N DEL 12
SRR1766463.5474017 chr18 56600456 N chr18 56600729 N DEL 10
SRR1766468.2214364 chr13 112913096 N chr13 112913290 N DEL 16
SRR1766482.1615913 chr13 112912925 N chr13 112913136 N DUP 10
SRR1766485.1254717 chr13 112912925 N chr13 112913136 N DUP 10
SRR1766468.1245468 chr13 112913196 N chr13 112913485 N DUP 13
SRR1766442.21004947 chr13 112913230 N chr13 112913441 N DUP 12
SRR1766477.11772392 chr13 112913030 N chr13 112913230 N DEL 10
SRR1766478.4786746 chr13 112912940 N chr13 112913261 N DEL 10
SRR1766472.1862328 chrX 2478837 N chrX 2479035 N DUP 10
SRR1766466.6429593 chrX 2479502 N chrX 2479824 N DEL 10
SRR1766467.372297 chrX 2479508 N chrX 2479830 N DEL 15
SRR1766474.4875424 chr1 4332511 N chr1 4332570 N DEL 10
SRR1766485.7883323 chr1 4332511 N chr1 4332570 N DEL 10
SRR1766471.1229517 chr1 4332511 N chr1 4332570 N DEL 17
SRR1766447.2595331 chr1 4332511 N chr1 4332570 N DEL 19
SRR1766471.6661709 chr1 4332511 N chr1 4332570 N DEL 10
SRR1766483.8087285 chr1 4332556 N chr1 4333518 N DEL 16
SRR1766465.10568007 chr1 4332511 N chr1 4332918 N DEL 15
SRR1766478.7511124 chr1 4332511 N chr1 4332570 N DEL 10
SRR1766454.9133928 chr1 4332614 N chr1 4333427 N DUP 10
SRR1766443.11094727 chr1 4332570 N chr1 4332627 N DUP 15
SRR1766479.12282309 chr1 4332511 N chr1 4332570 N DEL 12
SRR1766466.3535845 chr1 4332690 N chr1 4332777 N DEL 13
SRR1766462.4078557 chr1 4332645 N chr1 4332936 N DEL 10
SRR1766449.3611427 chr1 4332615 N chr1 4332991 N DUP 11
SRR1766478.828829 chr1 4332671 N chr1 4333517 N DEL 14
SRR1766485.2259402 chr1 4332570 N chr1 4332627 N DUP 10
SRR1766456.2953573 chr1 4332614 N chr1 4333048 N DUP 10
SRR1766471.1229517 chr1 4332614 N chr1 4332990 N DUP 10
SRR1766448.9216519 chr1 4332743 N chr1 4332976 N DEL 10
SRR1766460.5584371 chr1 4332700 N chr1 4333194 N DEL 10
SRR1766464.1642681 chr1 4333001 N chr1 4333584 N DUP 10
SRR1766463.8403608 chr1 4332614 N chr1 4333576 N DEL 10
SRR1766450.2795016 chr1 4333020 N chr1 4333489 N DEL 15
SRR1766459.7560099 chr1 4333049 N chr1 4333371 N DEL 10
SRR1766444.5549244 chr1 4333240 N chr1 4333448 N DEL 10
SRR1766443.2989947 chr1 4333182 N chr1 4333448 N DEL 10
SRR1766465.7261728 chr1 4332556 N chr1 4333460 N DEL 10
SRR1766454.10890745 chr1 4333054 N chr1 4333523 N DEL 10
SRR1766479.6270613 chr1 4333021 N chr1 4333575 N DUP 15
SRR1766484.9888651 chr1 4332515 N chr1 4333448 N DEL 15
SRR1766448.1485734 chr1 4332565 N chr1 4333146 N DEL 10
SRR1766472.7361104 chr1 4332631 N chr1 4333448 N DEL 12
SRR1766486.5451510 chr1 4332936 N chr1 4333167 N DUP 15
SRR1766444.2797920 chr1 4333112 N chr1 4333256 N DUP 10
SRR1766470.9585706 chr1 4332614 N chr1 4333108 N DEL 10
SRR1766472.10639638 chr1 4333133 N chr1 4333457 N DEL 10
SRR1766466.6107027 chr1 4332562 N chr1 4333085 N DEL 10
SRR1766474.1894881 chr1 4332556 N chr1 4333137 N DEL 10
SRR1766466.10153244 chr1 4332642 N chr1 4333136 N DEL 12
SRR1766467.849919 chr1 4333166 N chr1 4333310 N DUP 10
SRR1766464.5114633 chr1 4333053 N chr1 4333141 N DEL 12
SRR1766467.1043592 chr1 4333053 N chr1 4333493 N DEL 12
SRR1766442.32457730 chr1 4332614 N chr1 4333222 N DUP 10
SRR1766459.7560099 chr1 4332590 N chr1 4333169 N DUP 10
SRR1766481.11062883 chr1 4332590 N chr1 4333169 N DUP 10
SRR1766442.16313221 chr1 4332502 N chr1 4333226 N DUP 10
SRR1766462.1269920 chr1 4332560 N chr1 4333170 N DEL 10
SRR1766471.1038908 chr1 4333252 N chr1 4333489 N DEL 10
SRR1766469.3524751 chr1 4333066 N chr1 4333359 N DEL 10
SRR1766449.8726051 chr1 4333252 N chr1 4333489 N DEL 10
SRR1766466.3741585 chr1 4333223 N chr1 4333489 N DEL 10
SRR1766481.3825966 chr1 4333240 N chr1 4333448 N DEL 10
SRR1766450.792823 chr1 4333085 N chr1 4333229 N DUP 10
SRR1766442.20683542 chr1 4332560 N chr1 4333170 N DEL 10
SRR1766483.11597062 chr1 4332992 N chr1 4333165 N DUP 10
SRR1766483.8250848 chr1 4333228 N chr1 4333285 N DUP 10
SRR1766469.8345969 chr1 4333223 N chr1 4333489 N DEL 10
SRR1766458.7649016 chr1 4333049 N chr1 4333371 N DEL 10
SRR1766469.677256 chr1 4332555 N chr1 4333604 N DEL 10
SRR1766483.7481342 chr1 4333169 N chr1 4333493 N DEL 10
SRR1766442.8407769 chr1 4333240 N chr1 4333359 N DEL 10
SRR1766464.5741593 chr1 4333285 N chr1 4333464 N DEL 12
SRR1766442.34375501 chr1 4333053 N chr1 4333464 N DEL 14
SRR1766442.46233639 chr1 4333227 N chr1 4333433 N DEL 10
SRR1766443.3753855 chr1 4332564 N chr1 4333468 N DEL 12
SRR1766467.9049772 chr1 4333326 N chr1 4333447 N DEL 12
SRR1766485.286538 chr1 4332564 N chr1 4333468 N DEL 12
SRR1766474.7774313 chr1 4333136 N chr1 4333489 N DEL 10
SRR1766466.10153244 chr1 4332642 N chr1 4333136 N DEL 15
SRR1766478.4413525 chr1 4332502 N chr1 4333255 N DUP 10
SRR1766466.3741585 chr1 4332875 N chr1 4333489 N DEL 10
SRR1766450.2510119 chr1 4333136 N chr1 4333489 N DEL 10
SRR1766473.3704186 chr1 4332614 N chr1 4333545 N DUP 10
SRR1766481.12841215 chr1 4332874 N chr1 4333459 N DEL 15
SRR1766465.2185972 chr1 4332562 N chr1 4333085 N DEL 10
SRR1766479.6994666 chr1 4333053 N chr1 4333522 N DEL 10
SRR1766447.620163 chr1 4333240 N chr1 4333448 N DEL 10
SRR1766447.2251398 chr1 4333090 N chr1 4333731 N DUP 10
SRR1766480.8000657 chr1 4332874 N chr1 4333517 N DEL 10
SRR1766465.2185972 chr1 4333078 N chr1 4333489 N DEL 10
SRR1766467.9049772 chr1 4333547 N chr1 4333691 N DUP 10
SRR1766481.6779784 chr1 4333092 N chr1 4333588 N DUP 10
SRR1766465.7261728 chr1 4333371 N chr1 4333575 N DUP 10
SRR1766483.4148876 chr1 4333166 N chr1 4333575 N DUP 12
SRR1766479.2559879 chr1 4332879 N chr1 4333493 N DEL 10
SRR1766465.5208960 chr1 4332544 N chr1 4333448 N DEL 10
SRR1766455.346619 chr1 4333053 N chr1 4333522 N DEL 10
SRR1766458.7629482 chr1 4333460 N chr1 4333575 N DUP 10
SRR1766469.10592314 chr1 4333371 N chr1 4333575 N DUP 10
SRR1766474.8228594 chr1 4332999 N chr1 4333172 N DUP 10
SRR1766482.1670418 chr1 4332544 N chr1 4333448 N DEL 10
SRR1766449.1687719 chr1 4333310 N chr1 4333460 N DEL 15
SRR1766484.3692511 chr1 4333170 N chr1 4333579 N DUP 10
SRR1766468.4864345 chr1 4332875 N chr1 4333576 N DEL 10
SRR1766474.670863 chr1 4332556 N chr1 4333460 N DEL 10
SRR1766465.9274606 chr1 4332560 N chr1 4333170 N DEL 10
SRR1766458.7629482 chr1 4332556 N chr1 4333460 N DEL 10
SRR1766484.4761812 chr1 4333048 N chr1 4333604 N DEL 10
SRR1766442.43738499 chr1 4333048 N chr1 4333604 N DEL 10
SRR1766444.1054712 chr1 4332556 N chr1 4333460 N DEL 10
SRR1766454.10890745 chr1 4333053 N chr1 4333141 N DEL 15
SRR1766462.8971630 chr20 39587209 N chr20 39587258 N DUP 13
SRR1766457.4544417 chr20 39587209 N chr20 39587258 N DUP 16
SRR1766468.154946 chr2 16394934 N chr2 16395048 N DEL 11
SRR1766472.3984521 chr16 30168723 N chr16 30168880 N DEL 12
SRR1766454.8041988 chr1 240562858 N chr1 240563056 N DUP 17
SRR1766468.7033252 chr1 240562859 N chr1 240563099 N DUP 10
SRR1766466.8439118 chr1 240562859 N chr1 240563115 N DUP 16
SRR1766468.4875062 chr1 240563121 N chr1 240563285 N DEL 15
SRR1766458.7703655 chr1 240562882 N chr1 240563235 N DEL 15
SRR1766453.912378 chr1 240562873 N chr1 240563318 N DEL 11
SRR1766446.2314478 chr5 2082060 N chr5 2082754 N DEL 10
SRR1766476.5724190 chr5 2082097 N chr5 2082350 N DEL 10
SRR1766465.9617330 chr5 2082132 N chr5 2082196 N DEL 15
SRR1766451.2121864 chr5 2082182 N chr5 2082750 N DEL 10
SRR1766454.1259899 chr5 2082132 N chr5 2082196 N DEL 10
SRR1766453.6838218 chr5 2082191 N chr5 2082255 N DEL 10
SRR1766472.11871052 chr5 2082196 N chr5 2082258 N DUP 10
SRR1766456.182501 chr5 2082197 N chr5 2082385 N DUP 11
SRR1766443.1616175 chr5 2082209 N chr5 2082964 N DUP 16
SRR1766469.5317302 chr5 2082227 N chr5 2082478 N DUP 10
SRR1766481.1004632 chr5 2082250 N chr5 2082879 N DUP 10
SRR1766459.5443341 chr5 2082209 N chr5 2082964 N DUP 10
SRR1766450.5480536 chr5 2082209 N chr5 2082964 N DUP 12
SRR1766481.11384315 chr5 2082161 N chr5 2082286 N DUP 10
SRR1766475.6634289 chr5 2082209 N chr5 2082964 N DUP 10
SRR1766450.5453203 chr5 2082308 N chr5 2082750 N DEL 10
SRR1766475.6634289 chr5 2082227 N chr5 2082478 N DUP 10
SRR1766477.11119298 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766444.3096530 chr5 2082164 N chr5 2082352 N DUP 10
SRR1766453.3350555 chr5 2082196 N chr5 2082447 N DUP 10
SRR1766477.11550512 chr5 2082227 N chr5 2082478 N DUP 10
SRR1766442.22977030 chr5 2082227 N chr5 2082478 N DUP 15
SRR1766469.5618666 chr5 2082350 N chr5 2082475 N DUP 10
SRR1766470.6372347 chr5 2082075 N chr5 2082263 N DUP 13
SRR1766453.3543145 chr5 2082192 N chr5 2082254 N DUP 10
SRR1766485.4625684 chr5 2082136 N chr5 2082200 N DEL 10
SRR1766474.531252 chr5 2082209 N chr5 2082964 N DUP 13
SRR1766485.8949923 chr5 2082447 N chr5 2082700 N DEL 15
SRR1766450.5255427 chr5 2082196 N chr5 2082384 N DUP 11
SRR1766442.36890550 chr5 2082291 N chr5 2082733 N DEL 10
SRR1766461.9669304 chr5 2082731 N chr5 2082793 N DUP 10
SRR1766465.4384166 chr5 2082226 N chr5 2082353 N DEL 10
SRR1766467.11307747 chr5 2082316 N chr5 2082821 N DEL 10
SRR1766455.148065 chr5 2082190 N chr5 2082821 N DEL 15
SRR1766442.25830866 chr5 2082316 N chr5 2082821 N DEL 18
SRR1766468.1486245 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766457.7798515 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766442.35123216 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766456.2077572 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766478.10028038 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766481.6592463 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766453.9884496 chr5 2082196 N chr5 2082888 N DUP 10
SRR1766461.5710385 chr5 2082338 N chr5 2082906 N DEL 15
SRR1766486.2088918 chr5 2082317 N chr5 2082885 N DEL 10
SRR1766446.2988791 chr5 2082906 N chr5 2082968 N DUP 10
SRR1766458.9252244 chr5 2082906 N chr5 2082968 N DUP 18
SRR1766471.8172915 chr5 2082474 N chr5 2082916 N DEL 10
SRR1766447.4250475 chr7 132646995 N chr7 132647208 N DUP 10
SRR1766442.37684280 chr12 82640372 N chr12 82640563 N DEL 14
SRR1766461.10673178 chr12 82639946 N chr12 82640282 N DEL 16
SRR1766457.3600 chr12 82639946 N chr12 82640282 N DEL 15
SRR1766454.7802014 chr12 82640266 N chr12 82640401 N DUP 13
SRR1766462.8806091 chr4 38880239 N chr4 38880295 N DEL 18
SRR1766456.5791334 chr1 169273385 N chr1 169273788 N DEL 14
SRR1766454.7421730 chr1 169273377 N chr1 169273780 N DEL 10
SRR1766466.8733007 chr5 144847782 N chr5 144848047 N DEL 10
SRR1766479.11080116 chr12 110867472 N chr12 110867649 N DEL 10
SRR1766442.25827805 chr12 110867120 N chr12 110867747 N DUP 11
SRR1766486.5346696 chr12 110867266 N chr12 110867494 N DEL 10
SRR1766480.6170934 chr12 110867266 N chr12 110867494 N DEL 10
SRR1766475.6125733 chr12 110867109 N chr12 110867562 N DEL 10
SRR1766486.7937904 chr3 198076499 N chr3 198076566 N DEL 15
SRR1766486.695665 chr4 36484994 N chr4 36485105 N DEL 19
SRR1766469.7818746 chr4 36484995 N chr4 36485106 N DEL 14
SRR1766443.2206782 chr2 164818738 N chr2 164818797 N DEL 10
SRR1766467.3610157 chr12 130055314 N chr12 130055455 N DEL 10
SRR1766455.5570942 chr12 130055276 N chr12 130055438 N DEL 10
SRR1766467.739141 chr12 130055532 N chr12 130055663 N DUP 13
SRR1766459.4947587 chr16 22939832 N chr16 22939986 N DEL 15
SRR1766471.9068161 chr16 22939832 N chr16 22939986 N DEL 15
SRR1766485.4627710 chr16 22939878 N chr16 22940083 N DEL 14
SRR1766467.1384458 chr16 22939939 N chr16 22940042 N DEL 10
SRR1766457.6908869 chr16 22939832 N chr16 22939986 N DEL 10
SRR1766466.8348564 chr16 22939832 N chr16 22939986 N DEL 10
SRR1766443.1096478 chr16 22940075 N chr16 22940176 N DUP 10
SRR1766445.3124665 chr16 22939981 N chr16 22940339 N DEL 10
SRR1766486.8558441 chr16 22940059 N chr16 22940417 N DEL 10
SRR1766443.7356166 chr16 22939859 N chr16 22940472 N DEL 10
SRR1766475.7297021 chr2 203067146 N chr2 203067218 N DEL 12
SRR1766485.43942 chr14 85847716 N chr14 85847797 N DEL 17
SRR1766452.5001147 chr14 85847716 N chr14 85847797 N DEL 17
SRR1766452.6262241 chr14 85847716 N chr14 85847797 N DEL 17
SRR1766448.8686377 chr14 85847842 N chr14 85848173 N DEL 14
SRR1766475.513567 chr14 85847980 N chr14 85848239 N DEL 11
SRR1766468.5553988 chr14 85847980 N chr14 85848239 N DEL 13
SRR1766456.615286 chr14 85847948 N chr14 85848239 N DEL 14
SRR1766460.9172 chr14 85847948 N chr14 85848239 N DEL 14
SRR1766486.4783513 chr14 85847948 N chr14 85848239 N DEL 14
SRR1766479.8146751 chr14 85847916 N chr14 85848239 N DEL 14
SRR1766459.10919837 chr14 85847850 N chr14 85848239 N DEL 14
SRR1766461.4501618 chr14 85847850 N chr14 85848239 N DEL 14
SRR1766445.6889230 chr16 88798349 N chr16 88798495 N DUP 10
SRR1766446.5048959 chr7 56758269 N chr7 56758328 N DUP 10
SRR1766473.8006928 chrX 41507258 N chrX 41507388 N DUP 19
SRR1766459.3109839 chr18 41577578 N chr18 41577669 N DUP 17
SRR1766448.356980 chr1 191089495 N chr1 191089549 N DEL 10
SRR1766465.9799946 chr8 142991129 N chr8 142991326 N DEL 13
SRR1766451.1754076 chr17 83172625 N chr17 83172776 N DEL 10
SRR1766452.4099532 chr17 83172538 N chr17 83172725 N DUP 15
SRR1766445.132210 chr17 83172598 N chr17 83172749 N DEL 10
SRR1766486.3638211 chr17 83172560 N chr17 83172749 N DEL 13
SRR1766443.5260056 chr17 83172788 N chr17 83172863 N DUP 10
SRR1766481.8658521 chr17 83172625 N chr17 83172776 N DEL 10
SRR1766482.8305591 chr17 83172784 N chr17 83173538 N DUP 11
SRR1766474.8876135 chr17 83173214 N chr17 83173669 N DEL 19
SRR1766485.329596 chr17 83172521 N chr17 83172860 N DUP 14
SRR1766472.9689428 chr17 83172619 N chr17 83172694 N DUP 19
SRR1766442.30436134 chr17 83172580 N chr17 83173069 N DEL 16
SRR1766463.8855270 chr10 46136056 N chr10 46136105 N DUP 10
SRR1766452.2129119 chr10 46136056 N chr10 46136105 N DUP 12
SRR1766455.4201587 chr10 46136103 N chr10 46136168 N DEL 15
SRR1766455.1355315 chr10 46136090 N chr10 46136153 N DEL 11
SRR1766463.5064477 chr10 46136090 N chr10 46136153 N DEL 13
SRR1766470.1464109 chr10 46136090 N chr10 46136153 N DEL 13
SRR1766451.2805452 chr10 46136131 N chr10 46136200 N DUP 11
SRR1766465.9136980 chr10 46136136 N chr10 46136205 N DUP 16
SRR1766471.10465404 chr13 18944211 N chr13 18944429 N DEL 10
SRR1766485.5811589 chr2 129735720 N chr2 129735994 N DUP 13
SRR1766483.5615626 chr5 175051170 N chr5 175051227 N DEL 12
SRR1766452.9684565 chr4 6660611 N chr4 6660937 N DEL 14
SRR1766473.2455928 chr9 65825571 N chr9 65825760 N DEL 13
SRR1766481.8013694 chr9 65825571 N chr9 65825760 N DEL 18
SRR1766470.1526337 chr17 79827460 N chr17 79827583 N DEL 12
SRR1766477.6147934 chr17 79827460 N chr17 79827583 N DEL 12
SRR1766454.10340797 chr16 89196426 N chr16 89196613 N DEL 10
SRR1766474.4587026 chr14 48710863 N chr14 48710946 N DEL 11
SRR1766483.6730716 chr14 48710845 N chr14 48710959 N DEL 19
SRR1766484.3931912 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766462.3532246 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766470.3292467 chr14 48710863 N chr14 48710946 N DEL 11
SRR1766463.5167162 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766484.11328190 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766445.5006 chr14 48710815 N chr14 48710876 N DUP 12
SRR1766481.2252587 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766448.3439606 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766476.7842206 chr14 48710753 N chr14 48710904 N DUP 19
SRR1766457.4773511 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766442.36294710 chr14 48710753 N chr14 48710904 N DUP 19
SRR1766457.4441503 chr14 48710863 N chr14 48710946 N DEL 11
SRR1766472.5072988 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766479.13419391 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766470.5542698 chr14 48710815 N chr14 48710876 N DUP 19
SRR1766476.5459174 chr14 48710753 N chr14 48710904 N DUP 19
SRR1766448.3881858 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766468.4399353 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766478.689995 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766445.4807957 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766471.7338370 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766463.5102635 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766482.383305 chr14 48710815 N chr14 48710876 N DUP 16
SRR1766471.6801776 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766475.11458987 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766466.11132086 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766468.719585 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766457.2583891 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766448.974867 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766442.14276195 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766454.1977085 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766461.7484242 chr14 48710815 N chr14 48710876 N DUP 10
SRR1766475.496564 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766479.2762163 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766457.5768050 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766448.5798599 chr14 48710753 N chr14 48710904 N DUP 12
SRR1766484.1647397 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766442.17306690 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766479.7892122 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766472.187545 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766467.3508269 chr14 48710753 N chr14 48710904 N DUP 19
SRR1766442.26609313 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766467.5431639 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766446.3022653 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766442.38357669 chr14 48710753 N chr14 48710811 N DUP 19
SRR1766470.5233128 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766470.1748001 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766458.4095278 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766467.5431639 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766481.9557509 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766457.2534100 chr14 48710757 N chr14 48710818 N DUP 11
SRR1766469.531006 chr14 48710782 N chr14 48710840 N DUP 10
SRR1766473.5600841 chr14 48710783 N chr14 48710959 N DEL 15
SRR1766449.6067038 chr4 48104431 N chr4 48104684 N DEL 16
SRR1766466.8418436 chr4 48104421 N chr4 48104514 N DEL 18
SRR1766464.5030637 chr4 48104368 N chr4 48104462 N DUP 11
SRR1766448.7504018 chr4 48104464 N chr4 48104691 N DEL 17
SRR1766456.6177428 chr4 48104356 N chr4 48104442 N DUP 18
SRR1766450.6373742 chr4 48104464 N chr4 48104691 N DEL 19
SRR1766450.9514644 chr4 48104367 N chr4 48104632 N DUP 14
SRR1766452.4658940 chr4 48104365 N chr4 48104651 N DUP 13
SRR1766478.2343450 chr4 48104365 N chr4 48104651 N DUP 18
SRR1766445.4609705 chr4 48104383 N chr4 48104518 N DUP 12
SRR1766482.7192643 chr4 48104638 N chr4 48104715 N DUP 10
SRR1766482.3702258 chr4 48104403 N chr4 48104702 N DEL 15
SRR1766482.3483891 chr4 48104436 N chr4 48104691 N DEL 14
SRR1766477.6422413 chr4 48104399 N chr4 48104693 N DEL 11
SRR1766442.24635555 chr4 48104403 N chr4 48104702 N DEL 17
SRR1766468.5239912 chr4 48104403 N chr4 48104702 N DEL 17
SRR1766481.13074124 chr4 48104406 N chr4 48104705 N DEL 12
SRR1766463.9799838 chr4 48104408 N chr4 48104707 N DEL 10
SRR1766461.8010174 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766449.134392 chr17 77562775 N chr17 77562882 N DEL 18
SRR1766453.1980992 chr17 77562776 N chr17 77562934 N DUP 10
SRR1766449.2517215 chr17 77562775 N chr17 77562882 N DEL 16
SRR1766463.9843627 chr17 77562763 N chr17 77562870 N DEL 10
SRR1766480.7103607 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766481.4453507 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766470.2058659 chr17 77562769 N chr17 77562876 N DEL 10
SRR1766464.9796395 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766477.2284814 chr17 77562763 N chr17 77562870 N DEL 10
SRR1766448.4375654 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766477.5833728 chrY 11027124 N chrY 11027215 N DEL 11
SRR1766475.383348 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766454.9040902 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766484.5579563 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766443.7825574 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766484.1915601 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766450.8357767 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766480.6669082 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766442.4901217 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766446.4301961 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766486.2854498 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766484.4024732 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766482.3149900 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766455.1044501 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766474.2176121 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766482.6394426 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766447.8510608 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766477.1943205 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766442.38150251 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766454.1763559 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766454.6799396 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766452.8968949 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766484.1915601 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766446.9023220 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766442.9013655 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766467.9667718 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766453.10777787 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766477.4797036 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766482.282476 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766461.8985552 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766463.1766339 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766459.165027 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766442.28691290 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766475.1115337 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766451.9399581 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766450.1020368 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766456.6118378 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766442.8908181 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766457.3041478 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766474.8798753 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766460.6682335 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766473.5338326 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766481.2458626 chr6 106542759 N chr6 106543134 N DEL 10
SRR1766443.1400077 chr6 106542760 N chr6 106543135 N DEL 10
SRR1766483.9491190 chr2 57548080 N chr2 57548145 N DUP 11
SRR1766448.6682300 chr2 57548108 N chr2 57548161 N DEL 17
SRR1766454.6806192 chrX 136451176 N chrX 136451305 N DUP 19
SRR1766458.8746635 chrX 136451149 N chrX 136451220 N DEL 14
SRR1766464.8944529 chrX 136451220 N chrX 136451269 N DUP 19
SRR1766443.1096536 chrX 136451149 N chrX 136451220 N DEL 14
SRR1766449.7977451 chrX 136451114 N chrX 136451303 N DUP 18
SRR1766461.361617 chrX 136451222 N chrX 136451295 N DUP 12
SRR1766455.7313870 chrX 136451258 N chrX 136451319 N DUP 13
SRR1766442.43014644 chrX 136451145 N chrX 136451256 N DEL 18
SRR1766472.8105755 chrX 136451145 N chrX 136451256 N DEL 17
SRR1766456.952375 chrX 136451145 N chrX 136451256 N DEL 16
SRR1766463.7868411 chr5 180297014 N chr5 180297105 N DEL 19
SRR1766449.7751472 chr1 143258312 N chr1 143258458 N DUP 12
SRR1766475.10773090 chr16 7229895 N chr16 7230004 N DEL 13
SRR1766475.306879 chr14 89567556 N chr14 89567720 N DUP 13
SRR1766442.43901911 chr6 22836799 N chr6 22836928 N DEL 10
SRR1766457.769618 chr6 22837027 N chr6 22837377 N DEL 10
SRR1766474.6762309 chr6 22836737 N chr6 22837089 N DUP 10
SRR1766473.7352866 chr14 73023364 N chr14 73023473 N DUP 10
SRR1766484.7356431 chr14 73023333 N chr14 73023471 N DUP 12
SRR1766451.1833916 chr14 73023333 N chr14 73023471 N DUP 13
SRR1766475.449926 chr14 73023333 N chr14 73023471 N DUP 13
SRR1766442.34510338 chr14 73023333 N chr14 73023471 N DUP 15
SRR1766448.9732904 chr14 73023333 N chr14 73023471 N DUP 17
SRR1766484.7564148 chr14 73023400 N chr14 73023455 N DEL 17
SRR1766444.2549652 chr14 73023401 N chr14 73023454 N DUP 13
SRR1766469.5986209 chr14 73023401 N chr14 73023454 N DUP 13
SRR1766483.1305459 chr14 73023401 N chr14 73023454 N DUP 13
SRR1766464.9278956 chr14 73023401 N chr14 73023454 N DUP 15
SRR1766463.7845313 chr14 73023401 N chr14 73023454 N DUP 15
SRR1766446.7593408 chr14 73023401 N chr14 73023454 N DUP 15
SRR1766443.9294079 chr14 73023401 N chr14 73023454 N DUP 15
SRR1766446.1327521 chr14 73023400 N chr14 73023455 N DEL 15
SRR1766446.7965769 chr14 73023400 N chr14 73023455 N DEL 15
SRR1766442.22081457 chr14 73023400 N chr14 73023455 N DEL 15
SRR1766458.1247687 chr14 73023400 N chr14 73023455 N DEL 15
SRR1766447.6500876 chr14 73023400 N chr14 73023455 N DEL 14
SRR1766452.3441462 chr14 73023400 N chr14 73023455 N DEL 13
SRR1766457.4836368 chr12 124416701 N chr12 124416880 N DEL 16
SRR1766476.4800941 chr12 124416743 N chr12 124416957 N DEL 10
SRR1766452.4302792 chr5 142075446 N chr5 142075623 N DUP 14
SRR1766484.4528833 chr5 142075637 N chr5 142075937 N DEL 10
SRR1766480.7340283 chr5 142075637 N chr5 142075937 N DEL 10
SRR1766472.6419271 chr5 142075446 N chr5 142075623 N DUP 10
SRR1766468.2833133 chr5 142075664 N chr5 142075965 N DEL 11
SRR1766442.13700379 chr5 142075662 N chr5 142075962 N DEL 11
SRR1766467.10704287 chr5 142075767 N chr5 142076495 N DUP 13
SRR1766461.3811885 chr5 142075724 N chr5 142075823 N DUP 12
SRR1766442.23039326 chr5 142075621 N chr5 142075724 N DEL 12
SRR1766473.9003948 chr5 142075621 N chr5 142075724 N DEL 12
SRR1766448.1539612 chr5 142075629 N chr5 142075731 N DEL 11
SRR1766461.3811885 chr5 142075724 N chr5 142075823 N DUP 18
SRR1766473.6757673 chr5 142075722 N chr5 142075774 N DEL 13
SRR1766464.4547729 chr5 142075440 N chr5 142075725 N DEL 16
SRR1766458.4332305 chr5 142075715 N chr5 142075767 N DEL 18
SRR1766478.4332944 chr5 142075421 N chr5 142075757 N DEL 11
SRR1766451.9203540 chr5 142075437 N chr5 142075865 N DUP 12
SRR1766448.8697066 chr5 142075434 N chr5 142075867 N DEL 16
SRR1766473.10887337 chr5 142075434 N chr5 142075867 N DEL 16
SRR1766469.3578124 chr5 142075434 N chr5 142075867 N DEL 16
SRR1766476.1049434 chr5 142075435 N chr5 142075868 N DEL 14
SRR1766469.3578124 chr5 142075507 N chr5 142075983 N DUP 10
SRR1766482.2601077 chr5 142075610 N chr5 142076011 N DEL 16
SRR1766471.2889692 chr5 142075610 N chr5 142076011 N DEL 16
SRR1766485.9762040 chr5 142075756 N chr5 142076128 N DUP 10
SRR1766462.2882869 chr5 142076099 N chr5 142076377 N DEL 10
SRR1766446.212741 chr5 142076099 N chr5 142076327 N DEL 14
SRR1766483.4753866 chr5 142076099 N chr5 142076327 N DEL 13
SRR1766465.2076561 chr5 142075605 N chr5 142075956 N DEL 10
SRR1766460.1780949 chr5 142075603 N chr5 142075757 N DEL 10
SRR1766452.3788665 chr5 142075802 N chr5 142076580 N DEL 11
SRR1766450.5226772 chr2 240357809 N chr2 240357930 N DEL 17
SRR1766486.10854292 chr12 122731874 N chr12 122732098 N DUP 14
SRR1766459.11200037 chr19 28114323 N chr19 28114386 N DUP 17
SRR1766445.3464747 chr19 28114323 N chr19 28114386 N DUP 16
SRR1766465.4292348 chr8 116297695 N chr8 116297929 N DEL 12
SRR1766472.9166088 chr6 166955879 N chr6 166956030 N DEL 11
SRR1766470.347213 chr14 86443422 N chr14 86443494 N DEL 14
SRR1766477.11133941 chr14 86443635 N chr14 86443737 N DEL 17
SRR1766457.8113491 chr14 86443635 N chr14 86443737 N DEL 17
SRR1766442.42952005 chr14 86443635 N chr14 86443737 N DEL 17
SRR1766478.5238000 chr14 86443435 N chr14 86443685 N DEL 18
SRR1766483.407243 chr14 86443438 N chr14 86443688 N DEL 12
SRR1766450.8836247 chr14 86443661 N chr14 86443737 N DEL 16
SRR1766442.22992507 chr14 86443691 N chr14 86443767 N DEL 16
SRR1766479.4639488 chr14 86443661 N chr14 86443737 N DEL 11
SRR1766459.3077224 chr14 86443661 N chr14 86443737 N DEL 11
SRR1766474.8929750 chr14 86443661 N chr14 86443737 N DEL 11
SRR1766473.8607299 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766452.7161305 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766482.5713540 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766469.2243889 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766484.2829057 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766442.24853383 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766451.2672792 chr14 86444057 N chr14 86444117 N DEL 15
SRR1766442.22992507 chr14 86444057 N chr14 86444117 N DEL 16
SRR1766463.349530 chr14 86443590 N chr14 86444058 N DUP 16
SRR1766454.2140418 chr14 86444059 N chr14 86444112 N DEL 16
SRR1766483.3498350 chr14 86444059 N chr14 86444112 N DEL 16
SRR1766473.9157197 chr14 86443397 N chr14 86444095 N DUP 10
SRR1766461.6828702 chr14 86443959 N chr14 86444072 N DEL 19
SRR1766464.8581884 chr14 86443425 N chr14 86444072 N DEL 11
SRR1766479.10343351 chr14 86443425 N chr14 86444072 N DEL 10
SRR1766460.3863870 chr14 86443523 N chr14 86444112 N DEL 17
SRR1766442.6134313 chr14 86443525 N chr14 86444114 N DEL 13
SRR1766445.8947762 chr12 127166345 N chr12 127166404 N DUP 16
SRR1766477.9796204 chr12 127166345 N chr12 127166404 N DUP 17
SRR1766467.4660244 chr12 127166345 N chr12 127166404 N DUP 19
SRR1766473.4510760 chr12 127166395 N chr12 127166484 N DUP 10
SRR1766446.4228944 chr12 127166395 N chr12 127166484 N DUP 10
SRR1766480.6313399 chr18 48221288 N chr18 48221536 N DEL 15
SRR1766482.11101854 chr5 174522637 N chr5 174522704 N DEL 12
SRR1766443.2661640 chr5 174522603 N chr5 174522705 N DEL 10
SRR1766485.5863310 chr5 174522603 N chr5 174522707 N DEL 12
SRR1766475.4721310 chr2 16143671 N chr2 16145308 N DUP 10
SRR1766442.25173893 chr2 16143762 N chr2 16145266 N DEL 13
SRR1766478.6518221 chr2 16144013 N chr2 16145309 N DUP 13
SRR1766442.19880547 chr17 42123845 N chr17 42124168 N DUP 13
SRR1766443.7451191 chr3 93470409 N chr3 93470458 N DUP 17
SRR1766463.4981021 chr3 93470409 N chr3 93470458 N DUP 16
SRR1766475.5824442 chr3 93470409 N chr3 93470458 N DUP 18
SRR1766480.3157736 chr19 49612047 N chr19 49612354 N DEL 10
SRR1766442.16666031 chr10 7378306 N chr10 7378355 N DUP 15
SRR1766442.22774063 chr10 7378306 N chr10 7378355 N DUP 12
SRR1766452.1763621 chr10 7378306 N chr10 7378355 N DUP 12
SRR1766475.1516451 chr15 66381223 N chr15 66381852 N DEL 10
SRR1766442.32608465 chr2 239421632 N chr2 239421816 N DEL 10
SRR1766442.31053216 chr2 239421632 N chr2 239421816 N DEL 14
SRR1766444.1848128 chr2 239421591 N chr2 239421775 N DEL 13
SRR1766460.3406860 chr3 35748213 N chr3 35748434 N DEL 13
SRR1766462.5665021 chr3 35748113 N chr3 35748280 N DEL 10
SRR1766442.6201418 chr3 35748432 N chr3 35748636 N DUP 10
SRR1766486.1735191 chr12 34301311 N chr12 34301733 N DEL 15
SRR1766445.8880094 chr12 34301305 N chr12 34301727 N DEL 10
SRR1766485.9240589 chr12 34301349 N chr12 34302190 N DEL 12
SRR1766478.6052757 chr12 34301422 N chr12 34302475 N DEL 15
SRR1766477.895066 chr2 33911356 N chr2 33911419 N DEL 12
SRR1766480.8159475 chr1 220012938 N chr1 220013042 N DUP 16
SRR1766478.4506607 chr1 220012938 N chr1 220013042 N DUP 13
SRR1766457.8397286 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766450.7496326 chr1 220012938 N chr1 220013042 N DUP 14
SRR1766484.5501658 chr1 220012938 N chr1 220013042 N DUP 14
SRR1766461.2699270 chr1 220012938 N chr1 220013042 N DUP 11
SRR1766472.11486622 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766447.7842760 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766474.8348644 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766442.29118002 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766482.4618864 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766442.37559474 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766447.1280491 chr1 220012938 N chr1 220013042 N DUP 11
SRR1766466.5201590 chr1 220012938 N chr1 220013042 N DUP 11
SRR1766485.7704134 chr1 11135798 N chr1 11136100 N DEL 14
SRR1766469.8596490 chr7 138174569 N chr7 138174662 N DEL 13
SRR1766474.9648697 chr7 138174569 N chr7 138174662 N DEL 13
SRR1766442.23752160 chr7 138174569 N chr7 138174662 N DEL 13
SRR1766472.8479695 chr6 23802191 N chr6 23802302 N DEL 12
SRR1766484.7172295 chr6 23802192 N chr6 23802303 N DEL 11
SRR1766445.1875357 chr12 116652096 N chr12 116652199 N DUP 13
SRR1766480.3500644 chr12 116652096 N chr12 116652199 N DUP 13
SRR1766476.2952469 chr12 116652002 N chr12 116652198 N DUP 12
SRR1766469.8966842 chr12 116652032 N chr12 116652178 N DEL 12
SRR1766470.878799 chr12 116652025 N chr12 116652175 N DEL 15
SRR1766462.7735033 chr12 116652114 N chr12 116652175 N DEL 17
SRR1766465.326487 chr12 116652110 N chr12 116652175 N DEL 15
SRR1766478.2955197 chr12 116652110 N chr12 116652179 N DEL 11
SRR1766478.767736 chr4 163894706 N chr4 163894774 N DUP 18
SRR1766483.4538915 chr4 163894780 N chr4 163894840 N DEL 18
SRR1766486.11865358 chr4 163894780 N chr4 163894840 N DEL 18
SRR1766466.5281676 chr4 163894706 N chr4 163894774 N DUP 19
SRR1766479.8449256 chr4 163894706 N chr4 163894774 N DUP 19
SRR1766444.2914134 chr4 163894706 N chr4 163894774 N DUP 19
SRR1766448.2239811 chr4 163894821 N chr4 163894904 N DUP 11
SRR1766451.6251880 chr4 163894734 N chr4 163894840 N DEL 12
SRR1766463.8626599 chr4 163894713 N chr4 163894779 N DUP 16
SRR1766453.6990199 chrX 57698243 N chrX 57698806 N DUP 15
SRR1766479.1250646 chrX 57698279 N chrX 57698704 N DEL 15
SRR1766447.11392507 chrX 57698303 N chrX 57698402 N DUP 17
SRR1766472.11492922 chrX 57698191 N chrX 57698743 N DUP 19
SRR1766480.8317691 chrX 57697517 N chrX 57698793 N DUP 16
SRR1766447.8639660 chrX 57698637 N chrX 57698711 N DUP 19
SRR1766455.3622714 chrX 57698385 N chrX 57698792 N DEL 11
SRR1766464.6462547 chrX 57698325 N chrX 57698800 N DEL 15
SRR1766443.9148985 chr12 163361 N chr12 163520 N DUP 10
SRR1766463.1360890 chr8 675298 N chr8 676149 N DEL 10
SRR1766448.3331198 chr8 675381 N chr8 675545 N DUP 10
SRR1766460.1098885 chr8 675381 N chr8 675545 N DUP 10
SRR1766472.9457855 chr8 676177 N chr8 676312 N DUP 10
SRR1766471.265141 chr8 676153 N chr8 676209 N DEL 10
SRR1766448.5518291 chr8 675994 N chr8 676377 N DUP 17
SRR1766479.6653007 chr8 675814 N chr8 676388 N DUP 10
SRR1766448.10430876 chr8 675511 N chr8 676388 N DUP 13
SRR1766460.8211552 chr8 675511 N chr8 676388 N DUP 10
SRR1766477.3212384 chr8 675994 N chr8 676377 N DUP 17
SRR1766454.2962923 chr8 675511 N chr8 676388 N DUP 12
SRR1766447.6296919 chr8 675867 N chr8 676637 N DEL 16
SRR1766454.4311037 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766442.23620487 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766444.1123921 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766461.3364703 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766474.11180459 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766474.4132836 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766477.5017017 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766477.7916256 chr1 118319485 N chr1 118319548 N DUP 14
SRR1766442.40045430 chr2 131754522 N chr2 131754918 N DEL 10
SRR1766474.640842 chr2 131754646 N chr2 131755480 N DEL 15
SRR1766448.8849974 chr2 131755218 N chr2 131755438 N DEL 10
SRR1766471.5055056 chr2 131754091 N chr2 131755332 N DEL 14
SRR1766462.8268510 chr2 131754562 N chr2 131755396 N DEL 10
SRR1766451.1949286 chr2 131754236 N chr2 131755480 N DUP 10
SRR1766478.8628814 chr2 131754236 N chr2 131755679 N DUP 10
SRR1766442.438630 chrY 10924454 N chrY 10924538 N DUP 15
SRR1766474.11222621 chr7 121088825 N chr7 121088942 N DUP 10
SRR1766442.35404240 chr4 3809314 N chr4 3809470 N DEL 12
SRR1766466.8611578 chr3 84516559 N chr3 84516737 N DUP 12
SRR1766467.2451381 chr3 84516559 N chr3 84516737 N DUP 12
SRR1766484.399139 chr3 84516559 N chr3 84516737 N DUP 12
SRR1766443.8950394 chr3 84516559 N chr3 84516737 N DUP 12
SRR1766478.7061796 chr3 84516729 N chr3 84516792 N DUP 16
SRR1766479.10019109 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766473.706836 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766485.912074 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766452.5053281 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766465.2700061 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766471.10810924 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766453.4648880 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766480.6438425 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766485.2059701 chr17 77920548 N chr17 77920681 N DUP 15
SRR1766446.5387252 chr10 445895 N chr10 446152 N DEL 10
SRR1766472.4128835 chr22 10629003 N chr22 10629082 N DEL 15
SRR1766452.2375989 chr22 10629003 N chr22 10629082 N DEL 15
SRR1766455.8706832 chr17 8052954 N chr17 8053049 N DEL 11
SRR1766485.6518993 chr17 8052954 N chr17 8053049 N DEL 12
SRR1766484.9768915 chr17 8052954 N chr17 8053049 N DEL 13
SRR1766465.1484519 chr17 8052954 N chr17 8053049 N DEL 13
SRR1766454.10234852 chr17 8052954 N chr17 8053049 N DEL 13
SRR1766456.1296154 chr17 8052954 N chr17 8053049 N DEL 13
SRR1766452.10404207 chr17 8053023 N chr17 8053112 N DEL 13
SRR1766484.3957709 chr17 8053007 N chr17 8053114 N DEL 13
SRR1766486.4365436 chr17 8053010 N chr17 8053117 N DEL 10
SRR1766448.8630962 chr17 8052848 N chr17 8053257 N DEL 15
SRR1766451.6944760 chr8 35305719 N chr8 35305931 N DEL 13
SRR1766449.9118938 chr19 3988963 N chr19 3989266 N DEL 10
SRR1766450.4700379 chr19 3988752 N chr19 3989056 N DEL 18
SRR1766481.8708133 chr19 3989084 N chr19 3989384 N DEL 10
SRR1766449.10330924 chr3 159680789 N chr3 159680851 N DUP 11
SRR1766442.21337461 chr3 159680771 N chr3 159680878 N DEL 12
SRR1766482.3744270 chr3 159680752 N chr3 159680887 N DUP 10
SRR1766484.3109046 chr3 159680738 N chr3 159680865 N DEL 14
SRR1766465.8793087 chrX 72179191 N chrX 72179359 N DEL 15
SRR1766474.3696003 chrX 72179191 N chrX 72179359 N DEL 15
SRR1766477.11008970 chr10 25241326 N chr10 25241398 N DUP 13
SRR1766467.7692096 chr10 25241351 N chr10 25241429 N DEL 13
SRR1766460.3490834 chr10 25241352 N chr10 25241430 N DEL 12
SRR1766476.9861398 chr10 25241351 N chr10 25241429 N DEL 14
SRR1766476.1574992 chr11 68861420 N chr11 68861577 N DEL 10
SRR1766448.3072456 chrX 40236844 N chrX 40237012 N DEL 11
SRR1766445.9416049 chr3 143449252 N chr3 143449760 N DEL 19
SRR1766464.5327466 chr3 143449252 N chr3 143449760 N DEL 19
SRR1766447.6856747 chr3 143449252 N chr3 143449760 N DEL 16
SRR1766455.391530 chr3 143449252 N chr3 143449760 N DEL 16
SRR1766461.9614609 chr3 143449198 N chr3 143449763 N DEL 18
SRR1766460.2179095 chr3 143449252 N chr3 143449760 N DEL 19
SRR1766473.7367585 chr3 143449196 N chr3 143449760 N DEL 17
SRR1766469.10897100 chr3 143449198 N chr3 143449763 N DEL 18
SRR1766461.682331 chr3 143449198 N chr3 143449763 N DEL 18
SRR1766475.8273833 chr3 143449133 N chr3 143449810 N DUP 14
SRR1766473.5147936 chr3 143449234 N chr3 143449799 N DEL 15
SRR1766462.3324729 chr3 143449198 N chr3 143449763 N DEL 19
SRR1766462.1510450 chr3 143449763 N chr3 143449874 N DUP 12
SRR1766464.6039803 chr3 143449133 N chr3 143449810 N DUP 14
SRR1766475.10552202 chr3 143449763 N chr3 143449874 N DUP 12
SRR1766473.5033895 chr3 143449493 N chr3 143449632 N DUP 19
SRR1766475.6857724 chr3 143449750 N chr3 143449847 N DEL 19
SRR1766470.2228423 chr3 143449056 N chr3 143449826 N DEL 10
SRR1766447.3401251 chr3 143450052 N chr3 143450294 N DEL 10
SRR1766465.10431200 chr3 143450052 N chr3 143450294 N DEL 11
SRR1766481.10440938 chr11 104791539 N chr11 104791655 N DUP 12
SRR1766442.42910138 chr2 241628894 N chr2 241629075 N DEL 10
SRR1766452.10635577 chr18 54780361 N chr18 54780619 N DEL 10
SRR1766475.2950261 chr12 39713044 N chr12 39713141 N DEL 12
SRR1766477.5568562 chr12 39713045 N chr12 39713142 N DEL 11
SRR1766474.3725297 chr12 39712968 N chr12 39713175 N DEL 14
SRR1766464.4222708 chr17 47666647 N chr17 47666705 N DEL 10
SRR1766442.18831192 chr11 47657874 N chr11 47658177 N DUP 12
SRR1766463.8817437 chr7 100995441 N chr7 100996112 N DEL 12
SRR1766442.2648770 chr7 100995188 N chr7 100995936 N DEL 15
SRR1766467.8370489 chr10 126947606 N chr10 126948140 N DUP 16
SRR1766462.3225095 chr10 126947499 N chr10 126947633 N DEL 10
SRR1766455.9689092 chr10 126947496 N chr10 126948194 N DUP 11
SRR1766470.1317365 chr10 126947489 N chr10 126948090 N DEL 10
SRR1766444.6514218 chr10 126947529 N chr10 126947598 N DEL 13
SRR1766452.10600804 chr10 126947693 N chr10 126947895 N DEL 11
SRR1766456.5088505 chr10 126947625 N chr10 126948056 N DEL 10
SRR1766458.1373923 chr10 126947464 N chr10 126948096 N DEL 10
SRR1766473.4331467 chr10 126947439 N chr10 126948341 N DUP 13
SRR1766449.2965602 chr10 126947761 N chr10 126948130 N DEL 11
SRR1766452.10414938 chr10 126947663 N chr10 126947996 N DUP 10
SRR1766481.10877174 chr10 126947668 N chr10 126948569 N DEL 16
SRR1766472.11832695 chr10 126947950 N chr10 126948087 N DEL 15
SRR1766482.1453658 chr10 126947653 N chr10 126948087 N DEL 10
SRR1766455.5821830 chr10 126947524 N chr10 126947953 N DUP 13
SRR1766457.2896017 chr10 126948070 N chr10 126948140 N DUP 16
SRR1766442.21048004 chr10 126947576 N chr10 126948072 N DEL 16
SRR1766442.31900206 chr10 126948056 N chr10 126948358 N DUP 10
SRR1766473.252871 chr10 126947524 N chr10 126948355 N DUP 10
SRR1766468.1270051 chr10 126947979 N chr10 126948244 N DUP 13
SRR1766484.3945647 chr10 126947791 N chr10 126948189 N DUP 10
SRR1766455.7700498 chr10 126947462 N chr10 126948060 N DEL 10
SRR1766442.43338461 chr10 126947854 N chr10 126948056 N DEL 10
SRR1766471.5691776 chr10 126947597 N chr10 126947861 N DEL 10
SRR1766442.24107140 chr10 126947589 N chr10 126947984 N DUP 11
SRR1766465.2860578 chr10 126947524 N chr10 126947919 N DUP 13
SRR1766473.6500454 chr10 126947496 N chr10 126948160 N DUP 11
SRR1766469.9360861 chr10 126947640 N chr10 126948174 N DUP 19
SRR1766478.9289682 chr10 126948065 N chr10 126948129 N DUP 10
SRR1766484.3775872 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766463.5343559 chr10 126947422 N chr10 126947591 N DUP 11
SRR1766464.8723702 chr10 126947456 N chr10 126948191 N DUP 19
SRR1766462.816657 chr10 126947792 N chr10 126948162 N DUP 10
SRR1766458.6555825 chr10 126947554 N chr10 126947855 N DEL 13
SRR1766473.9671552 chr10 126947467 N chr10 126947762 N DEL 16
SRR1766458.5078900 chr10 126947983 N chr10 126948568 N DEL 10
SRR1766446.4487313 chr10 126947497 N chr10 126947796 N DUP 11
SRR1766443.10323761 chr10 126947458 N chr10 126948155 N DEL 11
SRR1766442.18391058 chr10 126947600 N chr10 126948569 N DEL 16
SRR1766470.1057442 chr10 126947538 N chr10 126947602 N DUP 10
SRR1766456.2981003 chr10 126947492 N chr10 126947589 N DEL 14
SRR1766451.8791147 chr10 126948056 N chr10 126948358 N DUP 10
SRR1766456.3242720 chr10 126947472 N chr10 126948073 N DEL 15
SRR1766443.9825540 chr10 126947586 N chr10 126947981 N DUP 13
SRR1766468.5746192 chr10 126947492 N chr10 126948087 N DEL 14
SRR1766481.12493910 chr10 126947422 N chr10 126947758 N DUP 11
SRR1766463.4334193 chr10 126947612 N chr10 126948074 N DEL 15
SRR1766464.10586500 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766464.10354857 chr10 126947560 N chr10 126948062 N DEL 10
SRR1766465.6816635 chr10 126947529 N chr10 126947700 N DEL 13
SRR1766476.7715033 chr10 126947490 N chr10 126948058 N DUP 10
SRR1766479.6760768 chr10 126947555 N chr10 126948259 N DUP 16
SRR1766452.1086251 chr10 126947829 N chr10 126947998 N DUP 10
SRR1766476.9192109 chr10 126947690 N chr10 126948056 N DEL 10
SRR1766447.10618584 chr10 126947567 N chr10 126948197 N DUP 13
SRR1766476.6964575 chr10 126947490 N chr10 126947690 N DUP 10
SRR1766483.8768564 chr10 126947490 N chr10 126947724 N DUP 10
SRR1766463.10781725 chr10 126947458 N chr10 126947688 N DEL 11
SRR1766464.9185707 chr10 126947461 N chr10 126947530 N DEL 10
SRR1766486.3159852 chr10 126947496 N chr10 126947665 N DUP 10
SRR1766476.5666329 chr10 126947524 N chr10 126947953 N DUP 13
SRR1766477.7448786 chr10 126947464 N chr10 126948099 N DEL 10
SRR1766483.8061414 chr10 126947687 N chr10 126947957 N DEL 11
SRR1766476.8762156 chr10 126947453 N chr10 126947553 N DEL 10
SRR1766480.4180718 chr10 126947928 N chr10 126948065 N DEL 10
SRR1766467.3799356 chr10 126947854 N chr10 126948056 N DEL 10
SRR1766455.9053641 chr10 126947600 N chr10 126948569 N DEL 16
SRR1766486.7105853 chr10 126948154 N chr10 126948294 N DEL 11
SRR1766463.7227385 chr10 126947885 N chr10 126948090 N DEL 13
SRR1766484.5083173 chr10 126947854 N chr10 126948056 N DEL 10
SRR1766477.10130098 chr10 126947473 N chr10 126947673 N DUP 14
SRR1766458.6555825 chr10 126947554 N chr10 126948192 N DEL 13
SRR1766476.7878364 chr10 126947458 N chr10 126948087 N DEL 11
SRR1766473.5082680 chr10 126947619 N chr10 126948087 N DEL 10
SRR1766474.6464341 chr10 126947467 N chr10 126947762 N DEL 11
SRR1766445.8873658 chr10 126947487 N chr10 126947687 N DUP 10
SRR1766447.3414984 chr10 126947537 N chr10 126948070 N DEL 10
SRR1766465.7527784 chr10 126947464 N chr10 126948065 N DEL 10
SRR1766479.2610269 chr10 126947601 N chr10 126947696 N DUP 13
SRR1766442.26515337 chr10 126947690 N chr10 126948056 N DEL 10
SRR1766466.5228074 chr10 126947557 N chr10 126948022 N DEL 13
SRR1766447.9463604 chr10 126948030 N chr10 126948130 N DEL 10
SRR1766481.4694938 chr10 126947588 N chr10 126948294 N DEL 13
SRR1766476.3797964 chr10 126947526 N chr10 126947632 N DEL 13
SRR1766474.8064010 chr10 126947762 N chr10 126947897 N DUP 11
SRR1766478.6182520 chr10 126947632 N chr10 126947693 N DUP 15
SRR1766463.10450632 chr10 126947589 N chr10 126947659 N DUP 16
SRR1766463.172660 chr10 126947589 N chr10 126948321 N DUP 10
SRR1766453.9252034 chr10 126947623 N chr10 126947890 N DEL 10
SRR1766472.11290418 chr10 126947499 N chr10 126948197 N DUP 13
SRR1766482.1000987 chr10 126947625 N chr10 126948155 N DEL 11
SRR1766457.2011452 chr10 126948087 N chr10 126948185 N DUP 15
SRR1766473.1787874 chr10 126947574 N chr10 126948176 N DUP 12
SRR1766454.5842197 chr10 126947608 N chr10 126948070 N DEL 16
SRR1766479.12517576 chr10 126947537 N chr10 126948070 N DEL 10
SRR1766442.743146 chr10 126947479 N chr10 126948080 N DEL 15
SRR1766459.7799527 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766447.4034789 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766466.8330554 chr10 126947928 N chr10 126948065 N DEL 10
SRR1766460.1682100 chr10 126947416 N chr10 126948049 N DUP 10
SRR1766465.3944793 chr10 126947461 N chr10 126948056 N DEL 13
SRR1766469.7597183 chr10 126947998 N chr10 126948132 N DEL 10
SRR1766468.3568200 chr10 126947625 N chr10 126948056 N DEL 10
SRR1766473.4539366 chr10 126947424 N chr10 126948056 N DEL 10
SRR1766471.6935264 chr10 126947684 N chr10 126947988 N DEL 13
SRR1766442.35813991 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766445.6817241 chr10 126947475 N chr10 126947774 N DUP 13
SRR1766452.5933781 chr10 126947692 N chr10 126948129 N DEL 12
SRR1766470.6100919 chr10 126948073 N chr10 126948174 N DUP 10
SRR1766483.800063 chr10 126947521 N chr10 126947659 N DUP 16
SRR1766449.8384614 chr10 126948090 N chr10 126948188 N DUP 10
SRR1766463.10450632 chr10 126947467 N chr10 126948062 N DEL 13
SRR1766446.54148 chr10 126947600 N chr10 126948569 N DEL 16
SRR1766473.332021 chr10 126947965 N chr10 126948569 N DEL 16
SRR1766442.33223973 chr10 126947483 N chr10 126948118 N DEL 10
SRR1766469.7094554 chr10 126947557 N chr10 126948121 N DEL 16
SRR1766473.9135770 chr10 126947560 N chr10 126947756 N DEL 19
SRR1766443.4926066 chr10 126947600 N chr10 126948569 N DEL 16
SRR1766442.7834194 chr4 146008342 N chr4 146008432 N DEL 10
SRR1766455.6878962 chr9 95083489 N chr9 95083585 N DUP 10
SRR1766459.4254733 chr22 12571521 N chr22 12571575 N DEL 16
SRR1766451.2501926 chr14 65692608 N chr14 65692659 N DEL 11
SRR1766473.5567176 chr14 65692608 N chr14 65692659 N DEL 11
SRR1766451.9326935 chr14 65692608 N chr14 65692659 N DEL 11
SRR1766450.9586330 chr14 65692608 N chr14 65692659 N DEL 11
SRR1766486.1974416 chr14 65692559 N chr14 65692659 N DEL 11
SRR1766477.11545340 chr14 65692560 N chr14 65692660 N DEL 11
SRR1766460.1278588 chr14 65692558 N chr14 65692658 N DEL 11
SRR1766486.11290209 chr10 52834578 N chr10 52834717 N DEL 12
SRR1766446.10614688 chr10 52834357 N chr10 52835506 N DUP 16
SRR1766482.3501267 chr10 52834343 N chr10 52834494 N DUP 16
SRR1766449.8174668 chr10 52835303 N chr10 52835477 N DEL 10
SRR1766457.8165387 chr10 52834976 N chr10 52835039 N DUP 18
SRR1766475.6106743 chr10 52835035 N chr10 52835450 N DEL 16
SRR1766449.968100 chr10 52834920 N chr10 52835443 N DEL 18
SRR1766475.897889 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766469.4864618 chr10 52834137 N chr10 52834343 N DEL 12
SRR1766443.10336536 chr10 52834262 N chr10 52834925 N DUP 17
SRR1766459.3416325 chr10 52834566 N chr10 52834751 N DEL 11
SRR1766445.998017 chr10 52834902 N chr10 52834959 N DEL 12
SRR1766461.8929824 chr10 52834328 N chr10 52834861 N DUP 10
SRR1766481.9970168 chr10 52835344 N chr10 52835516 N DUP 10
SRR1766450.5499935 chr10 52834845 N chr10 52834903 N DEL 10
SRR1766442.1991002 chr10 52835233 N chr10 52835477 N DEL 14
SRR1766481.7605879 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766470.4965910 chr10 52834920 N chr10 52835443 N DEL 11
SRR1766469.7981130 chr10 52834159 N chr10 52834344 N DEL 10
SRR1766477.6236954 chr10 52834513 N chr10 52834668 N DUP 16
SRR1766483.8037494 chr10 52834271 N chr10 52834472 N DUP 18
SRR1766447.5677813 chr10 52834663 N chr10 52834932 N DUP 17
SRR1766443.1483430 chr10 52834262 N chr10 52834925 N DUP 14
SRR1766451.4111021 chr10 52834352 N chr10 52834901 N DUP 11
SRR1766482.2991508 chr10 52834307 N chr10 52834538 N DEL 11
SRR1766459.10529944 chr10 52834299 N chr10 52834675 N DEL 13
SRR1766484.1379780 chr10 52834190 N chr10 52834464 N DUP 12
SRR1766476.9776208 chr10 52834578 N chr10 52834717 N DEL 13
SRR1766486.8024372 chr10 52834357 N chr10 52834419 N DUP 16
SRR1766486.5568017 chr10 52834468 N chr10 52835479 N DEL 14
SRR1766482.7760437 chr10 52834451 N chr10 52835482 N DEL 11
SRR1766473.7015063 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766455.8223662 chr10 52834663 N chr10 52834932 N DUP 17
SRR1766461.4776924 chr10 52834904 N chr10 52834961 N DEL 12
SRR1766444.6733059 chr10 52835062 N chr10 52835477 N DEL 11
SRR1766448.6669711 chr10 52834180 N chr10 52834262 N DUP 19
SRR1766476.3496000 chr10 52834228 N chr10 52834360 N DEL 12
SRR1766475.3720762 chr10 52834217 N chr10 52834899 N DEL 12
SRR1766460.37586 chr10 52834606 N chr10 52834886 N DUP 19
SRR1766462.8407781 chr10 52835233 N chr10 52835477 N DEL 14
SRR1766452.5180251 chr10 52834527 N chr10 52834878 N DUP 11
SRR1766442.41431891 chr10 52834333 N chr10 52834392 N DUP 15
SRR1766459.4892629 chr10 52834527 N chr10 52834878 N DUP 11
SRR1766454.3397677 chr10 52834348 N chr10 52834444 N DUP 10
SRR1766457.451781 chr10 52834513 N chr10 52834668 N DUP 15
SRR1766485.2831073 chr10 52834180 N chr10 52834262 N DUP 19
SRR1766450.9493129 chr10 52834213 N chr10 52834296 N DUP 15
SRR1766472.7631750 chr10 52834219 N chr10 52834352 N DEL 11
SRR1766475.5829802 chr10 52834282 N chr10 52834479 N DEL 18
SRR1766479.744178 chr10 52834299 N chr10 52834675 N DEL 14
SRR1766442.14019273 chr10 52834527 N chr10 52834878 N DUP 11
SRR1766454.4786326 chr10 52834468 N chr10 52835479 N DEL 15
SRR1766478.2839191 chr10 52834529 N chr10 52834587 N DEL 14
SRR1766442.42273243 chr10 52834343 N chr10 52834400 N DUP 11
SRR1766479.5222674 chr10 52834248 N chr10 52834457 N DUP 18
SRR1766448.2894725 chr10 52834573 N chr10 52834758 N DEL 11
SRR1766446.10614688 chr10 52834180 N chr10 52834262 N DUP 16
SRR1766449.5184961 chr10 52834462 N chr10 52834649 N DEL 17
SRR1766477.8918353 chr10 52835062 N chr10 52835477 N DEL 14
SRR1766471.5208502 chr10 52834309 N chr10 52834385 N DUP 14
SRR1766481.10193444 chr10 52835128 N chr10 52835477 N DEL 14
SRR1766453.3279804 chr10 52834663 N chr10 52834932 N DUP 12
SRR1766475.9590094 chr10 52834171 N chr10 52834445 N DUP 16
SRR1766448.1365620 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766482.5479155 chr10 52834959 N chr10 52835506 N DUP 17
SRR1766468.4270493 chr10 52834196 N chr10 52834313 N DUP 16
SRR1766449.3394212 chr10 52834329 N chr10 52834501 N DEL 10
SRR1766454.8238494 chr10 52834214 N chr10 52834333 N DEL 14
SRR1766458.2707345 chr10 52834309 N chr10 52834433 N DUP 10
SRR1766483.3848811 chr10 52834959 N chr10 52835506 N DUP 15
SRR1766448.5502724 chr10 52834468 N chr10 52835479 N DEL 14
SRR1766483.4662958 chr10 52834235 N chr10 52834755 N DEL 13
SRR1766448.6012014 chr10 52835316 N chr10 52835500 N DEL 14
SRR1766457.6722196 chr10 52834215 N chr10 52834348 N DEL 15
SRR1766467.961717 chr10 52834208 N chr10 52834341 N DEL 17
SRR1766473.3750949 chr10 52834246 N chr10 52834302 N DUP 15
SRR1766470.2999087 chr10 52834262 N chr10 52834423 N DUP 13
SRR1766448.10886233 chr10 52835128 N chr10 52835477 N DEL 14
SRR1766462.8407781 chr10 52834272 N chr10 52835317 N DUP 12
SRR1766459.4380243 chr10 52834526 N chr10 52834663 N DUP 17
SRR1766464.6430532 chr10 52834343 N chr10 52834494 N DUP 12
SRR1766442.14654078 chr10 52834343 N chr10 52834494 N DUP 15
SRR1766459.11359956 chr10 52834348 N chr10 52834444 N DUP 15
SRR1766459.141569 chr10 52834985 N chr10 52835480 N DEL 11
SRR1766442.27176991 chr10 52834399 N chr10 52834662 N DEL 19
SRR1766442.18310656 chr10 52834374 N chr10 52834538 N DEL 16
SRR1766461.2952880 chr10 52834592 N chr10 52834669 N DUP 14
SRR1766458.5578702 chr10 52834215 N chr10 52834348 N DEL 15
SRR1766469.4913358 chr10 52834302 N chr10 52834512 N DEL 15
SRR1766482.3501267 chr10 52834364 N chr10 52834435 N DEL 16
SRR1766469.4130133 chr10 52834606 N chr10 52834886 N DUP 18
SRR1766476.5757096 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766465.8571054 chr10 52834287 N chr10 52834636 N DUP 16
SRR1766442.6349846 chr10 52834211 N chr10 52834528 N DUP 11
SRR1766459.4207964 chr10 52834222 N chr10 52834896 N DEL 15
SRR1766464.46233 chr10 52834566 N chr10 52834751 N DEL 11
SRR1766448.5519213 chr10 52834307 N chr10 52834538 N DEL 10
SRR1766454.1715984 chr7 152487421 N chr7 152487490 N DEL 11
SRR1766455.7967884 chr18 1747201 N chr18 1747262 N DUP 15
SRR1766482.5069586 chr18 1747189 N chr18 1747282 N DUP 19
SRR1766470.774084 chr18 1747179 N chr18 1747252 N DUP 18
SRR1766464.8511475 chr18 1747181 N chr18 1747280 N DUP 17
SRR1766485.11357864 chr18 1747179 N chr18 1747270 N DUP 14
SRR1766464.8756450 chr18 1747223 N chr18 1747310 N DUP 12
SRR1766453.1027038 chr18 1747206 N chr18 1747323 N DEL 13
SRR1766452.2782993 chr18 1747219 N chr18 1747402 N DEL 18
SRR1766467.2550308 chr5 38832207 N chr5 38832338 N DEL 12
SRR1766470.4484859 chr5 38832209 N chr5 38832338 N DEL 13
SRR1766474.7799439 chr5 38832255 N chr5 38832348 N DUP 12
SRR1766456.508299 chr5 38832212 N chr5 38832289 N DEL 10
SRR1766457.5919399 chr5 38832251 N chr5 38832338 N DEL 12
SRR1766472.6618929 chr17 83120066 N chr17 83120165 N DEL 12
SRR1766442.12402026 chr10 6413688 N chr10 6413832 N DEL 14
SRR1766469.7269358 chr10 6413688 N chr10 6413832 N DEL 15
SRR1766477.3440084 chr10 6413686 N chr10 6413883 N DEL 12
SRR1766442.36883666 chr10 6413631 N chr10 6413791 N DEL 11
SRR1766479.7530171 chr10 6413786 N chr10 6413838 N DUP 13
SRR1766474.9353504 chr10 6413686 N chr10 6413883 N DEL 12
SRR1766484.4952826 chr10 6413786 N chr10 6413881 N DUP 13
SRR1766446.8155806 chr10 6413789 N chr10 6413925 N DUP 13
SRR1766462.7981236 chr10 6413786 N chr10 6413881 N DUP 14
SRR1766447.3135905 chr10 6413687 N chr10 6413884 N DEL 13
SRR1766451.6067218 chr10 6413688 N chr10 6413885 N DEL 13
SRR1766482.8213441 chr10 6413690 N chr10 6413887 N DEL 11
SRR1766476.9245016 chr7 112391550 N chr7 112391785 N DEL 10
SRR1766442.24644621 chr7 112391530 N chr7 112392025 N DEL 10
SRR1766474.1414707 chr7 112391668 N chr7 112392059 N DEL 10
SRR1766477.3642909 chr7 112391612 N chr7 112391819 N DUP 15
SRR1766472.5536930 chr7 112391659 N chr7 112392258 N DEL 15
SRR1766443.8510253 chrX 2446459 N chrX 2446947 N DEL 15
SRR1766484.4524200 chrX 2446432 N chrX 2446672 N DEL 11
SRR1766474.5856253 chr16 3062628 N chr16 3063352 N DEL 10
SRR1766449.148659 chr16 3062774 N chr16 3063498 N DEL 17
SRR1766453.2487347 chr9 64773276 N chr9 64773393 N DEL 10
SRR1766463.6339014 chr9 64773482 N chr9 64773754 N DUP 11
SRR1766481.3218934 chr2 70149051 N chr2 70149171 N DEL 12
SRR1766443.10182651 chr3 195710912 N chr3 195711138 N DEL 10
SRR1766455.5079765 chr3 195710833 N chr3 195711237 N DUP 10
SRR1766486.10732033 chr3 195710880 N chr3 195710971 N DEL 10
SRR1766450.10621828 chr3 195710594 N chr3 195710773 N DUP 10
SRR1766457.3462539 chr3 195710507 N chr3 195711574 N DEL 15
SRR1766474.8942288 chr3 195710672 N chr3 195711168 N DEL 18
SRR1766475.5597405 chr3 195710910 N chr3 195711572 N DEL 15
SRR1766448.9376852 chr3 195711152 N chr3 195711376 N DUP 10
SRR1766455.9004478 chr3 195710727 N chr3 195711133 N DEL 10
SRR1766474.1491531 chr3 195710912 N chr3 195711138 N DEL 10
SRR1766460.4964616 chr3 195710427 N chr3 195710516 N DUP 10
SRR1766484.9848909 chr3 195711168 N chr3 195711347 N DUP 10
SRR1766449.5724436 chr3 195710912 N chr3 195711273 N DEL 15
SRR1766483.4753288 chr3 195710745 N chr3 195710881 N DEL 10
SRR1766442.19981783 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766477.10566214 chr3 195710833 N chr3 195711327 N DUP 10
SRR1766465.5826697 chr3 195710594 N chr3 195711223 N DUP 10
SRR1766469.3467702 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766447.7067491 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766455.5079765 chr3 195710475 N chr3 195711286 N DEL 10
SRR1766467.10289914 chr3 195710700 N chr3 195710836 N DEL 18
SRR1766452.6045983 chr3 195710745 N chr3 195711106 N DEL 15
SRR1766442.20460302 chr3 195710746 N chr3 195711330 N DUP 10
SRR1766478.6919910 chr3 195710704 N chr3 195710840 N DEL 10
SRR1766476.5840858 chr3 195711103 N chr3 195711372 N DUP 15
SRR1766442.16760103 chr3 195710653 N chr3 195710967 N DUP 10
SRR1766473.1854743 chr3 195711012 N chr3 195711148 N DEL 15
SRR1766457.9207961 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766481.401328 chr3 195710880 N chr3 195710971 N DEL 10
SRR1766469.3986800 chr3 195710925 N chr3 195711331 N DEL 10
SRR1766450.9305504 chr3 195710913 N chr3 195711227 N DUP 10
SRR1766474.8532251 chr3 195710970 N chr3 195711151 N DEL 15
SRR1766472.4780329 chr3 195710912 N chr3 195711093 N DEL 10
SRR1766442.12486994 chr3 195710672 N chr3 195711213 N DEL 10
SRR1766476.6082131 chr3 195710732 N chr3 195711273 N DEL 10
SRR1766459.9666726 chr3 195710732 N chr3 195711273 N DEL 10
SRR1766470.8672911 chr3 195710656 N chr3 195710745 N DUP 13
SRR1766478.8736120 chr3 195710633 N chr3 195711262 N DUP 12
SRR1766474.7567723 chr3 195711103 N chr3 195711372 N DUP 15
SRR1766444.3503240 chr3 195710722 N chr3 195711308 N DEL 19
SRR1766454.2024097 chr3 195710836 N chr3 195710925 N DUP 12
SRR1766465.553161 chr3 195710970 N chr3 195711106 N DEL 10
SRR1766450.394408 chr3 195710638 N chr3 195711177 N DUP 10
SRR1766473.10829557 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766477.7248460 chr3 195710426 N chr3 195711057 N DEL 10
SRR1766466.6654618 chr3 195711013 N chr3 195711192 N DUP 11
SRR1766479.12475779 chr3 195711088 N chr3 195711357 N DUP 10
SRR1766447.5846248 chr3 195710833 N chr3 195710967 N DUP 11
SRR1766485.5620443 chr3 195710745 N chr3 195710836 N DEL 12
SRR1766462.7946574 chr3 195711182 N chr3 195711273 N DEL 10
SRR1766474.7022316 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766443.4603466 chr3 195710970 N chr3 195711061 N DEL 10
SRR1766455.9004478 chr3 195710427 N chr3 195710741 N DUP 10
SRR1766466.1081679 chr3 195710745 N chr3 195711286 N DEL 19
SRR1766463.7189814 chr3 195710777 N chr3 195711093 N DEL 10
SRR1766474.532605 chr3 195710913 N chr3 195711227 N DUP 10
SRR1766479.8854023 chr3 195710878 N chr3 195711372 N DUP 17
SRR1766463.8865853 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766476.7856287 chr3 195710639 N chr3 195711133 N DUP 10
SRR1766468.5751723 chr3 195710628 N chr3 195710897 N DUP 10
SRR1766449.6616360 chr3 195710833 N chr3 195711192 N DUP 14
SRR1766450.887153 chr3 195711148 N chr3 195711372 N DUP 11
SRR1766447.408951 chr3 195710926 N chr3 195711375 N DUP 15
SRR1766449.6367427 chr3 195710732 N chr3 195711273 N DEL 10
SRR1766459.7609795 chr3 195710777 N chr3 195711093 N DEL 10
SRR1766466.3648164 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766483.75109 chr3 195710913 N chr3 195711227 N DUP 10
SRR1766466.5914983 chr3 195710475 N chr3 195711286 N DEL 10
SRR1766457.8172859 chr3 195711229 N chr3 195711363 N DUP 10
SRR1766486.3483938 chr3 195710913 N chr3 195711227 N DUP 10
SRR1766468.5959020 chr3 195710923 N chr3 195711104 N DEL 10
SRR1766464.3221854 chr3 195711078 N chr3 195711347 N DUP 10
SRR1766479.2256567 chr3 195710652 N chr3 195711283 N DEL 15
SRR1766480.7694544 chr3 195710745 N chr3 195710836 N DEL 10
SRR1766465.8842441 chr3 195710459 N chr3 195711405 N DEL 19
SRR1766467.10289914 chr3 195710862 N chr3 195711268 N DEL 15
SRR1766484.8928592 chr3 195710789 N chr3 195711373 N DUP 10
SRR1766476.2866907 chr3 195710656 N chr3 195710745 N DUP 11
SRR1766448.837598 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766465.553161 chr3 195711140 N chr3 195711319 N DUP 10
SRR1766445.9596139 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766471.169227 chr3 195710868 N chr3 195711182 N DUP 12
SRR1766480.7559984 chr3 195710457 N chr3 195711133 N DEL 10
SRR1766458.189902 chr3 195710727 N chr3 195711133 N DEL 10
SRR1766483.10796568 chr3 195710475 N chr3 195711151 N DEL 10
SRR1766464.8428911 chr3 195710547 N chr3 195710863 N DEL 15
SRR1766460.8663933 chr3 195710911 N chr3 195711137 N DEL 15
SRR1766468.6262396 chr3 195710475 N chr3 195711061 N DEL 14
SRR1766460.6925891 chr3 195711078 N chr3 195711347 N DUP 10
SRR1766463.8588399 chr3 195710898 N chr3 195711032 N DUP 10
SRR1766442.14751536 chr3 195710547 N chr3 195710863 N DEL 15
SRR1766460.10106805 chr3 195710789 N chr3 195711148 N DUP 17
SRR1766450.1336038 chr3 195710745 N chr3 195711286 N DEL 10
SRR1766482.10001994 chr3 195710878 N chr3 195711372 N DUP 10
SRR1766455.2201857 chr3 195711012 N chr3 195711148 N DEL 15
SRR1766485.984262 chr3 195710732 N chr3 195711138 N DEL 10
SRR1766463.7304346 chr3 195710633 N chr3 195711217 N DUP 10
SRR1766449.8188394 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766444.2574313 chr3 195711012 N chr3 195711283 N DEL 10
SRR1766465.5399817 chr3 195710789 N chr3 195711373 N DUP 16
SRR1766482.4252815 chr3 195710652 N chr3 195711103 N DEL 10
SRR1766483.8839114 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766455.781242 chr3 195710833 N chr3 195711237 N DUP 10
SRR1766453.258496 chr3 195710732 N chr3 195710868 N DEL 10
SRR1766447.11282149 chr3 195710926 N chr3 195711105 N DUP 15
SRR1766442.33584866 chr3 195710912 N chr3 195711138 N DEL 15
SRR1766471.11641451 chr3 195710833 N chr3 195711192 N DUP 17
SRR1766478.7676866 chr3 195710897 N chr3 195711123 N DEL 10
SRR1766452.1746923 chr3 195710507 N chr3 195711273 N DEL 10
SRR1766450.887153 chr3 195710912 N chr3 195711273 N DEL 15
SRR1766458.2233427 chr3 195710590 N chr3 195710949 N DUP 17
SRR1766471.11429162 chr3 195711058 N chr3 195711372 N DUP 10
SRR1766485.135474 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766468.3137871 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766470.10029457 chr3 195710779 N chr3 195711363 N DUP 15
SRR1766455.2498048 chr3 195710475 N chr3 195710836 N DEL 10
SRR1766467.2743063 chr3 195710777 N chr3 195711093 N DEL 15
SRR1766469.3750314 chr3 195710745 N chr3 195710881 N DEL 12
SRR1766461.655496 chr3 195710789 N chr3 195711013 N DUP 15
SRR1766442.40725359 chr3 195710907 N chr3 195711133 N DEL 10
SRR1766472.4723707 chr3 195710542 N chr3 195710633 N DEL 15
SRR1766462.10039965 chr3 195710701 N chr3 195711240 N DUP 13
SRR1766460.9110915 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766485.7394197 chr3 195711008 N chr3 195711232 N DUP 10
SRR1766443.4940134 chr3 195710628 N chr3 195710897 N DUP 12
SRR1766484.9848909 chr3 195710832 N chr3 195711238 N DEL 15
SRR1766481.10232930 chr3 195710826 N chr3 195711142 N DEL 10
SRR1766477.11193780 chr3 195710475 N chr3 195711061 N DEL 10
SRR1766467.3593080 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766476.6082131 chr3 195711140 N chr3 195711319 N DUP 10
SRR1766475.11050212 chr3 195710912 N chr3 195711228 N DEL 14
SRR1766474.7596352 chr3 195710735 N chr3 195711141 N DEL 10
SRR1766451.1034834 chr3 195710511 N chr3 195711142 N DEL 10
SRR1766480.8347394 chr3 195710912 N chr3 195711138 N DEL 15
SRR1766482.5996566 chr3 195710912 N chr3 195711273 N DEL 15
SRR1766468.5127411 chr3 195710746 N chr3 195711240 N DUP 14
SRR1766442.29999421 chr3 195710475 N chr3 195711061 N DEL 10
SRR1766478.8736120 chr3 195710652 N chr3 195711148 N DEL 10
SRR1766442.22842530 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766479.10878674 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766481.808784 chr3 195710626 N chr3 195711165 N DUP 10
SRR1766442.44460459 chr3 195710745 N chr3 195711286 N DEL 15
SRR1766442.44343984 chr3 195710998 N chr3 195711087 N DUP 10
SRR1766475.6189519 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766482.8002010 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766483.6659795 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766467.8598360 chr3 195711078 N chr3 195711347 N DUP 10
SRR1766477.2482102 chr3 195710833 N chr3 195711192 N DUP 12
SRR1766474.9856445 chr3 195711103 N chr3 195711372 N DUP 15
SRR1766457.7812382 chr3 195711023 N chr3 195711202 N DUP 11
SRR1766477.7248460 chr3 195710673 N chr3 195711167 N DUP 14
SRR1766457.6375563 chr3 195710745 N chr3 195711061 N DEL 10
SRR1766459.6172648 chr3 195710656 N chr3 195710745 N DUP 10
SRR1766458.6590782 chr3 195710728 N chr3 195710819 N DEL 19
SRR1766463.8429951 chr3 195710633 N chr3 195711262 N DUP 14
SRR1766479.4039026 chr3 195710431 N chr3 195711150 N DUP 10
SRR1766477.937789 chr3 195710701 N chr3 195711195 N DUP 10
SRR1766457.1670099 chr3 195711023 N chr3 195711202 N DUP 11
SRR1766453.7617469 chr3 195711013 N chr3 195711192 N DUP 10
SRR1766477.5150813 chr3 195710537 N chr3 195710853 N DEL 10
SRR1766471.5020912 chr3 195710789 N chr3 195711373 N DUP 10
SRR1766468.6262396 chr3 195710907 N chr3 195711133 N DEL 12
SRR1766443.6423575 chr3 195710547 N chr3 195710863 N DEL 15
SRR1766461.214453 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766470.635997 chr3 195710925 N chr3 195711061 N DEL 10
SRR1766473.6701931 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766451.7364049 chr3 195710897 N chr3 195711213 N DEL 10
SRR1766472.6537572 chr3 195710925 N chr3 195711331 N DEL 10
SRR1766467.2489668 chr3 195711058 N chr3 195711372 N DUP 10
SRR1766467.6409670 chr3 195710907 N chr3 195711133 N DEL 15
SRR1766471.169227 chr3 195710548 N chr3 195711089 N DEL 12
SRR1766463.3808006 chr3 195710833 N chr3 195711237 N DUP 11
SRR1766475.10734632 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766467.11909659 chr3 195710459 N chr3 195711405 N DEL 19
SRR1766447.408951 chr3 195710878 N chr3 195711012 N DUP 10
SRR1766485.3535942 chr3 195710836 N chr3 195710970 N DUP 17
SRR1766472.2927865 chr3 195710656 N chr3 195710745 N DUP 11
SRR1766455.8921189 chr3 195710745 N chr3 195711331 N DEL 10
SRR1766475.11201508 chr3 195710732 N chr3 195711093 N DEL 10
SRR1766466.6347383 chr3 195710626 N chr3 195711210 N DUP 13
SRR1766453.934597 chr3 195710907 N chr3 195711133 N DEL 11
SRR1766472.7658271 chr3 195710672 N chr3 195711168 N DEL 11
SRR1766445.6863892 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766459.5970256 chr3 195710475 N chr3 195711061 N DEL 10
SRR1766485.4252295 chr3 195710475 N chr3 195711151 N DEL 10
SRR1766477.4833033 chr3 195710833 N chr3 195710922 N DUP 17
SRR1766482.7511894 chr3 195710595 N chr3 195711406 N DEL 10
SRR1766467.7695697 chr3 195711048 N chr3 195711362 N DUP 10
SRR1766470.1238586 chr3 195710457 N chr3 195711133 N DEL 10
SRR1766442.44460459 chr3 195710788 N chr3 195710879 N DEL 15
SRR1766453.6263591 chr3 195710590 N chr3 195710814 N DUP 15
SRR1766456.6505169 chr3 195710886 N chr3 195711020 N DUP 10
SRR1766481.401328 chr3 195711048 N chr3 195711362 N DUP 10
SRR1766442.36079111 chr3 195710454 N chr3 195710590 N DEL 10
SRR1766444.2118210 chr3 195710427 N chr3 195711236 N DUP 10
SRR1766484.2346909 chr3 195710652 N chr3 195711058 N DEL 10
SRR1766454.4427009 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766484.2182020 chr3 195710898 N chr3 195710987 N DUP 14
SRR1766442.29532329 chr3 195711452 N chr3 195711619 N DEL 10
SRR1766447.4999222 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766442.24904724 chr3 195711140 N chr3 195711319 N DUP 10
SRR1766463.9254572 chr3 195710475 N chr3 195711061 N DEL 10
SRR1766481.3123362 chr3 195710459 N chr3 195711405 N DEL 19
SRR1766469.10933803 chr3 195710897 N chr3 195711123 N DEL 10
SRR1766454.5799610 chr3 195710701 N chr3 195711150 N DUP 15
SRR1766477.6908917 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766446.4027275 chr3 195710897 N chr3 195711258 N DEL 10
SRR1766449.9872863 chr3 195710745 N chr3 195711106 N DEL 10
SRR1766451.1444838 chr3 195710833 N chr3 195711327 N DUP 10
SRR1766474.3832772 chr3 195711355 N chr3 195711477 N DEL 11
SRR1766467.1984014 chr3 195710732 N chr3 195711273 N DEL 10
SRR1766467.3277409 chr3 195710457 N chr3 195711133 N DEL 13
SRR1766485.10768266 chr3 195710912 N chr3 195711273 N DEL 13
SRR1766442.46715952 chr3 195710789 N chr3 195711013 N DUP 11
SRR1766474.10077014 chr3 195711452 N chr3 195711619 N DEL 10
SRR1766456.3324189 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766459.7117162 chr3 195710745 N chr3 195710881 N DEL 11
SRR1766455.3351269 chr3 195710907 N chr3 195711133 N DEL 15
SRR1766480.5745705 chr3 195710624 N chr3 195711030 N DEL 10
SRR1766464.4828612 chr3 195710833 N chr3 195711192 N DUP 16
SRR1766446.3366022 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766462.493625 chr3 195710475 N chr3 195710656 N DEL 10
SRR1766472.6838449 chr3 195710878 N chr3 195711012 N DUP 10
SRR1766470.3593366 chr3 195710916 N chr3 195711097 N DEL 10
SRR1766450.7953199 chr3 195710672 N chr3 195711168 N DEL 10
SRR1766471.11163655 chr3 195710653 N chr3 195711192 N DUP 10
SRR1766449.8359246 chr3 195710925 N chr3 195711286 N DEL 10
SRR1766454.8857819 chr3 195710867 N chr3 195711048 N DEL 15
SRR1766470.5933755 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766442.43840210 chr3 195711078 N chr3 195711347 N DUP 10
SRR1766448.9248612 chr3 195710672 N chr3 195711168 N DEL 10
SRR1766474.3832772 chr3 195711360 N chr3 195711572 N DEL 13
SRR1766455.5643578 chr3 195710742 N chr3 195711013 N DEL 10
SRR1766446.7445980 chr3 195711183 N chr3 195711409 N DEL 15
SRR1766464.1659129 chr3 195710700 N chr3 195710836 N DEL 15
SRR1766473.2465703 chr3 195710878 N chr3 195711012 N DUP 10
SRR1766485.12053858 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766478.5473077 chr3 195710682 N chr3 195711133 N DEL 10
SRR1766472.9674977 chr3 195710643 N chr3 195711272 N DUP 10
SRR1766454.535141 chr3 195710925 N chr3 195711151 N DEL 10
SRR1766442.21983193 chr3 195710619 N chr3 195711158 N DUP 10
SRR1766473.10023160 chr3 195711012 N chr3 195711148 N DEL 16
SRR1766467.9978162 chr3 195710517 N chr3 195710833 N DEL 15
SRR1766472.3839632 chr3 195710628 N chr3 195711347 N DUP 15
SRR1766442.12466967 chr3 195710507 N chr3 195711408 N DEL 12
SRR1766469.3711865 chr3 195710542 N chr3 195710633 N DEL 10
SRR1766465.1693275 chr3 195710700 N chr3 195710836 N DEL 10
SRR1766442.44332938 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766486.7315157 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766457.8737280 chr3 195710897 N chr3 195711258 N DEL 10
SRR1766462.9596106 chr3 195710833 N chr3 195711237 N DUP 10
SRR1766448.4758028 chr3 195711058 N chr3 195711372 N DUP 10
SRR1766465.8004613 chr3 195710480 N chr3 195710661 N DEL 10
SRR1766444.4464954 chr14 64895053 N chr14 64895178 N DUP 12
SRR1766470.3710924 chr1 79571577 N chr1 79571638 N DEL 11
SRR1766483.9491342 chr1 79571577 N chr1 79571638 N DEL 12
SRR1766462.2485562 chr1 79571577 N chr1 79571638 N DEL 18
SRR1766447.9312595 chr1 79571577 N chr1 79571638 N DEL 18
SRR1766468.2163352 chr1 79571577 N chr1 79571638 N DEL 11
SRR1766471.5590163 chr1 79571738 N chr1 79572271 N DEL 11
SRR1766451.6894104 chr1 79571738 N chr1 79572271 N DEL 11
SRR1766442.34987791 chr1 79571818 N chr1 79572324 N DEL 12
SRR1766442.34633864 chr1 79571738 N chr1 79572271 N DEL 13
SRR1766471.11304270 chr1 79571546 N chr1 79572271 N DEL 13
SRR1766468.4178449 chr1 79571546 N chr1 79572271 N DEL 13
SRR1766459.9780871 chr1 79571546 N chr1 79572271 N DEL 13
SRR1766448.10726856 chr9 90694423 N chr9 90694568 N DEL 10
SRR1766484.11213057 chr9 90694623 N chr9 90694744 N DUP 10
SRR1766474.4940835 chr9 90694646 N chr9 90694824 N DUP 11
SRR1766479.13054677 chr9 90694440 N chr9 90694848 N DEL 12
SRR1766454.76778 chr8 138805414 N chr8 138805682 N DEL 13
SRR1766480.1881716 chr8 138805448 N chr8 138805740 N DEL 12
SRR1766486.7169460 chr8 138805175 N chr8 138805798 N DEL 10
SRR1766446.9095398 chr8 138805054 N chr8 138805994 N DUP 10
SRR1766480.4933065 chr8 138805462 N chr8 138805968 N DEL 12
SRR1766449.6096411 chr8 138805315 N chr8 138806197 N DUP 14
SRR1766482.4581115 chr8 138805094 N chr8 138806180 N DEL 19
SRR1766442.6216434 chr8 138805147 N chr8 138806181 N DEL 10
SRR1766461.361097 chr8 138806218 N chr8 138806279 N DEL 17
SRR1766478.10005766 chr8 138806005 N chr8 138806287 N DUP 11
SRR1766480.679171 chr8 138806199 N chr8 138806308 N DUP 14
SRR1766468.4190891 chr8 138805441 N chr8 138806328 N DEL 15
SRR1766479.7239807 chr8 138806070 N chr8 138806329 N DEL 10
SRR1766459.5658021 chr8 138805088 N chr8 138806366 N DEL 10
SRR1766483.272223 chr8 138805780 N chr8 138806364 N DEL 15
SRR1766442.32097664 chr16 9676239 N chr16 9676324 N DEL 10
SRR1766477.5740264 chr16 9676241 N chr16 9676326 N DEL 10
SRR1766442.37291015 chr22 18387819 N chr22 18389317 N DEL 14
SRR1766478.1374096 chr22 18387819 N chr22 18389317 N DEL 13
SRR1766451.5862318 chr22 18387815 N chr22 18389190 N DEL 12
SRR1766480.3894290 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766461.10893418 chr22 18387821 N chr22 18389216 N DEL 16
SRR1766449.6324853 chr22 18387753 N chr22 18388498 N DUP 11
SRR1766463.10308022 chr22 18387821 N chr22 18389216 N DEL 16
SRR1766454.5110384 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766449.6285817 chr22 18387821 N chr22 18389216 N DEL 16
SRR1766442.6786160 chr22 18387819 N chr22 18389317 N DEL 13
SRR1766486.2857285 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766459.3491401 chr22 18387819 N chr22 18389317 N DEL 13
SRR1766486.5100544 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766464.10167303 chr22 18387819 N chr22 18389317 N DEL 13
SRR1766442.627522 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766459.8404462 chr22 18388339 N chr22 18389057 N DUP 12
SRR1766485.9898568 chr22 18387821 N chr22 18389216 N DEL 16
SRR1766462.295527 chr22 18387821 N chr22 18389216 N DEL 17
SRR1766466.9704657 chr22 18387815 N chr22 18389190 N DEL 12
SRR1766467.4444426 chr12 58598054 N chr12 58598123 N DEL 11
SRR1766483.2597789 chr12 58598058 N chr12 58598127 N DEL 11
SRR1766471.9749542 chr8 502871 N chr8 503915 N DEL 10
SRR1766469.6440352 chr8 502890 N chr8 503881 N DEL 15
SRR1766476.9458167 chr8 502747 N chr8 502905 N DUP 10
SRR1766484.1851163 chr8 502898 N chr8 503889 N DEL 15
SRR1766468.411684 chr8 502914 N chr8 503956 N DUP 10
SRR1766451.7719733 chr8 502860 N chr8 502914 N DEL 10
SRR1766478.6657668 chr8 502754 N chr8 502914 N DEL 13
SRR1766452.3233212 chr8 502868 N chr8 503079 N DUP 10
SRR1766453.3917157 chr8 502745 N chr8 503062 N DUP 15
SRR1766474.7086772 chr8 503083 N chr8 503913 N DUP 15
SRR1766474.8472392 chr8 503209 N chr8 503582 N DEL 11
SRR1766469.3854778 chr8 503201 N chr8 503874 N DEL 10
SRR1766454.4203599 chr8 503201 N chr8 503874 N DEL 10
SRR1766483.7222789 chr8 502840 N chr8 503159 N DEL 10
SRR1766455.7355902 chr8 503183 N chr8 503607 N DUP 10
SRR1766456.3322045 chr8 503108 N chr8 503268 N DEL 15
SRR1766475.2914781 chr8 502842 N chr8 503214 N DEL 10
SRR1766470.8872816 chr8 502764 N chr8 503295 N DEL 14
SRR1766483.5664643 chr8 503304 N chr8 503922 N DUP 10
SRR1766478.1782770 chr8 503400 N chr8 504020 N DEL 10
SRR1766476.2152719 chr8 502745 N chr8 503487 N DUP 11
SRR1766473.5118661 chr8 502978 N chr8 503508 N DUP 10
SRR1766486.2540170 chr8 503467 N chr8 504085 N DUP 10
SRR1766473.9919515 chr8 502778 N chr8 503522 N DEL 10
SRR1766450.1299375 chr8 502778 N chr8 503522 N DEL 10
SRR1766448.4247165 chr8 502725 N chr8 503575 N DEL 19
SRR1766455.8063520 chr8 503765 N chr8 503905 N DUP 10
SRR1766445.6372168 chr8 503037 N chr8 503975 N DEL 12
SRR1766478.3420881 chr8 503791 N chr8 504093 N DEL 10
SRR1766486.5961332 chr8 503957 N chr8 504118 N DEL 15
SRR1766474.5890640 chr8 503958 N chr8 504119 N DEL 17
SRR1766474.2170047 chr6 21924857 N chr6 21925146 N DEL 10
SRR1766457.2101709 chr12 132533240 N chr12 132533435 N DEL 15
SRR1766447.10099578 chr19 14314284 N chr19 14314435 N DEL 10
SRR1766460.7025797 chr9 134729779 N chr9 134729880 N DUP 15
SRR1766451.8778622 chr4 110267179 N chr4 110267313 N DEL 10
SRR1766455.4441729 chr16 938438 N chr16 938605 N DEL 10
SRR1766460.2212240 chr20 51961825 N chr20 51961881 N DEL 17
SRR1766484.8808183 chr20 51961808 N chr20 51961869 N DUP 13
SRR1766448.9185081 chr20 51961808 N chr20 51961869 N DUP 14
SRR1766478.4537233 chr20 51961808 N chr20 51961869 N DUP 11
SRR1766482.5816062 chr20 51961860 N chr20 51961918 N DEL 13
SRR1766445.5371765 chr20 51961860 N chr20 51961918 N DEL 14
SRR1766442.12650950 chr20 51961827 N chr20 51961918 N DEL 12
SRR1766481.9655942 chr5 139446617 N chr5 139446678 N DUP 16
SRR1766469.4138406 chr21 30210368 N chr21 30210452 N DEL 18
SRR1766442.23746175 chr21 30210368 N chr21 30210452 N DEL 18
SRR1766474.3070299 chr21 30210368 N chr21 30210452 N DEL 18
SRR1766460.2600477 chr21 30210328 N chr21 30210459 N DUP 11
SRR1766442.26075966 chr21 30210443 N chr21 30210505 N DEL 11
SRR1766477.5122969 chr21 30210443 N chr21 30210505 N DEL 11
SRR1766442.47170639 chr21 30210441 N chr21 30210505 N DEL 13
SRR1766472.5054308 chr1 152910467 N chr1 152910676 N DUP 15
SRR1766474.2656039 chr1 152910467 N chr1 152910586 N DUP 10
SRR1766475.4591905 chr1 152910598 N chr1 152910959 N DEL 10
SRR1766470.4229988 chr1 152910467 N chr1 152910676 N DUP 12
SRR1766476.2082186 chr1 152910718 N chr1 152910959 N DEL 10
SRR1766442.6346928 chr1 152910725 N chr1 152910876 N DEL 10
SRR1766469.1778429 chr1 152910722 N chr1 152910963 N DEL 10
SRR1766461.10997945 chr1 152910702 N chr1 152910943 N DEL 18
SRR1766473.7020687 chr1 152910460 N chr1 152910579 N DUP 10
SRR1766482.10614598 chr1 152910812 N chr1 152910963 N DEL 10
SRR1766442.8667672 chr1 152910468 N chr1 152910857 N DUP 14
SRR1766443.2486898 chr1 152910474 N chr1 152910833 N DUP 15
SRR1766485.8810549 chr1 152910808 N chr1 152910897 N DUP 10
SRR1766468.2904263 chr1 152910904 N chr1 152911085 N DEL 12
SRR1766467.9626364 chr1 152910495 N chr1 152910856 N DEL 18
SRR1766483.2051446 chr1 152910545 N chr1 152910876 N DEL 15
SRR1766442.34098364 chr1 152910515 N chr1 152910876 N DEL 18
SRR1766455.6899229 chr1 152910916 N chr1 152911005 N DUP 10
SRR1766468.2073554 chr1 152910492 N chr1 152910943 N DEL 10
SRR1766477.438229 chr1 152910474 N chr1 152911013 N DUP 15
SRR1766447.6054186 chr1 152910510 N chr1 152910961 N DEL 17
SRR1766451.6599576 chr1 152910500 N chr1 152911071 N DEL 14
SRR1766477.8541968 chr1 152910498 N chr1 152911099 N DEL 10
SRR1766483.3118710 chr1 152911016 N chr1 152911137 N DEL 16
SRR1766481.13058358 chr1 152910988 N chr1 152911139 N DEL 10
SRR1766473.1929648 chr1 152910986 N chr1 152911137 N DEL 10
SRR1766455.6368920 chr1 152911003 N chr1 152911205 N DEL 10
SRR1766444.126691 chr1 152911161 N chr1 152911513 N DEL 12
SRR1766480.5367214 chr8 53948069 N chr8 53948492 N DEL 10
SRR1766458.4485813 chr8 53948469 N chr8 53948534 N DEL 12
SRR1766442.3697057 chr8 53948546 N chr8 53948702 N DUP 19
SRR1766457.1535324 chr8 53948546 N chr8 53948702 N DUP 15
SRR1766484.975708 chr8 53948681 N chr8 53948775 N DEL 10
SRR1766451.734687 chr8 53948694 N chr8 53949379 N DEL 19
SRR1766474.8039837 chr8 53948546 N chr8 53948671 N DUP 14
SRR1766443.2383968 chr8 53948546 N chr8 53948671 N DUP 14
SRR1766483.1400840 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766459.4283077 chr8 53948546 N chr8 53948702 N DUP 10
SRR1766443.3007941 chr8 53948546 N chr8 53948671 N DUP 14
SRR1766472.10061483 chr8 53948546 N chr8 53948702 N DUP 12
SRR1766480.5367214 chr8 53948546 N chr8 53948702 N DUP 12
SRR1766471.3337781 chr8 53948546 N chr8 53948702 N DUP 15
SRR1766477.10730121 chr8 53948681 N chr8 53948775 N DEL 14
SRR1766451.10491113 chr8 53948579 N chr8 53948640 N DUP 10
SRR1766482.3077480 chr8 53948546 N chr8 53948702 N DUP 18
SRR1766459.7983865 chr8 53948546 N chr8 53948671 N DUP 14
SRR1766472.6925159 chr8 53948681 N chr8 53948775 N DEL 14
SRR1766472.3520083 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766478.7083075 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766477.7993044 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766453.6186332 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766486.8335902 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766451.9742482 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766458.6096115 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766467.3611520 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766452.9734761 chr8 53948635 N chr8 53949039 N DEL 10
SRR1766479.524443 chr8 53948635 N chr8 53949039 N DEL 12
SRR1766442.11481844 chr8 53948813 N chr8 53949469 N DUP 10
SRR1766472.3450154 chr8 53948568 N chr8 53948790 N DEL 10
SRR1766460.5722005 chr8 53949349 N chr8 53949414 N DUP 15
SRR1766442.3386806 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766454.3170456 chr8 53949349 N chr8 53949414 N DUP 16
SRR1766475.6495258 chr8 53949349 N chr8 53949414 N DUP 18
SRR1766485.4518706 chr8 53949349 N chr8 53949414 N DUP 18
SRR1766442.26590434 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766443.2522726 chr8 53949349 N chr8 53949414 N DUP 18
SRR1766482.3077480 chr8 53949349 N chr8 53949414 N DUP 18
SRR1766486.11420708 chr8 53949349 N chr8 53949414 N DUP 17
SRR1766451.10491113 chr8 53949349 N chr8 53949414 N DUP 15
SRR1766479.1620539 chr8 53949349 N chr8 53949414 N DUP 15
SRR1766470.2756996 chr8 53949349 N chr8 53949414 N DUP 16
SRR1766465.9141214 chr8 53949349 N chr8 53949414 N DUP 17
SRR1766451.32847 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766451.3859206 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766474.8039837 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766481.11739291 chr8 53949193 N chr8 53949382 N DEL 12
SRR1766465.5298271 chr8 53949193 N chr8 53949382 N DEL 12
SRR1766472.3378987 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766448.8703754 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766478.3222391 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766452.5856556 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766458.6502372 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766481.6853877 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766442.39466710 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766455.4331222 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766476.5927921 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766460.8989042 chr8 53948503 N chr8 53949382 N DEL 12
SRR1766478.231747 chr8 53947542 N chr8 53949383 N DEL 12
SRR1766442.2788552 chr8 53947544 N chr8 53949385 N DEL 12
SRR1766473.3207979 chr3 68370513 N chr3 68370588 N DUP 13
SRR1766463.4837440 chr3 68370481 N chr3 68370544 N DUP 10
SRR1766475.4698443 chr1 193564152 N chr1 193564215 N DUP 18
SRR1766473.10071648 chr1 193564152 N chr1 193564215 N DUP 18
SRR1766442.25832369 chr1 193564152 N chr1 193564215 N DUP 18
SRR1766486.4843192 chr1 193564094 N chr1 193564157 N DUP 14
SRR1766483.11307293 chr1 193564152 N chr1 193564215 N DUP 17
SRR1766485.7714912 chr1 193564152 N chr1 193564215 N DUP 10
SRR1766451.4404855 chr1 193564152 N chr1 193564215 N DUP 11
SRR1766447.11444853 chr1 193564108 N chr1 193564235 N DEL 13
SRR1766457.8214793 chr1 193564109 N chr1 193564236 N DEL 12
SRR1766450.3142331 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766442.4206423 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766463.6903386 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766466.6520294 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766482.4059033 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766455.6058643 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766483.9242974 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766473.7538231 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766478.85808 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766485.11068888 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766464.7524560 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766476.8699710 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766442.36381810 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766472.8079996 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766477.6387356 chr1 193564454 N chr1 193564513 N DUP 12
SRR1766451.7150110 chr1 193564447 N chr1 193564506 N DUP 10
SRR1766482.7926549 chr1 193564447 N chr1 193564506 N DUP 10
SRR1766454.10975702 chr1 193564454 N chr1 193564513 N DUP 11
SRR1766473.7800479 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766485.11732669 chr1 193564447 N chr1 193564506 N DUP 10
SRR1766442.12520589 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766474.8652019 chr1 193564447 N chr1 193564506 N DUP 11
SRR1766476.5950297 chr4 47123656 N chr4 47123728 N DEL 10
SRR1766466.8043261 chr4 47123656 N chr4 47123728 N DEL 11
SRR1766481.6991814 chr4 47123656 N chr4 47123728 N DEL 12
SRR1766458.6776830 chr4 47123656 N chr4 47123728 N DEL 16
SRR1766462.5339398 chr4 47123656 N chr4 47123728 N DEL 16
SRR1766473.7989262 chr4 47123656 N chr4 47123728 N DEL 16
SRR1766461.7605809 chr4 47123591 N chr4 47123729 N DEL 14
SRR1766442.5011230 chr4 47123591 N chr4 47123729 N DEL 14
SRR1766447.8537721 chr4 47123615 N chr4 47123731 N DEL 12
SRR1766479.3554254 chr4 47123616 N chr4 47123732 N DEL 11
SRR1766447.2263748 chr4 47123616 N chr4 47123732 N DEL 11
SRR1766486.7116022 chr7 98548101 N chr7 98548218 N DEL 10
SRR1766466.2612322 chr7 98548115 N chr7 98548360 N DEL 10
SRR1766460.11162023 chr7 98548043 N chr7 98548146 N DUP 10
SRR1766461.6444505 chr7 98548147 N chr7 98548220 N DEL 10
SRR1766442.13887972 chr7 98548164 N chr7 98548669 N DEL 10
SRR1766461.9124717 chr7 98548157 N chr7 98548598 N DEL 15
SRR1766486.6817236 chr7 98548163 N chr7 98548768 N DEL 14
SRR1766442.27465266 chr7 98548139 N chr7 98548224 N DEL 15
SRR1766448.71091 chr7 98548139 N chr7 98548224 N DEL 15
SRR1766458.9403477 chr7 98548212 N chr7 98548309 N DEL 14
SRR1766442.5942859 chr7 98548148 N chr7 98548243 N DUP 10
SRR1766477.383737 chr7 98548043 N chr7 98548242 N DUP 10
SRR1766470.5566145 chr7 98548268 N chr7 98548329 N DEL 10
SRR1766483.169293 chr7 98548200 N chr7 98548703 N DUP 17
SRR1766471.11487128 chr7 98548208 N chr7 98548263 N DUP 14
SRR1766442.40470313 chr7 98548220 N chr7 98548283 N DUP 12
SRR1766466.4977195 chr7 98548186 N chr7 98548645 N DUP 17
SRR1766471.630374 chr7 98548186 N chr7 98548645 N DUP 16
SRR1766453.720103 chr7 98548296 N chr7 98548765 N DEL 16
SRR1766463.8036211 chr7 98548267 N chr7 98548344 N DEL 18
SRR1766446.8319032 chr7 98548045 N chr7 98548304 N DUP 12
SRR1766484.3714467 chr7 98548322 N chr7 98548771 N DEL 12
SRR1766453.5406955 chr7 98548221 N chr7 98548324 N DUP 10
SRR1766466.8379930 chr7 98548190 N chr7 98548301 N DUP 10
SRR1766481.6867636 chr7 98548211 N chr7 98548326 N DUP 14
SRR1766467.6559650 chr7 98548219 N chr7 98548350 N DUP 10
SRR1766457.5098205 chr7 98548200 N chr7 98548335 N DUP 12
SRR1766470.10609240 chr7 98548376 N chr7 98548749 N DEL 17
SRR1766458.8643213 chr7 98548395 N chr7 98548756 N DEL 10
SRR1766478.10878121 chr7 98548262 N chr7 98548347 N DEL 10
SRR1766481.11251140 chr7 98548244 N chr7 98548309 N DEL 11
SRR1766481.4296496 chr7 98548247 N chr7 98548332 N DEL 18
SRR1766467.6559650 chr7 98548162 N chr7 98548339 N DEL 10
SRR1766448.4562121 chr7 98548200 N chr7 98548407 N DUP 18
SRR1766462.5733748 chr7 98548244 N chr7 98548381 N DEL 15
SRR1766486.5726415 chr7 98548358 N chr7 98548441 N DUP 15
SRR1766451.6047935 chr7 98548488 N chr7 98548765 N DEL 13
SRR1766476.9806805 chr7 98548085 N chr7 98548484 N DUP 14
SRR1766478.5194205 chr7 98548043 N chr7 98548522 N DUP 13
SRR1766442.25488686 chr7 98548420 N chr7 98548523 N DUP 12
SRR1766442.6855979 chr7 98548248 N chr7 98548473 N DEL 18
SRR1766452.4814280 chr7 98548245 N chr7 98548466 N DEL 15
SRR1766484.2043011 chr7 98548472 N chr7 98548583 N DUP 15
SRR1766460.4659647 chr7 98548106 N chr7 98548569 N DUP 10
SRR1766464.7088058 chr7 98548143 N chr7 98548564 N DEL 15
SRR1766442.4903226 chr7 98548423 N chr7 98548674 N DUP 14
SRR1766452.2820528 chr7 98548488 N chr7 98548557 N DEL 15
SRR1766476.7130305 chr7 98548240 N chr7 98548589 N DEL 15
SRR1766462.7628201 chr7 98548106 N chr7 98548701 N DUP 10
SRR1766453.3469609 chr7 98548144 N chr7 98548627 N DUP 12
SRR1766443.5165035 chr7 98548124 N chr7 98548669 N DEL 10
SRR1766485.4716558 chr20 33115584 N chr20 33115740 N DEL 10
SRR1766472.1075631 chr8 72573698 N chr8 72573859 N DEL 15
SRR1766458.4594203 chr19 51944740 N chr19 51944993 N DEL 15
SRR1766480.6838663 chr19 51944794 N chr19 51945047 N DEL 18
SRR1766442.4047295 chr11 129671829 N chr11 129672176 N DEL 16
SRR1766462.7016405 chr11 129671834 N chr11 129672181 N DEL 10
SRR1766462.4809574 chr3 122252489 N chr3 122252560 N DEL 10
SRR1766457.6889164 chr6 59360836 N chr6 59361004 N DUP 10
SRR1766453.4173298 chr6 59360818 N chr6 59360986 N DUP 10
SRR1766442.21498640 chr11 131265291 N chr11 131265465 N DEL 15
SRR1766472.10859752 chr11 131265291 N chr11 131265465 N DEL 15
SRR1766451.10489424 chr11 131265291 N chr11 131265465 N DEL 16
SRR1766442.15356765 chr11 131265291 N chr11 131265465 N DEL 17
SRR1766465.2138958 chr11 131265291 N chr11 131265465 N DEL 17
SRR1766442.861060 chr11 131265291 N chr11 131265465 N DEL 17
SRR1766467.5413266 chr11 131265368 N chr11 131265417 N DUP 11
SRR1766481.234453 chr11 131265352 N chr11 131265544 N DUP 11
SRR1766468.2007970 chr4 15733383 N chr4 15733532 N DEL 18
SRR1766442.42863461 chr11 70119163 N chr11 70119388 N DUP 10
SRR1766483.7050024 chr11 70119432 N chr11 70119632 N DEL 10
SRR1766454.6137843 chr7 50459722 N chr7 50459916 N DEL 10
SRR1766481.2162972 chrX 120374757 N chrX 120374845 N DEL 17
SRR1766452.107015 chrX 120374810 N chrX 120374920 N DUP 15
SRR1766451.294699 chrX 120374788 N chrX 120374910 N DUP 16
SRR1766485.4373049 chrX 120374696 N chrX 120374907 N DEL 16
SRR1766450.10847777 chrX 54065345 N chrX 54065860 N DEL 10
SRR1766484.7672051 chr20 36976512 N chr20 36976860 N DUP 12
SRR1766447.1968733 chr20 36976512 N chr20 36976860 N DUP 12
SRR1766473.4263025 chr8 38508022 N chr8 38508089 N DEL 12
SRR1766469.6961169 chr8 38508008 N chr8 38508090 N DEL 14
SRR1766449.8636484 chr17 72189542 N chr17 72189697 N DUP 14
SRR1766472.2440465 chr9 43337167 N chr9 43337241 N DUP 12
SRR1766460.5617959 chr6 157870610 N chr6 157870819 N DUP 10
SRR1766466.6142338 chr10 27296559 N chr10 27296783 N DUP 15
SRR1766476.10091523 chr10 27296590 N chr10 27296716 N DUP 10
SRR1766482.980916 chr4 43451137 N chr4 43451231 N DEL 14
SRR1766442.27703620 chr4 43450920 N chr4 43451088 N DEL 10
SRR1766442.43901911 chr6 22836799 N chr6 22836928 N DEL 10
SRR1766457.769618 chr6 22836727 N chr6 22837030 N DUP 10
SRR1766474.6762309 chr6 22836737 N chr6 22837089 N DUP 10
SRR1766464.6026045 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766460.1982169 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766453.7066482 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766442.12203348 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766451.6880040 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766447.2945355 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766453.6237945 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766450.1838200 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766460.8339405 chr9 43321830 N chr9 43321923 N DUP 14
SRR1766472.5866829 chr9 43321846 N chr9 43321897 N DUP 10
SRR1766483.669286 chr9 43321798 N chr9 43321849 N DUP 11
SRR1766470.2513747 chr9 43321843 N chr9 43321894 N DUP 11
SRR1766453.5350190 chr9 43321843 N chr9 43321894 N DUP 12
SRR1766452.7524072 chr1 2960156 N chr1 2960247 N DEL 10
SRR1766471.10812301 chr1 2960156 N chr1 2960247 N DEL 10
SRR1766465.1854512 chr1 2960156 N chr1 2960277 N DEL 12
SRR1766482.4026133 chr1 2960156 N chr1 2960277 N DEL 12
SRR1766443.1192417 chr1 2960156 N chr1 2960277 N DEL 13
SRR1766470.8564719 chr1 2960156 N chr1 2960277 N DEL 15
SRR1766479.9203261 chr1 2960156 N chr1 2960277 N DEL 15
SRR1766466.6253184 chr1 2960156 N chr1 2960277 N DEL 14
SRR1766468.3661359 chr2 3844467 N chr2 3844526 N DUP 10
SRR1766453.829135 chr10 42171825 N chr10 42171966 N DEL 10
SRR1766472.11835266 chr11 62962001 N chr11 62962302 N DEL 19
SRR1766442.6779404 chr11 62962001 N chr11 62962302 N DEL 10
SRR1766478.3257918 chr6 4895431 N chr6 4895506 N DUP 16
SRR1766462.885501 chr15 57075906 N chr15 57075980 N DUP 12
SRR1766474.4160485 chr15 57075906 N chr15 57075980 N DUP 12
SRR1766471.436829 chr15 57075906 N chr15 57075980 N DUP 13
SRR1766474.9860200 chr15 57075924 N chr15 57075986 N DEL 14
SRR1766476.806376 chr2 197473565 N chr2 197473642 N DUP 15
SRR1766450.8830998 chr15 65864211 N chr15 65864551 N DEL 11
SRR1766451.5135594 chr15 65864193 N chr15 65864623 N DEL 11
SRR1766484.10435606 chr15 65864193 N chr15 65864623 N DEL 11
SRR1766484.9713825 chr6 169923983 N chr6 169924381 N DUP 16
SRR1766478.10214154 chr6 169923983 N chr6 169924381 N DUP 16
SRR1766469.5036537 chr6 169923983 N chr6 169924381 N DUP 12
SRR1766463.3411238 chr6 169923983 N chr6 169924381 N DUP 11
SRR1766479.5250248 chr6 169923959 N chr6 169924141 N DUP 14
SRR1766473.11177425 chr6 169923954 N chr6 169924136 N DUP 10
SRR1766485.449032 chr6 169924065 N chr6 169924283 N DUP 16
SRR1766455.6704533 chr6 169924033 N chr6 169924140 N DUP 18
SRR1766458.1423171 chr6 169923954 N chr6 169924136 N DUP 16
SRR1766445.2206256 chr6 169924033 N chr6 169924140 N DUP 18
SRR1766462.1454658 chr6 169923954 N chr6 169924136 N DUP 17
SRR1766456.3733458 chr6 169923954 N chr6 169924136 N DUP 17
SRR1766467.6218822 chr6 169923954 N chr6 169924136 N DUP 17
SRR1766477.7915747 chr6 169923959 N chr6 169924141 N DUP 17
SRR1766481.11745449 chr6 169923959 N chr6 169924141 N DUP 18
SRR1766443.7775524 chr6 169923989 N chr6 169924065 N DEL 13
SRR1766461.1697056 chr6 169923980 N chr6 169924056 N DEL 10
SRR1766442.938096 chr6 169923967 N chr6 169924091 N DEL 10
SRR1766455.10007880 chr12 42228188 N chr12 42228315 N DUP 10
SRR1766477.2080943 chr10 2392451 N chr10 2392570 N DEL 10
SRR1766444.5589195 chr10 2392454 N chr10 2392573 N DEL 10
SRR1766485.4708893 chr10 2392458 N chr10 2392577 N DEL 10
SRR1766458.4289321 chr10 2392482 N chr10 2392730 N DEL 12
SRR1766442.37383603 chr10 2392487 N chr10 2392647 N DUP 17
SRR1766469.1566032 chr10 2392515 N chr10 2392763 N DEL 11
SRR1766458.4056319 chr10 2392488 N chr10 2392648 N DUP 12
SRR1766456.2321708 chr10 2392488 N chr10 2392605 N DUP 16
SRR1766448.229427 chr10 2392488 N chr10 2392648 N DUP 12
SRR1766483.3160667 chr10 2392482 N chr10 2392730 N DEL 16
SRR1766444.656851 chr10 2392488 N chr10 2392736 N DEL 11
SRR1766485.9920992 chr10 2392600 N chr10 2392730 N DEL 15
SRR1766466.10126575 chr10 2392600 N chr10 2392730 N DEL 15
SRR1766451.3213089 chr10 2392605 N chr10 2392774 N DEL 15
SRR1766486.1121972 chr10 60240259 N chr10 60240368 N DEL 13
SRR1766477.8986785 chr10 60240259 N chr10 60240368 N DEL 13
SRR1766451.10459403 chr10 60240271 N chr10 60240402 N DUP 13
SRR1766474.7729092 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766442.20425156 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766467.6718301 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766466.3883400 chr10 60240205 N chr10 60240303 N DEL 14
SRR1766482.7427773 chr10 60240205 N chr10 60240303 N DEL 13
SRR1766442.812296 chr17 4933971 N chr17 4934050 N DEL 13
SRR1766452.2466527 chr17 4933973 N chr17 4934052 N DEL 18
SRR1766473.11825443 chrX 72179232 N chrX 72179400 N DEL 15
SRR1766458.9586774 chr21 8464379 N chr21 8464624 N DEL 10
SRR1766442.13676881 chr21 8464564 N chr21 8464736 N DUP 18
SRR1766445.9717491 chr21 8464376 N chr21 8464882 N DEL 10
SRR1766442.24267580 chr21 8464841 N chr21 8464900 N DUP 13
SRR1766442.10665647 chr21 8464524 N chr21 8464746 N DEL 11
SRR1766458.2189670 chr21 8464762 N chr21 8464854 N DUP 10
SRR1766471.2392060 chr21 8464341 N chr21 8464796 N DEL 13
SRR1766446.4101725 chr21 8464369 N chr21 8464869 N DEL 12
SRR1766482.7714200 chr21 8464343 N chr21 8464841 N DEL 10
SRR1766442.8810644 chr21 8464343 N chr21 8464712 N DEL 12
SRR1766483.4348363 chr21 8464400 N chr21 8464876 N DEL 12
SRR1766460.8874286 chr21 8464532 N chr21 8464690 N DEL 13
SRR1766486.2980316 chr21 8464276 N chr21 8464712 N DUP 13
SRR1766467.4832535 chr21 8464789 N chr21 8464855 N DUP 10
SRR1766452.21346 chr21 8464821 N chr21 8464969 N DUP 10
SRR1766442.11262696 chr21 8464309 N chr21 8464566 N DEL 14
SRR1766464.3757429 chr21 8464532 N chr21 8464690 N DEL 13
SRR1766449.2873499 chr21 8464841 N chr21 8464894 N DUP 10
SRR1766479.12120908 chr21 8464386 N chr21 8464671 N DUP 14
SRR1766461.6805265 chr21 8464525 N chr21 8464743 N DEL 10
SRR1766480.3699048 chr21 8464841 N chr21 8464894 N DUP 10
SRR1766461.6723246 chr21 8464316 N chr21 8464581 N DEL 13
SRR1766481.12563641 chr21 8464341 N chr21 8464790 N DEL 10
SRR1766460.1772583 chr21 8464820 N chr21 8464935 N DUP 11
SRR1766485.5818323 chr21 8464742 N chr21 8465013 N DUP 10
SRR1766444.1655131 chr21 8464385 N chr21 8464919 N DUP 10
SRR1766478.11848773 chr21 8464395 N chr21 8464841 N DEL 10
SRR1766461.8239120 chr21 8464399 N chr21 8464780 N DEL 14
SRR1766457.6639652 chr21 34670028 N chr21 34670329 N DEL 11
SRR1766466.5498767 chr6 16616704 N chr6 16616761 N DEL 11
SRR1766442.14279952 chr12 5929310 N chr12 5929453 N DUP 10
SRR1766442.11314633 chr12 5929310 N chr12 5929453 N DUP 10
SRR1766459.10593179 chr12 5929310 N chr12 5929453 N DUP 11
SRR1766472.8895753 chr12 5929310 N chr12 5929453 N DUP 15
SRR1766452.3700988 chr12 5929310 N chr12 5929453 N DUP 15
SRR1766458.7161007 chr12 5929487 N chr12 5929782 N DUP 10
SRR1766464.5984668 chr12 5929501 N chr12 5929650 N DEL 10
SRR1766443.2697334 chr12 5929403 N chr12 5929550 N DUP 10
SRR1766464.1168502 chr12 5929599 N chr12 5929746 N DUP 10
SRR1766485.6063647 chr12 5929599 N chr12 5929746 N DUP 10
SRR1766465.696922 chr12 5929413 N chr12 5929782 N DUP 18
SRR1766442.42200809 chr12 5929413 N chr12 5929782 N DUP 15
SRR1766465.3969839 chr12 5929413 N chr12 5929782 N DUP 15
SRR1766484.9151315 chr12 5929635 N chr12 5929782 N DUP 10
SRR1766448.6711066 chr12 5929413 N chr12 5929782 N DUP 15
SRR1766456.3939774 chr12 5929413 N chr12 5929782 N DUP 10
SRR1766443.1801683 chr12 5929429 N chr12 5929652 N DEL 10
SRR1766476.6140423 chr12 5929630 N chr12 5929703 N DUP 10
SRR1766466.621726 chr12 5929487 N chr12 5929782 N DUP 15
SRR1766477.10533136 chr12 5929310 N chr12 5929383 N DUP 15
SRR1766449.1295593 chr12 5929348 N chr12 5929641 N DEL 10
SRR1766442.36126599 chr12 5929481 N chr12 5929704 N DEL 10
SRR1766456.2078241 chr12 5929501 N chr12 5929650 N DEL 10
SRR1766470.10141030 chr12 5929413 N chr12 5929782 N DUP 15
SRR1766482.10295176 chr12 5929413 N chr12 5929782 N DUP 10
SRR1766473.4342316 chr12 5929413 N chr12 5929782 N DUP 12
SRR1766454.2961043 chr12 5929413 N chr12 5929782 N DUP 12
SRR1766442.31065082 chr10 132980618 N chr10 132980772 N DEL 10
SRR1766461.7176706 chr10 132980758 N chr10 132980836 N DEL 10
SRR1766481.4141272 chr10 132980702 N chr10 132980909 N DUP 10
SRR1766473.10628996 chr10 132980780 N chr10 132980954 N DUP 10
SRR1766460.9222259 chr10 132980592 N chr10 132980876 N DUP 10
SRR1766464.610714 chr10 132980639 N chr10 132980870 N DEL 10
SRR1766479.10310734 chr10 132980692 N chr10 132980890 N DEL 17
SRR1766447.10545792 chr10 132980648 N chr10 132980955 N DEL 10
SRR1766473.4107834 chrX 107204842 N chrX 107205043 N DEL 12
SRR1766483.2792806 chrX 107204842 N chrX 107205043 N DEL 13
SRR1766466.9635048 chrX 107204870 N chrX 107204967 N DEL 13
SRR1766471.7817743 chrX 107204870 N chrX 107204967 N DEL 13
SRR1766462.9059923 chrX 107204827 N chrX 107204882 N DUP 19
SRR1766484.7167012 chrX 107204827 N chrX 107204882 N DUP 19
SRR1766478.11061727 chrX 107204922 N chrX 107205043 N DEL 15
SRR1766480.8300932 chrX 107204922 N chrX 107205043 N DEL 14
SRR1766470.4514772 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766464.7782581 chrX 107204898 N chrX 107205019 N DEL 13
SRR1766457.7288802 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766486.3641391 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766453.6069706 chrX 107204827 N chrX 107204906 N DUP 15
SRR1766475.5690233 chrX 107204827 N chrX 107204906 N DUP 19
SRR1766459.5660222 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766465.2885075 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766477.6988972 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766462.11206093 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766468.4946384 chrX 107204842 N chrX 107205043 N DEL 13
SRR1766447.6559092 chrX 107204846 N chrX 107205047 N DEL 11
SRR1766472.5999522 chr3 887332 N chr3 887388 N DEL 10
SRR1766476.8866578 chr3 887332 N chr3 887388 N DEL 10
SRR1766453.7127672 chr1 34102722 N chr1 34102818 N DEL 19
SRR1766477.4047385 chr1 34102728 N chr1 34102784 N DUP 15
SRR1766481.12021832 chr1 34102728 N chr1 34102784 N DUP 19
SRR1766443.1788655 chr1 34102722 N chr1 34102818 N DEL 18
SRR1766457.6683676 chr1 34102722 N chr1 34102818 N DEL 17
SRR1766464.5833726 chr1 34102722 N chr1 34102818 N DEL 17
SRR1766475.2411998 chr1 34102712 N chr1 34102827 N DEL 12
SRR1766459.10498539 chr1 34102714 N chr1 34102829 N DEL 10
SRR1766478.5525424 chr1 34102714 N chr1 34102829 N DEL 10
SRR1766458.7095308 chr8 28463387 N chr8 28463520 N DEL 10
SRR1766485.1236663 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766461.7417626 chr16 77713978 N chr16 77714221 N DUP 14
SRR1766471.5530269 chr16 77713978 N chr16 77714221 N DUP 11
SRR1766468.1127984 chr16 77713974 N chr16 77714217 N DUP 10
SRR1766470.4539864 chr16 77714034 N chr16 77714279 N DEL 10
SRR1766471.7393756 chr16 77713945 N chr16 77714249 N DUP 14
SRR1766477.10337537 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766458.7741035 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766446.7094752 chr16 77713978 N chr16 77714221 N DUP 15
SRR1766449.9990780 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766485.2350102 chr16 77714062 N chr16 77714246 N DEL 10
SRR1766442.8319229 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766442.8142213 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766465.3766743 chr16 77713977 N chr16 77714222 N DEL 10
SRR1766476.4967565 chr16 77713845 N chr16 77714225 N DEL 10
SRR1766468.3943243 chr16 77713978 N chr16 77714221 N DUP 10
SRR1766472.11653910 chr16 77714100 N chr16 77714221 N DUP 10
SRR1766442.22500358 chr16 77713978 N chr16 77714221 N DUP 10
SRR1766473.5310134 chr16 77713978 N chr16 77714221 N DUP 10
SRR1766464.9869033 chr16 77713978 N chr16 77714221 N DUP 11
SRR1766486.469049 chr16 77714218 N chr16 77714339 N DUP 10
SRR1766484.6934444 chr9 24100027 N chr9 24100088 N DUP 10
SRR1766459.141951 chr9 24100087 N chr9 24100163 N DEL 15
SRR1766464.7146132 chr3 22379398 N chr3 22379489 N DUP 10
SRR1766457.1895463 chr3 22379397 N chr3 22379472 N DUP 12
SRR1766460.4027190 chr5 1272722 N chr5 1273234 N DEL 10
SRR1766448.9611073 chr5 1272688 N chr5 1272901 N DEL 14
SRR1766482.8219950 chr5 1272688 N chr5 1273270 N DEL 14
SRR1766452.1353494 chr5 1272828 N chr5 1273883 N DEL 10
SRR1766455.188779 chr5 1273738 N chr5 1273850 N DUP 14
SRR1766462.10635448 chr5 1272759 N chr5 1273117 N DUP 10
SRR1766482.3332762 chr5 1272761 N chr5 1273673 N DUP 13
SRR1766482.11112772 chr5 1272921 N chr5 1273217 N DUP 12
SRR1766469.6686642 chr5 1272915 N chr5 1273095 N DUP 12
SRR1766482.11883006 chr5 1272880 N chr5 1273940 N DEL 10
SRR1766474.5045022 chr5 1272950 N chr5 1273940 N DEL 12
SRR1766451.4002328 chr5 1272646 N chr5 1272824 N DUP 18
SRR1766478.6070231 chr5 1272828 N chr5 1273738 N DEL 11
SRR1766448.8659739 chr5 1272705 N chr5 1273941 N DEL 14
SRR1766462.11127400 chr5 1272709 N chr5 1273945 N DEL 10
SRR1766450.6397588 chr5 1272707 N chr5 1273943 N DEL 12
SRR1766452.1028794 chr5 1272706 N chr5 1273942 N DEL 13
SRR1766442.12861091 chr7 1295473 N chr7 1295557 N DUP 12
SRR1766480.6512380 chr7 1295517 N chr7 1295603 N DUP 13
SRR1766451.1278231 chr7 1295428 N chr7 1295702 N DEL 14
SRR1766478.11455743 chr7 1295443 N chr7 1295717 N DEL 10
SRR1766452.6331120 chr7 45813283 N chr7 45813382 N DEL 10
SRR1766444.91059 chr7 45813324 N chr7 45813505 N DEL 18
SRR1766482.488163 chr7 45813249 N chr7 45813444 N DUP 11
SRR1766445.3513444 chr19 57138016 N chr19 57138178 N DUP 14
SRR1766465.6743129 chr19 57138060 N chr19 57138116 N DUP 13
SRR1766475.7586315 chr19 57137986 N chr19 57138146 N DUP 12
SRR1766469.10762129 chr19 57138052 N chr19 57138155 N DUP 10
SRR1766474.60635 chr19 57138024 N chr19 57138099 N DUP 13
SRR1766463.3412795 chr19 57138057 N chr19 57138133 N DUP 12
SRR1766442.35089032 chr19 57138028 N chr19 57138152 N DUP 12
SRR1766442.38839232 chr19 57138011 N chr19 57138242 N DUP 14
SRR1766470.9249561 chr19 57138052 N chr19 57138231 N DUP 15
SRR1766470.4003522 chr3 198168301 N chr3 198169088 N DEL 10
SRR1766482.9253841 chr3 198168416 N chr3 198168888 N DEL 10
SRR1766486.5983349 chr3 198168324 N chr3 198169046 N DUP 12
SRR1766479.7923151 chr3 198168324 N chr3 198169046 N DUP 11
SRR1766447.6382140 chr3 198168328 N chr3 198169050 N DUP 10
SRR1766473.4993679 chr3 198168364 N chr3 198168836 N DEL 15
SRR1766451.1147388 chr3 198168513 N chr3 198169396 N DEL 10
SRR1766442.2697693 chr3 198168513 N chr3 198169396 N DEL 10
SRR1766458.8507277 chr3 198168595 N chr3 198169100 N DEL 10
SRR1766470.1585656 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766462.2847133 chr3 198169225 N chr3 198169415 N DEL 10
SRR1766454.7751465 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766483.7964676 chr3 198168595 N chr3 198169415 N DEL 10
SRR1766443.3857864 chr3 198168626 N chr3 198169129 N DUP 10
SRR1766442.40805581 chr3 198168355 N chr3 198168701 N DEL 10
SRR1766464.8444301 chr3 198168292 N chr3 198168701 N DEL 10
SRR1766480.8407238 chr3 198168752 N chr3 198169129 N DUP 10
SRR1766442.34123755 chr3 198168406 N chr3 198168752 N DEL 12
SRR1766478.8185470 chr3 198168752 N chr3 198168940 N DUP 10
SRR1766484.9415166 chr3 198168752 N chr3 198168940 N DUP 10
SRR1766448.1998186 chr3 198168802 N chr3 198169307 N DEL 10
SRR1766482.5096010 chr3 198168773 N chr3 198169150 N DUP 15
SRR1766442.25227893 chr3 198168773 N chr3 198169150 N DUP 15
SRR1766442.18645038 chr3 198168773 N chr3 198169150 N DUP 13
SRR1766445.4493860 chr3 198168773 N chr3 198169150 N DUP 11
SRR1766442.23240159 chr3 198168688 N chr3 198169319 N DEL 15
SRR1766486.5983349 chr3 198168420 N chr3 198168829 N DEL 10
SRR1766454.1401927 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766471.1101035 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766442.8618175 chr3 198168428 N chr3 198168837 N DEL 10
SRR1766465.4324141 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766444.6857119 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766455.6253367 chr3 198168428 N chr3 198168837 N DEL 10
SRR1766480.6787953 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766467.9442482 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766464.832250 chr3 198168591 N chr3 198169535 N DUP 10
SRR1766442.34604789 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766477.7101214 chr3 198168815 N chr3 198169066 N DUP 10
SRR1766446.4642990 chr3 198168595 N chr3 198168848 N DEL 10
SRR1766485.776469 chr3 198168355 N chr3 198168827 N DEL 10
SRR1766471.2064196 chr3 198168353 N chr3 198168825 N DEL 10
SRR1766462.1723348 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766463.7625470 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766482.3827695 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766473.1681528 chr3 198168848 N chr3 198168910 N DUP 10
SRR1766477.1343927 chr3 198168299 N chr3 198169525 N DUP 10
SRR1766485.12100895 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766459.1218682 chr3 198168888 N chr3 198169139 N DUP 10
SRR1766484.4162833 chr3 198168794 N chr3 198169047 N DEL 10
SRR1766472.2526073 chr3 198168762 N chr3 198168950 N DUP 10
SRR1766482.9253841 chr3 198168636 N chr3 198168950 N DUP 10
SRR1766452.6384526 chr3 198168762 N chr3 198168950 N DUP 10
SRR1766453.10082429 chr3 198168338 N chr3 198169186 N DUP 15
SRR1766442.31879319 chr3 198168825 N chr3 198168950 N DUP 10
SRR1766454.6879471 chr3 198168513 N chr3 198168953 N DUP 10
SRR1766447.9921110 chr3 198168427 N chr3 198168836 N DEL 10
SRR1766462.4508420 chr3 198168580 N chr3 198168959 N DEL 10
SRR1766470.9600531 chr3 198168972 N chr3 198169288 N DEL 10
SRR1766451.1147388 chr3 198168580 N chr3 198168959 N DEL 10
SRR1766452.1424623 chr3 198169224 N chr3 198169288 N DEL 10
SRR1766457.503391 chr3 198168428 N chr3 198168837 N DEL 10
SRR1766448.2303111 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766474.2192381 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766478.11096723 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766475.4682199 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766473.4683580 chr3 198169048 N chr3 198169362 N DUP 10
SRR1766468.2547939 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766486.7845216 chr3 198169047 N chr3 198169361 N DUP 10
SRR1766449.3403725 chr3 198169369 N chr3 198169433 N DEL 10
SRR1766473.9311745 chr3 198169055 N chr3 198169117 N DUP 10
SRR1766442.16936494 chr3 198168794 N chr3 198169047 N DEL 10
SRR1766458.8507277 chr3 198168676 N chr3 198169055 N DEL 10
SRR1766446.2005536 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766442.37051932 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766462.8845260 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766459.7820729 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766478.8149081 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766448.10141482 chr3 198168762 N chr3 198168950 N DUP 10
SRR1766443.3217929 chr3 198168394 N chr3 198169055 N DEL 10
SRR1766442.5783748 chr3 198168762 N chr3 198168950 N DUP 10
SRR1766443.7510034 chr3 198168457 N chr3 198169055 N DEL 10
SRR1766467.4594022 chr3 198168395 N chr3 198169056 N DEL 10
SRR1766460.4744481 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766446.9440374 chr3 198169098 N chr3 198169288 N DEL 10
SRR1766450.6116059 chr3 198169098 N chr3 198169288 N DEL 10
SRR1766465.10534219 chr3 198169098 N chr3 198169288 N DEL 10
SRR1766460.4744481 chr3 198168843 N chr3 198168905 N DUP 10
SRR1766460.9798777 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766444.6298511 chr3 198168825 N chr3 198168950 N DUP 10
SRR1766484.2970205 chr3 198168825 N chr3 198168950 N DUP 10
SRR1766479.13019236 chr3 198168825 N chr3 198168950 N DUP 10
SRR1766453.6561226 chr3 198168958 N chr3 198169148 N DEL 10
SRR1766451.5885465 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766442.13409660 chr3 198168420 N chr3 198169396 N DEL 10
SRR1766453.10136296 chr3 198168418 N chr3 198168638 N DEL 10
SRR1766470.6730709 chr3 198168613 N chr3 198169055 N DEL 10
SRR1766484.9748975 chr3 198168357 N chr3 198169396 N DEL 10
SRR1766447.10449885 chr3 198168420 N chr3 198169396 N DEL 10
SRR1766466.2801333 chr3 198168416 N chr3 198168825 N DEL 10
SRR1766442.28744001 chr3 198169181 N chr3 198169495 N DUP 10
SRR1766442.27572363 chr3 198168418 N chr3 198168638 N DEL 10
SRR1766446.8068417 chr3 198169047 N chr3 198169172 N DUP 10
SRR1766445.2284530 chr3 198168866 N chr3 198169180 N DUP 15
SRR1766471.747624 chr3 198169047 N chr3 198169172 N DUP 10
SRR1766473.7100442 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766479.6955620 chr3 198169047 N chr3 198169172 N DUP 10
SRR1766486.1130915 chr3 198169047 N chr3 198169172 N DUP 10
SRR1766451.5914311 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766472.2095336 chr3 198169180 N chr3 198169433 N DEL 15
SRR1766447.9827794 chr3 198168497 N chr3 198169252 N DUP 10
SRR1766465.671698 chr3 198169369 N chr3 198169433 N DEL 13
SRR1766466.2502959 chr3 198168513 N chr3 198169205 N DUP 10
SRR1766481.10912235 chr3 198169036 N chr3 198169226 N DEL 10
SRR1766454.5089271 chr3 198168549 N chr3 198169243 N DEL 10
SRR1766478.8688477 chr3 198168549 N chr3 198169243 N DEL 10
SRR1766479.3581095 chr3 198168909 N chr3 198169288 N DEL 12
SRR1766465.1965398 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766452.2248917 chr3 198168909 N chr3 198169288 N DEL 15
SRR1766459.4870445 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766476.8882488 chr3 198168928 N chr3 198169307 N DEL 15
SRR1766477.9288504 chr3 198168802 N chr3 198169307 N DEL 15
SRR1766460.8661718 chr3 198168676 N chr3 198169307 N DEL 15
SRR1766450.252618 chr3 198169140 N chr3 198169328 N DUP 10
SRR1766442.23240159 chr3 198168394 N chr3 198169307 N DEL 10
SRR1766446.10204673 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766459.4870445 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766460.5977806 chr3 198169224 N chr3 198169288 N DEL 14
SRR1766443.1207970 chr3 198169047 N chr3 198169361 N DUP 10
SRR1766447.3271600 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766449.9644855 chr3 198169047 N chr3 198169361 N DUP 10
SRR1766448.391205 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766453.1085413 chr3 198169224 N chr3 198169288 N DEL 15
SRR1766474.2192381 chr3 198169224 N chr3 198169288 N DEL 15
SRR1766442.38264626 chr3 198169224 N chr3 198169288 N DEL 15
SRR1766452.1424623 chr3 198169224 N chr3 198169288 N DEL 13
SRR1766442.12012906 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766465.10534219 chr3 198169369 N chr3 198169433 N DEL 10
SRR1766479.10326344 chr3 198169180 N chr3 198169433 N DEL 15
SRR1766461.2947535 chr3 198169369 N chr3 198169433 N DEL 10
SRR1766459.1759401 chr3 198168626 N chr3 198169192 N DUP 12
SRR1766459.10902306 chr3 198169140 N chr3 198169202 N DUP 10
SRR1766464.5484446 chr3 198168889 N chr3 198169394 N DEL 10
SRR1766475.1988528 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766452.10032623 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766452.10032623 chr3 198169224 N chr3 198169288 N DEL 12
SRR1766477.10850804 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766442.33436551 chr3 198169224 N chr3 198169288 N DEL 15
SRR1766486.1810069 chr3 198169224 N chr3 198169288 N DEL 13
SRR1766445.54561 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766447.1649448 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766461.2947535 chr3 198169224 N chr3 198169288 N DEL 10
SRR1766456.3346227 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766469.7577147 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766472.10629820 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766452.4383822 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766467.9003657 chr3 198169080 N chr3 198169396 N DEL 10
SRR1766463.1766669 chr3 198168823 N chr3 198169389 N DUP 10
SRR1766442.22820724 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766464.7279379 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766451.9781443 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766451.6884696 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766452.1509551 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766470.5199415 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766479.3818572 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766443.7224086 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766469.8352623 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766473.2918984 chr3 198168294 N chr3 198169396 N DEL 11
SRR1766473.6114207 chr3 198168297 N chr3 198169399 N DEL 11
SRR1766442.34082399 chr3 198168295 N chr3 198169397 N DEL 14
SRR1766454.6331897 chr3 198168295 N chr3 198169397 N DEL 14
SRR1766480.4875857 chr3 198168513 N chr3 198168890 N DUP 10
SRR1766460.9485661 chr3 198168676 N chr3 198169055 N DEL 10
SRR1766450.3205339 chr3 198169180 N chr3 198169433 N DEL 13
SRR1766452.9769942 chr3 198169369 N chr3 198169433 N DEL 10
SRR1766473.6968027 chr3 198168898 N chr3 198168962 N DEL 10
SRR1766481.7178966 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766447.433975 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766474.8529549 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766461.6468289 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766467.10458266 chr3 198168866 N chr3 198169369 N DUP 10
SRR1766452.2023421 chr3 198169307 N chr3 198169495 N DUP 10
SRR1766484.2144915 chr12 129388110 N chr12 129388275 N DUP 10
SRR1766482.2166763 chr19 47802706 N chr19 47802815 N DEL 12
SRR1766452.1172948 chr11 59632741 N chr11 59632802 N DUP 10
SRR1766472.11009848 chr11 59632741 N chr11 59632802 N DUP 11
SRR1766442.31034937 chr11 59632741 N chr11 59632802 N DUP 11
SRR1766479.2848175 chr11 59632741 N chr11 59632802 N DUP 11
SRR1766454.7510045 chr11 59632758 N chr11 59632896 N DUP 11
SRR1766453.10320305 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766450.7426073 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766464.8162357 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766449.2984884 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766475.10377551 chr11 59632745 N chr11 59632905 N DUP 10
SRR1766472.11075332 chr11 59632758 N chr11 59632896 N DUP 17
SRR1766447.891614 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766451.1611213 chr11 59632758 N chr11 59632896 N DUP 11
SRR1766476.6201423 chr11 59632758 N chr11 59632896 N DUP 14
SRR1766465.8666844 chr11 59632758 N chr11 59632896 N DUP 14
SRR1766479.5032663 chr11 59632755 N chr11 59632897 N DEL 15
SRR1766459.7519141 chr14 91044491 N chr14 91044542 N DEL 17
SRR1766484.11474737 chr1 81747030 N chr1 81747113 N DEL 14
SRR1766475.8965645 chr14 104325061 N chr14 104325190 N DUP 10
SRR1766477.1099365 chr14 104325126 N chr14 104325191 N DUP 14
SRR1766449.5620478 chr14 104325139 N chr14 104325266 N DUP 10
SRR1766466.8296672 chr14 104325139 N chr14 104325266 N DUP 10
SRR1766442.8660600 chr14 104325139 N chr14 104325266 N DUP 10
SRR1766479.12956037 chr14 104325140 N chr14 104325267 N DUP 10
SRR1766442.9005132 chr21 14261871 N chr21 14261948 N DUP 13
SRR1766443.5580810 chr21 14261873 N chr21 14261950 N DUP 13
SRR1766446.1585090 chr21 14261873 N chr21 14261950 N DUP 13
SRR1766449.1360291 chr21 14261871 N chr21 14261948 N DUP 13
SRR1766474.8544762 chr21 14261874 N chr21 14261951 N DUP 12
SRR1766460.18178 chr21 14261872 N chr21 14261949 N DUP 14
SRR1766452.6758425 chr21 14261871 N chr21 14261948 N DUP 17
SRR1766485.11016921 chr21 14261871 N chr21 14261948 N DUP 18
SRR1766442.41054206 chr4 4220180 N chr4 4220245 N DUP 14
SRR1766462.10518422 chrX 649100 N chrX 649153 N DEL 10
SRR1766446.10003 chrX 649094 N chrX 649167 N DUP 11
SRR1766481.7302533 chrX 649071 N chrX 649196 N DEL 11
SRR1766448.10642261 chr2 30263892 N chr2 30264211 N DEL 10
SRR1766485.10433661 chr21 45501821 N chr21 45501951 N DEL 10
SRR1766449.2761965 chr21 45501821 N chr21 45501951 N DEL 10
SRR1766475.1586005 chr21 45501821 N chr21 45501951 N DEL 10
SRR1766462.5933631 chr21 45501821 N chr21 45501951 N DEL 10
SRR1766449.10881995 chr21 45501840 N chr21 45502097 N DUP 10
SRR1766470.3741626 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766469.4529495 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766468.5392343 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766465.5211463 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766481.187727 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766442.35278987 chr21 45501808 N chr21 45502022 N DUP 14
SRR1766471.11294967 chr21 45501850 N chr21 45502023 N DEL 10
SRR1766475.10758435 chr21 45501850 N chr21 45502023 N DEL 10
SRR1766449.1431250 chr21 45501850 N chr21 45502023 N DEL 10
SRR1766465.2663227 chr21 45501849 N chr21 45502109 N DEL 13
SRR1766477.4743806 chr21 45501849 N chr21 45502109 N DEL 15
SRR1766448.1960208 chr21 45501914 N chr21 45502218 N DEL 16
SRR1766474.4879850 chr21 45501871 N chr21 45502218 N DEL 15
SRR1766442.44674105 chr21 45502108 N chr21 45502239 N DEL 15
SRR1766469.6628223 chr21 45502112 N chr21 45502243 N DEL 11
SRR1766470.912384 chr6 34683567 N chr6 34683648 N DUP 11
SRR1766473.688089 chr6 34683567 N chr6 34683648 N DUP 11
SRR1766442.8348651 chr6 34683567 N chr6 34683648 N DUP 13
SRR1766464.10567720 chr20 35539681 N chr20 35539732 N DEL 12
SRR1766463.9499511 chr20 35539681 N chr20 35539732 N DEL 12
SRR1766459.5517392 chr1 11522690 N chr1 11522911 N DEL 11
SRR1766448.4861640 chr1 11522690 N chr1 11522911 N DEL 18
SRR1766445.6787493 chr1 11522701 N chr1 11522790 N DEL 18
SRR1766469.6336979 chr1 11522911 N chr1 11522976 N DUP 15
SRR1766460.10284557 chr1 11522777 N chr1 11522866 N DEL 16
SRR1766448.2677992 chr1 11522766 N chr1 11523020 N DEL 18
SRR1766468.3122618 chr1 11522771 N chr1 11522836 N DUP 16
SRR1766476.3342138 chr1 11522723 N chr1 11522779 N DEL 16
SRR1766481.6948997 chr1 11522800 N chr1 11522856 N DEL 15
SRR1766474.2416296 chr1 11522778 N chr1 11522865 N DUP 15
SRR1766467.2864822 chr1 11522757 N chr1 11522855 N DUP 14
SRR1766442.47184389 chr1 11522705 N chr1 11522761 N DEL 10
SRR1766482.7986008 chr1 11522811 N chr1 11522964 N DUP 13
SRR1766455.766176 chr1 11522855 N chr1 11522999 N DEL 15
SRR1766462.1403498 chr1 11522722 N chr1 11522778 N DEL 12
SRR1766460.10284557 chr1 11522856 N chr1 11523020 N DUP 11
SRR1766477.3418572 chr1 11522801 N chr1 11522899 N DUP 11
SRR1766447.1021930 chr1 11522847 N chr1 11522901 N DUP 15
SRR1766482.3461498 chr1 11522833 N chr1 11522898 N DUP 15
SRR1766449.10815081 chr1 11522867 N chr1 11522954 N DUP 15
SRR1766474.2416296 chr1 11522724 N chr1 11522877 N DUP 14
SRR1766444.5884168 chr1 11522844 N chr1 11522911 N DEL 15
SRR1766459.11097738 chr1 11522837 N chr1 11522968 N DUP 10
SRR1766447.10571861 chr1 11522790 N chr1 11522912 N DEL 13
SRR1766477.3418572 chr1 11522834 N chr1 11522965 N DUP 10
SRR1766457.759551 chr1 11522834 N chr1 11522899 N DUP 15
SRR1766465.4579191 chr1 11522790 N chr1 11523064 N DUP 10
SRR1766444.1242946 chr1 11522889 N chr1 11522987 N DUP 10
SRR1766458.3373386 chr1 11522779 N chr1 11522921 N DUP 15
SRR1766462.9391873 chr1 11522887 N chr1 11522943 N DEL 17
SRR1766467.2534300 chr1 11522833 N chr1 11522898 N DUP 10
SRR1766447.966989 chr1 11522795 N chr1 11522871 N DUP 19
SRR1766445.2206400 chr1 11522756 N chr1 11522953 N DUP 16
SRR1766447.3775181 chr1 11522833 N chr1 11522898 N DUP 14
SRR1766458.8995500 chr1 11522682 N chr1 11522978 N DUP 11
SRR1766477.8399597 chr1 11522782 N chr1 11522990 N DUP 15
SRR1766472.2718692 chr1 11522728 N chr1 11522839 N DEL 11
SRR1766458.598827 chr1 11522834 N chr1 11522910 N DUP 10
SRR1766472.11932065 chr1 11522689 N chr1 11522888 N DEL 10
SRR1766457.1623244 chr1 11522933 N chr1 11522987 N DUP 10
SRR1766482.10486760 chr1 11522800 N chr1 11522900 N DEL 10
SRR1766471.7637015 chr1 11522673 N chr1 11522892 N DUP 15
SRR1766484.5106505 chr1 11522899 N chr1 11522999 N DEL 14
SRR1766471.2626925 chr1 11522876 N chr1 11522943 N DEL 10
SRR1766464.906067 chr1 11522683 N chr1 11522946 N DUP 16
SRR1766480.4017982 chr1 11522867 N chr1 11522954 N DUP 15
SRR1766484.5106505 chr1 11522713 N chr1 11522822 N DUP 15
SRR1766463.9240650 chr1 11522893 N chr1 11523004 N DEL 10
SRR1766460.1744327 chr1 11522746 N chr1 11522833 N DUP 10
SRR1766467.4875381 chr1 11522733 N chr1 11523029 N DUP 11
SRR1766442.32466797 chr1 11522943 N chr1 11523063 N DUP 10
SRR1766469.550113 chr1 11522909 N chr1 11522998 N DEL 12
SRR1766483.11554571 chr1 11522866 N chr1 11523087 N DEL 10
SRR1766442.36692428 chr1 11522807 N chr1 11523072 N DEL 10
SRR1766477.1710911 chr1 11522866 N chr1 11523087 N DEL 15
SRR1766446.6835560 chr1 11522877 N chr1 11523087 N DEL 15
SRR1766470.3235227 chr1 11522717 N chr1 11523103 N DEL 18
SRR1766479.4367259 chr1 11522888 N chr1 11523087 N DEL 17
SRR1766462.1512512 chr4 6512078 N chr4 6512181 N DEL 10
SRR1766464.1845413 chr4 6512032 N chr4 6512685 N DUP 17
SRR1766462.7118319 chr4 6511969 N chr4 6512046 N DUP 10
SRR1766451.4246617 chr4 6511751 N chr4 6512788 N DUP 15
SRR1766442.37250888 chr4 6511696 N chr4 6511964 N DEL 10
SRR1766442.32331045 chr4 6512514 N chr4 6512803 N DEL 17
SRR1766464.6617698 chr4 6512005 N chr4 6512174 N DEL 15
SRR1766443.946713 chr4 6511751 N chr4 6512059 N DUP 19
SRR1766480.44355 chr4 6511672 N chr4 6512157 N DUP 15
SRR1766463.9707609 chr4 6512061 N chr4 6512587 N DEL 15
SRR1766479.4778171 chr4 6511987 N chr4 6512391 N DUP 12
SRR1766462.1998124 chr4 6512040 N chr4 6512404 N DEL 16
SRR1766479.9659673 chr4 6512511 N chr4 6512803 N DEL 11
SRR1766482.7953450 chr4 6511565 N chr4 6512146 N DUP 15
SRR1766481.9635619 chr4 6512072 N chr4 6512595 N DEL 10
SRR1766486.4322751 chr4 6512011 N chr4 6512085 N DUP 11
SRR1766459.2358773 chr4 6511803 N chr4 6511909 N DEL 15
SRR1766449.9487334 chr4 6511719 N chr4 6512686 N DEL 15
SRR1766443.6249558 chr4 6511900 N chr4 6511967 N DEL 19
SRR1766480.1557525 chr4 6512001 N chr4 6512092 N DEL 10
SRR1766449.9019694 chr4 6512042 N chr4 6512166 N DEL 10
SRR1766476.884049 chr4 6511783 N chr4 6512681 N DEL 16
SRR1766474.11273852 chr4 6511751 N chr4 6512038 N DUP 18
SRR1766478.7571584 chr4 6512036 N chr4 6512310 N DEL 15
SRR1766479.13279782 chr4 6511684 N chr4 6512076 N DUP 15
SRR1766467.6755552 chr4 6512267 N chr4 6512625 N DEL 16
SRR1766483.11286513 chr4 6512436 N chr4 6512674 N DEL 17
SRR1766477.8968558 chr4 6511751 N chr4 6512068 N DUP 19
SRR1766484.3012884 chr4 6511688 N chr4 6512838 N DEL 10
SRR1766474.7706815 chr4 6511699 N chr4 6512073 N DUP 10
SRR1766442.46992958 chr4 6512445 N chr4 6512641 N DEL 18
SRR1766462.5307146 chr4 6512041 N chr4 6512390 N DEL 15
SRR1766467.2766808 chr4 6512334 N chr4 6512803 N DEL 17
SRR1766471.729973 chr4 6511727 N chr4 6512022 N DUP 11
SRR1766472.643150 chr4 6512238 N chr4 6512803 N DEL 17
SRR1766460.3690639 chr4 6511522 N chr4 6511655 N DEL 12
SRR1766481.5943877 chr4 6512014 N chr4 6512670 N DUP 12
SRR1766454.4584699 chr4 6511774 N chr4 6512067 N DUP 18
SRR1766442.18117396 chr4 6511963 N chr4 6512553 N DUP 17
SRR1766474.3663873 chr4 6511977 N chr4 6512075 N DUP 17
SRR1766484.1532911 chr4 6512238 N chr4 6512803 N DEL 17
SRR1766452.6525913 chr4 6512122 N chr4 6512642 N DEL 17
SRR1766458.6656436 chr4 6512064 N chr4 6512662 N DEL 15
SRR1766469.10460161 chr4 6512008 N chr4 6512079 N DUP 10
SRR1766442.15562102 chr4 6511800 N chr4 6512159 N DUP 14
SRR1766483.11340352 chr4 6512511 N chr4 6512803 N DEL 11
SRR1766478.5148229 chr4 6512029 N chr4 6512115 N DUP 17
SRR1766446.10068454 chr4 6511672 N chr4 6512064 N DUP 15
SRR1766449.10862705 chr4 6511522 N chr4 6511691 N DEL 10
SRR1766442.22326896 chr4 6511933 N chr4 6511983 N DUP 11
SRR1766466.4087488 chr4 6511541 N chr4 6512235 N DEL 16
SRR1766472.6267779 chr4 6512004 N chr4 6512326 N DEL 12
SRR1766444.2734046 chr4 6511722 N chr4 6512662 N DEL 10
SRR1766476.7290640 chr4 6512078 N chr4 6512628 N DEL 10
SRR1766474.3016922 chr4 6511761 N chr4 6512075 N DUP 11
SRR1766452.5242026 chr4 6512511 N chr4 6512803 N DEL 11
SRR1766454.1913741 chr4 6511756 N chr4 6512076 N DUP 18
SRR1766452.6525913 chr4 6512054 N chr4 6512475 N DEL 15
SRR1766442.25782208 chr11 134738880 N chr11 134739013 N DEL 19
SRR1766442.44233628 chr11 134738880 N chr11 134739013 N DEL 14
SRR1766481.8157875 chr11 134738883 N chr11 134739106 N DUP 10
SRR1766486.875628 chr11 134738867 N chr11 134739060 N DEL 15
SRR1766478.10230582 chr18 76896488 N chr18 76896537 N DUP 10
SRR1766451.9729379 chr4 2856748 N chr4 2857073 N DEL 10
SRR1766478.2437952 chr4 2856812 N chr4 2857134 N DEL 12
SRR1766479.4303626 chr4 2856796 N chr4 2857118 N DEL 10
SRR1766467.4065500 chrX 142126033 N chrX 142126097 N DEL 10
SRR1766469.5630912 chrX 142126115 N chrX 142126198 N DEL 12
SRR1766459.7612526 chrX 142126115 N chrX 142126198 N DEL 12
SRR1766476.6471060 chrX 142126133 N chrX 142126203 N DEL 11
SRR1766463.5107930 chrX 142126133 N chrX 142126203 N DEL 14
SRR1766452.7510255 chrX 142126133 N chrX 142126203 N DEL 15
SRR1766471.2454953 chr21 42591832 N chr21 42591903 N DEL 10
SRR1766449.330591 chr18 41349899 N chr18 41349967 N DUP 13
SRR1766451.4955734 chr18 41349886 N chr18 41349996 N DUP 12
SRR1766448.8984370 chr18 41349886 N chr18 41349996 N DUP 13
SRR1766451.6414193 chr18 41349886 N chr18 41349996 N DUP 14
SRR1766460.3994208 chr18 41349886 N chr18 41349996 N DUP 16
SRR1766485.4573420 chr18 41349886 N chr18 41349996 N DUP 16
SRR1766453.2523118 chr18 41349926 N chr18 41350003 N DUP 18
SRR1766485.12036142 chr5 173129190 N chr5 173129527 N DEL 10
SRR1766445.895049 chr9 40590175 N chr9 40590342 N DEL 13
SRR1766475.9732305 chr6 94711526 N chr6 94711888 N DUP 14
SRR1766442.30049145 chr6 94711526 N chr6 94711888 N DUP 14
SRR1766442.26998185 chr6 94711670 N chr6 94711854 N DUP 10
SRR1766454.8228689 chr6 94711525 N chr6 94711761 N DEL 11
SRR1766475.9732305 chr6 94711511 N chr6 94711888 N DUP 14
SRR1766466.9728593 chr5 162906168 N chr5 162906219 N DEL 14
SRR1766472.140325 chr10 73262122 N chr10 73262217 N DUP 12
SRR1766478.1726151 chr10 73262122 N chr10 73262217 N DUP 12
SRR1766484.9450932 chr10 73262122 N chr10 73262217 N DUP 12
SRR1766449.984472 chr10 73262172 N chr10 73262231 N DEL 10
SRR1766470.723184 chr9 69340774 N chr9 69340841 N DEL 10
SRR1766473.7764161 chr9 69340761 N chr9 69340856 N DEL 12
SRR1766475.2695665 chr9 69340785 N chr9 69340934 N DEL 10
SRR1766477.4935965 chr9 69340830 N chr9 69340951 N DEL 11
SRR1766480.8708878 chr9 69340818 N chr9 69340885 N DEL 16
SRR1766484.5103234 chr9 69340817 N chr9 69340886 N DUP 10
SRR1766445.6515273 chr9 69340897 N chr9 69340976 N DUP 10
SRR1766458.7064041 chr9 69340860 N chr9 69340913 N DEL 17
SRR1766476.10594913 chr9 69340870 N chr9 69340939 N DEL 19
SRR1766482.2451125 chr9 69340870 N chr9 69340939 N DEL 15
SRR1766463.9860548 chr9 69340774 N chr9 69340965 N DEL 12
SRR1766471.4633476 chr18 72675687 N chr18 72675778 N DEL 15
SRR1766481.11282398 chr18 72675797 N chr18 72675888 N DEL 10
SRR1766479.2750750 chr18 72675816 N chr18 72675907 N DEL 15
SRR1766479.3512450 chr18 72675811 N chr18 72675902 N DEL 10
SRR1766451.3483997 chr2 168631704 N chr2 168631765 N DUP 10
SRR1766457.4946375 chr2 168631704 N chr2 168631765 N DUP 11
SRR1766461.5970728 chr21 40498824 N chr21 40498885 N DEL 11
SRR1766484.6832801 chr21 40498824 N chr21 40498885 N DEL 17
SRR1766480.589887 chr21 40498824 N chr21 40498885 N DEL 13
SRR1766459.7914985 chr21 40498824 N chr21 40498885 N DEL 13
SRR1766471.9171108 chr21 40498824 N chr21 40498885 N DEL 16
SRR1766452.9452455 chr21 40498824 N chr21 40498885 N DEL 16
SRR1766460.8572665 chr21 40498864 N chr21 40498955 N DEL 10
SRR1766451.8221494 chr21 40498828 N chr21 40498889 N DEL 11
SRR1766462.3425978 chr21 40498864 N chr21 40498955 N DEL 15
SRR1766460.3089862 chr21 40498869 N chr21 40498960 N DEL 10
SRR1766447.1562684 chr12 121750661 N chr12 121751045 N DEL 11
SRR1766469.2479386 chr12 121750803 N chr12 121751030 N DEL 12
SRR1766463.6787856 chr12 121751023 N chr12 121751493 N DEL 11
SRR1766468.1780920 chr12 121750947 N chr12 121751177 N DEL 12
SRR1766480.7317745 chr12 121751272 N chr12 121751513 N DUP 11
SRR1766448.1816541 chr17 8829691 N chr17 8829742 N DUP 17
SRR1766471.5853055 chr17 8829514 N chr17 8829751 N DEL 15
SRR1766471.4697917 chr11 89112662 N chr11 89112823 N DEL 11
SRR1766479.7530684 chr6 168257712 N chr6 168257801 N DEL 10
SRR1766445.5859122 chr6 168257676 N chr6 168257745 N DEL 13
SRR1766462.3731772 chr20 64017391 N chr20 64017788 N DEL 16
SRR1766444.2643093 chr20 64017416 N chr20 64017769 N DEL 11
SRR1766465.3457480 chr22 49477091 N chr22 49477256 N DEL 10
SRR1766481.10478203 chr22 49477091 N chr22 49477948 N DEL 15
SRR1766467.7030489 chr22 49477091 N chr22 49477313 N DEL 12
SRR1766465.3457480 chr22 49477012 N chr22 49477325 N DEL 11
SRR1766448.10595125 chr22 49477081 N chr22 49477333 N DEL 10
SRR1766485.5525528 chr22 49477528 N chr22 49477623 N DEL 10
SRR1766467.2267873 chr22 49477610 N chr22 49477766 N DEL 14
SRR1766466.5081350 chr22 49476992 N chr22 49477661 N DUP 14
SRR1766462.11123785 chr22 49477070 N chr22 49477868 N DUP 10
SRR1766457.3349760 chr22 49477354 N chr22 49477892 N DUP 10
SRR1766481.12591158 chr22 49477502 N chr22 49477953 N DEL 11
SRR1766467.6876468 chr22 49477092 N chr22 49477979 N DEL 11
SRR1766460.8446611 chr18 9887642 N chr18 9887823 N DEL 17
SRR1766442.21531532 chr18 9887525 N chr18 9887749 N DUP 14
SRR1766456.3273218 chr18 9887604 N chr18 9887695 N DEL 10
SRR1766448.8387519 chr6 157283053 N chr6 157283466 N DUP 10
SRR1766486.1596459 chr1 228631234 N chr1 228631293 N DUP 12
SRR1766444.4096235 chr2 118305297 N chr2 118305361 N DEL 12
SRR1766465.11120104 chr2 118305296 N chr2 118305358 N DUP 10
SRR1766461.5992344 chr2 118305297 N chr2 118305361 N DEL 19
SRR1766448.6374881 chr2 118305687 N chr2 118305766 N DUP 15
SRR1766464.10849360 chr2 118305687 N chr2 118305766 N DUP 15
SRR1766445.2480899 chr2 118305687 N chr2 118305766 N DUP 15
SRR1766485.7484538 chr16 48932387 N chr16 48932500 N DUP 16
SRR1766455.3653124 chr2 105210478 N chr2 105211118 N DEL 10
SRR1766481.7362363 chr18 79237007 N chr18 79237117 N DEL 10
SRR1766464.1524448 chr18 79236956 N chr18 79237117 N DEL 10
SRR1766471.4802654 chr18 79236902 N chr18 79237061 N DUP 10
SRR1766474.2101939 chr18 79237069 N chr18 79237499 N DEL 10
SRR1766470.9526081 chr3 127154843 N chr3 127155086 N DEL 11
SRR1766446.7547004 chr1 232368459 N chr1 232368722 N DUP 15
SRR1766442.26787874 chr19 53990572 N chr19 53990683 N DEL 13
SRR1766442.39206125 chr19 53991199 N chr19 53991271 N DUP 11
SRR1766454.2721593 chr19 53990751 N chr19 53991263 N DEL 17
SRR1766448.9487496 chr19 53990753 N chr19 53991265 N DEL 17
SRR1766455.4415555 chr19 53990716 N chr19 53991265 N DEL 17
SRR1766466.1766866 chr19 53990713 N chr19 53991262 N DEL 13
SRR1766474.6535639 chr19 53990713 N chr19 53991262 N DEL 10
SRR1766445.2330495 chr19 53990713 N chr19 53991262 N DEL 10
SRR1766461.6559010 chr19 53990677 N chr19 53991263 N DEL 10
SRR1766481.4076187 chr19 53990677 N chr19 53991263 N DEL 10
SRR1766442.11489316 chrX 23523383 N chrX 23523497 N DEL 15
SRR1766465.10783745 chr4 168793335 N chr4 168793434 N DEL 11
SRR1766483.11265334 chr4 168793311 N chr4 168793410 N DEL 12
SRR1766472.232346 chr4 168793359 N chr4 168793458 N DEL 11
SRR1766474.2549351 chr4 168793311 N chr4 168793410 N DEL 11
SRR1766459.9212335 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766481.2024056 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766455.1325294 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766442.8588090 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766467.11788071 chr4 168793418 N chr4 168793516 N DEL 11
SRR1766444.833047 chr4 168793418 N chr4 168793516 N DEL 11
SRR1766463.8305745 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766459.9267253 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766459.9982881 chr4 168793284 N chr4 168793532 N DUP 10
SRR1766445.2189057 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766443.2235559 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766479.2134224 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766486.82444 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766453.8348741 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766481.3212651 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766443.904725 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766466.881151 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766447.598630 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766460.10706412 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766442.19349917 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766443.6213861 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766471.2318564 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766458.2755623 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766449.9613880 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766477.399156 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766454.4999230 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766479.13870801 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766458.2553896 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766450.189355 chr4 168793322 N chr4 168793516 N DEL 11
SRR1766453.6179082 chr4 168793323 N chr4 168793517 N DEL 16
SRR1766479.9068621 chr4 168793322 N chr4 168793516 N DEL 11
SRR1766456.2709829 chr4 168793322 N chr4 168793516 N DEL 11
SRR1766449.5797437 chr4 168793322 N chr4 168793516 N DEL 11
SRR1766442.32762427 chr4 168793298 N chr4 168793516 N DEL 11
SRR1766460.3374870 chr4 168793298 N chr4 168793516 N DEL 11
SRR1766452.3058440 chr4 168793298 N chr4 168793516 N DEL 11
SRR1766479.5943555 chr4 168793298 N chr4 168793516 N DEL 11
SRR1766476.868937 chr7 158950530 N chr7 158950836 N DEL 10
SRR1766453.2591929 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766473.144859 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766444.6055709 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766475.6087177 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766459.9278196 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766442.29821866 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766478.9747975 chr7 158950737 N chr7 158950919 N DUP 10
SRR1766467.4728417 chr7 158950920 N chr7 158951041 N DUP 10
SRR1766462.7581550 chr17 82009748 N chr17 82009920 N DEL 11
SRR1766457.1322557 chr17 82009753 N chr17 82009807 N DUP 10
SRR1766459.8869696 chr19 54770329 N chr19 54770465 N DEL 10
SRR1766469.8213701 chr19 54770300 N chr19 54770608 N DUP 11
SRR1766479.10274469 chr19 54770331 N chr19 54770563 N DEL 14
SRR1766466.8709599 chr19 54770459 N chr19 54770691 N DEL 15
SRR1766450.9543883 chr17 44984425 N chr17 44985186 N DUP 13
SRR1766478.2121904 chr17 44984590 N chr17 44985327 N DUP 14
SRR1766480.7793587 chr17 44984600 N chr17 44985229 N DUP 10
SRR1766469.2935742 chr17 44984707 N chr17 44985140 N DEL 15
SRR1766463.7427346 chr17 44984359 N chr17 44984630 N DEL 11
SRR1766447.7352218 chr17 44984749 N chr17 44985270 N DUP 16
SRR1766482.4546937 chr17 44984644 N chr17 44985156 N DUP 10
SRR1766466.2394144 chr17 44984909 N chr17 44985268 N DUP 10
SRR1766457.914526 chr17 44984774 N chr17 44985178 N DUP 10
SRR1766450.5937451 chr17 44984585 N chr17 44985178 N DUP 11
SRR1766442.10596442 chr17 44984692 N chr17 44985242 N DEL 13
SRR1766478.6794463 chr17 44984680 N chr17 44985284 N DEL 10
SRR1766464.8921506 chr17 44984653 N chr17 44985257 N DEL 18
SRR1766477.3929566 chr17 44985184 N chr17 44985302 N DEL 10
SRR1766464.6843622 chrY 10646342 N chrY 10646672 N DEL 10
SRR1766465.9847987 chr10 102637416 N chr10 102637532 N DUP 12
SRR1766442.1763377 chr10 102637718 N chr10 102637807 N DUP 11
SRR1766464.960101 chr10 102637701 N chr10 102637823 N DUP 14
SRR1766442.33601028 chr10 102637739 N chr10 102637833 N DUP 16
SRR1766472.4239913 chr10 102637740 N chr10 102637797 N DUP 14
SRR1766465.7725181 chr10 102637718 N chr10 102637807 N DUP 11
SRR1766459.7466408 chr10 102637739 N chr10 102637833 N DUP 19
SRR1766445.3651237 chrX 35600911 N chrX 35601011 N DUP 14
SRR1766450.4639613 chrX 35600886 N chrX 35601030 N DUP 10
SRR1766470.5548123 chrX 35600889 N chrX 35601037 N DUP 14
SRR1766473.714143 chrX 35600898 N chrX 35601070 N DUP 14
SRR1766458.1716387 chrX 35600936 N chrX 35601011 N DUP 17
SRR1766465.2637436 chrX 35600939 N chrX 35601007 N DUP 12
SRR1766480.1051086 chrX 35600939 N chrX 35601007 N DUP 11
SRR1766442.17847578 chrX 35600949 N chrX 35601017 N DUP 19
SRR1766452.10449664 chrX 35600972 N chrX 35601077 N DUP 18
SRR1766442.11179291 chrX 35600897 N chrX 35601030 N DUP 10
SRR1766459.4268173 chrX 35600887 N chrX 35601054 N DUP 13
SRR1766442.30999057 chrX 35600949 N chrX 35601006 N DUP 16
SRR1766484.415740 chrX 35600949 N chrX 35601006 N DUP 16
SRR1766451.4261790 chrX 35600981 N chrX 35601095 N DUP 17
SRR1766469.8810954 chrX 35600974 N chrX 35601135 N DUP 10
SRR1766446.1977179 chrX 35600927 N chrX 35600986 N DUP 11
SRR1766446.3687907 chrX 35600927 N chrX 35600986 N DUP 11
SRR1766473.9910788 chrX 35600914 N chrX 35600969 N DUP 17
SRR1766474.7604554 chrX 35600949 N chrX 35601010 N DUP 16
SRR1766462.4034393 chrX 35600925 N chrX 35601009 N DUP 11
SRR1766457.4979407 chrX 35600873 N chrX 35600944 N DEL 13
SRR1766452.2239816 chrX 35600789 N chrX 35600928 N DEL 16
SRR1766449.8215278 chrX 35600913 N chrX 35601041 N DUP 10
SRR1766442.36879467 chrX 35600888 N chrX 35601021 N DUP 19
SRR1766463.4124714 chrX 35600919 N chrX 35601063 N DUP 12
SRR1766475.8228710 chrX 35600919 N chrX 35601063 N DUP 18
SRR1766485.3403172 chrX 35600919 N chrX 35601063 N DUP 19
SRR1766474.6117537 chrX 35600765 N chrX 35601085 N DUP 15
SRR1766465.1754152 chr16 17167628 N chr16 17167753 N DEL 10
SRR1766483.1193136 chr16 17167662 N chr16 17167725 N DEL 10
SRR1766465.8383353 chr16 17167662 N chr16 17167725 N DEL 10
SRR1766455.9858731 chr16 17167562 N chr16 17167685 N DUP 15
SRR1766446.2438935 chr16 17167662 N chr16 17167725 N DEL 10
SRR1766455.9858804 chr16 17167562 N chr16 17167716 N DUP 10
SRR1766479.6327442 chr16 17167753 N chr16 17167814 N DUP 10
SRR1766458.9053629 chr16 17167628 N chr16 17167753 N DEL 13
SRR1766444.3103207 chr16 17167799 N chr16 17167862 N DEL 15
SRR1766472.3250424 chr16 17167843 N chr16 17167999 N DEL 19
SRR1766455.779315 chr16 17167613 N chr16 17167862 N DEL 10
SRR1766472.7347093 chr7 105433769 N chr7 105433905 N DEL 19
SRR1766445.1717709 chr11 101629020 N chr11 101629084 N DUP 19
SRR1766480.118460 chr5 43136640 N chr5 43136801 N DEL 11
SRR1766448.8068102 chr11 71362100 N chr11 71362485 N DEL 13
SRR1766442.17665723 chr11 71362165 N chr11 71363037 N DEL 15
SRR1766473.5157919 chr11 71362222 N chr11 71362671 N DEL 14
SRR1766447.5894118 chr11 71362257 N chr11 71362658 N DEL 16
SRR1766449.4645274 chr11 71362227 N chr11 71362939 N DEL 10
SRR1766465.11210800 chr11 71362307 N chr11 71362995 N DEL 15
SRR1766466.5005942 chr11 71362305 N chr11 71362658 N DEL 10
SRR1766471.9152596 chr11 71362311 N chr11 71362408 N DEL 14
SRR1766464.7570945 chr11 71362327 N chr11 71362807 N DEL 13
SRR1766449.2647419 chr11 71362461 N chr11 71363356 N DEL 11
SRR1766470.3575750 chr11 71362509 N chr11 71362965 N DEL 15
SRR1766460.1980267 chr11 71362515 N chr11 71362851 N DEL 14
SRR1766460.5861818 chr11 71362497 N chr11 71363321 N DEL 18
SRR1766472.10784921 chr11 71362464 N chr11 71362886 N DUP 11
SRR1766445.727329 chr11 71362549 N chr11 71362662 N DEL 10
SRR1766449.5479671 chr11 71362472 N chr11 71362870 N DUP 13
SRR1766456.4229224 chr11 71362543 N chr11 71362823 N DEL 15
SRR1766467.7172944 chr11 71362569 N chr11 71362658 N DEL 15
SRR1766446.5774531 chr11 71362569 N chr11 71362658 N DEL 16
SRR1766464.9570163 chr11 71362513 N chr11 71362991 N DUP 15
SRR1766485.5978334 chr11 71362190 N chr11 71362597 N DUP 10
SRR1766442.33072783 chr11 71362583 N chr11 71363167 N DEL 14
SRR1766469.2613072 chr11 71362214 N chr11 71362511 N DEL 15
SRR1766468.5177052 chr11 71362524 N chr11 71362834 N DUP 15
SRR1766465.5169907 chr11 71362591 N chr11 71362871 N DEL 12
SRR1766478.4976335 chr11 71362342 N chr11 71362511 N DEL 10
SRR1766445.8402921 chr11 71362529 N chr11 71362903 N DUP 12
SRR1766466.2328616 chr11 71362524 N chr11 71362834 N DUP 15
SRR1766460.7385137 chr11 71362605 N chr11 71362965 N DEL 10
SRR1766481.5419689 chr11 71362205 N chr11 71362550 N DEL 10
SRR1766485.9379500 chr11 71362560 N chr11 71362695 N DUP 10
SRR1766450.9315424 chr11 71362685 N chr11 71363356 N DEL 15
SRR1766479.12672498 chr11 71362236 N chr11 71362613 N DEL 17
SRR1766442.12162768 chr11 71362365 N chr11 71362700 N DUP 15
SRR1766478.3558518 chr11 71362679 N chr11 71363159 N DEL 15
SRR1766472.5416717 chr11 71362636 N chr11 71362890 N DUP 15
SRR1766449.6633775 chr11 71362636 N chr11 71362890 N DUP 15
SRR1766473.5110401 chr11 71362326 N chr11 71362639 N DEL 10
SRR1766474.4577651 chr11 71362641 N chr11 71363079 N DUP 10
SRR1766486.917352 chr11 71362652 N chr11 71362986 N DUP 10
SRR1766484.4953417 chr11 71362214 N chr11 71362655 N DEL 10
SRR1766485.9033971 chr11 71362658 N chr11 71362824 N DUP 10
SRR1766447.11179387 chr11 71362587 N chr11 71362779 N DEL 10
SRR1766481.5258286 chr11 71362868 N chr11 71363157 N DEL 13
SRR1766482.6952144 chr11 71362559 N chr11 71362861 N DUP 10
SRR1766446.4475112 chr11 71362619 N chr11 71362787 N DEL 10
SRR1766466.6559651 chr11 71362897 N chr11 71363186 N DEL 13
SRR1766473.1464989 chr11 71362894 N chr11 71363175 N DEL 15
SRR1766453.2445991 chr11 71362659 N chr11 71362897 N DUP 10
SRR1766461.8189875 chr11 71362205 N chr11 71362813 N DEL 13
SRR1766452.7927641 chr11 71362213 N chr11 71362813 N DEL 15
SRR1766457.2138614 chr11 71362813 N chr11 71362988 N DUP 11
SRR1766470.1359243 chr11 71362855 N chr11 71363166 N DUP 10
SRR1766484.8698302 chr11 71362863 N chr11 71363206 N DUP 15
SRR1766446.3196653 chr11 71362184 N chr11 71362990 N DUP 11
SRR1766456.1307408 chr11 71362901 N chr11 71363188 N DUP 15
SRR1766477.10958934 chr11 71362918 N chr11 71363181 N DUP 11
SRR1766465.11210800 chr11 71362207 N chr11 71362927 N DEL 15
SRR1766467.5595986 chr11 71362426 N chr11 71362938 N DEL 10
SRR1766471.2296894 chr11 71362674 N chr11 71362938 N DEL 10
SRR1766442.4336325 chr11 71362215 N chr11 71362959 N DEL 10
SRR1766448.9344259 chr11 71362965 N chr11 71363188 N DUP 12
SRR1766442.29131103 chr11 71363010 N chr11 71363081 N DUP 10
SRR1766448.2289497 chr11 71363031 N chr11 71363110 N DUP 17
SRR1766455.8415563 chr11 71363010 N chr11 71363081 N DUP 10
SRR1766475.4023532 chr11 71362842 N chr11 71362995 N DEL 11
SRR1766453.7954749 chr11 71362698 N chr11 71363010 N DEL 15
SRR1766459.916242 chr11 71363010 N chr11 71363345 N DUP 10
SRR1766442.27533844 chr11 71362213 N chr11 71363013 N DEL 10
SRR1766452.10412259 chr11 71363118 N chr11 71363374 N DEL 11
SRR1766445.3357383 chr11 71363067 N chr11 71363385 N DUP 15
SRR1766475.4358429 chr11 71362664 N chr11 71363142 N DUP 15
SRR1766484.3690769 chr11 71363151 N chr11 71363296 N DEL 15
SRR1766480.3540835 chr11 71363166 N chr11 71363436 N DUP 18
SRR1766445.7582500 chr11 71363097 N chr11 71363154 N DEL 10
SRR1766485.1435462 chr11 71362185 N chr11 71363183 N DUP 12
SRR1766471.10629522 chr11 71362988 N chr11 71363149 N DEL 16
SRR1766471.7148702 chr11 71362986 N chr11 71363163 N DEL 18
SRR1766478.3655375 chr11 71362938 N chr11 71363209 N DUP 12
SRR1766473.3677126 chr11 71363095 N chr11 71363152 N DEL 10
SRR1766444.1552354 chr11 71362843 N chr11 71363148 N DEL 10
SRR1766470.6829964 chr11 71362204 N chr11 71363164 N DEL 10
SRR1766446.7945186 chr11 71362988 N chr11 71363157 N DEL 16
SRR1766467.2515553 chr11 71363159 N chr11 71363278 N DUP 12
SRR1766447.1172997 chr11 71362893 N chr11 71363222 N DEL 10
SRR1766466.6559651 chr11 71363261 N chr11 71363427 N DUP 15
SRR1766467.1238712 chr11 71362382 N chr11 71363222 N DEL 10
SRR1766478.3558518 chr11 71362690 N chr11 71363250 N DEL 12
SRR1766450.8030381 chr11 71363185 N chr11 71363282 N DEL 12
SRR1766484.11211100 chr11 71363203 N chr11 71363284 N DEL 10
SRR1766455.8453985 chr11 71362215 N chr11 71363295 N DEL 10
SRR1766443.8525842 chr11 71363086 N chr11 71363366 N DEL 17
SRR1766445.3103884 chr19 55530597 N chr19 55530934 N DEL 11
SRR1766443.10812473 chr6 95502056 N chr6 95502163 N DUP 18
SRR1766473.6699064 chr6 95502056 N chr6 95502163 N DUP 19
SRR1766442.21787624 chr6 95502075 N chr6 95502146 N DUP 18
SRR1766463.1810392 chr6 95502102 N chr6 95502247 N DEL 12
SRR1766469.10892917 chr6 95502060 N chr6 95502332 N DUP 16
SRR1766452.3848279 chr6 95502225 N chr6 95502310 N DUP 18
SRR1766465.812864 chr6 95502326 N chr6 95502414 N DEL 16
SRR1766443.9439229 chr6 95502263 N chr6 95502324 N DUP 17
SRR1766445.325905 chr6 95502263 N chr6 95502324 N DUP 17
SRR1766455.9427814 chr6 95502522 N chr6 95503045 N DEL 15
SRR1766450.10426355 chr6 95502562 N chr6 95503099 N DEL 14
SRR1766450.98598 chr6 95502562 N chr6 95503099 N DEL 14
SRR1766451.8225970 chr6 95502531 N chr6 95503132 N DEL 10
SRR1766483.8520803 chr6 95502603 N chr6 95503268 N DUP 11
SRR1766474.3642564 chr6 95502603 N chr6 95503268 N DUP 10
SRR1766443.4658238 chr6 95502532 N chr6 95503205 N DEL 11
SRR1766478.5601427 chr6 95502533 N chr6 95503243 N DEL 10
SRR1766452.1068694 chr1 109654236 N chr1 109654340 N DEL 10
SRR1766464.9546549 chr1 109654236 N chr1 109654340 N DEL 10
SRR1766481.1909562 chr1 109654236 N chr1 109654340 N DEL 10
SRR1766467.2741961 chr1 109654236 N chr1 109654340 N DEL 18
SRR1766462.1217967 chr3 9639315 N chr3 9639364 N DUP 13
SRR1766476.6111175 chr7 60919991 N chr7 60920137 N DUP 10
SRR1766468.4353498 chr7 60919976 N chr7 60920122 N DUP 10
SRR1766455.9808171 chr7 60919991 N chr7 60920137 N DUP 15
SRR1766448.2413914 chr15 63547907 N chr15 63548006 N DUP 11
SRR1766468.3452328 chr15 63547953 N chr15 63548038 N DEL 15
SRR1766475.6928772 chr15 63547953 N chr15 63548038 N DEL 15
SRR1766461.1328256 chr15 63547956 N chr15 63548041 N DEL 12
SRR1766470.7748660 chr1 24907789 N chr1 24907863 N DUP 12
SRR1766462.9549874 chr1 24907853 N chr1 24907904 N DEL 19
SRR1766449.25683 chr1 24907798 N chr1 24907847 N DUP 15
SRR1766461.6646043 chr1 24907814 N chr1 24907888 N DUP 10
SRR1766448.4688978 chr1 24907883 N chr1 24908259 N DEL 15
SRR1766476.4593966 chr1 24907958 N chr1 24908384 N DEL 17
SRR1766463.9151774 chr1 24907839 N chr1 24908013 N DUP 10
SRR1766471.10855959 chr1 24908063 N chr1 24908139 N DEL 10
SRR1766461.1487471 chr1 24907797 N chr1 24908071 N DUP 15
SRR1766464.5546754 chr1 24908123 N chr1 24908224 N DEL 10
SRR1766442.45998972 chr1 24908113 N chr1 24908214 N DEL 12
SRR1766479.9220674 chr1 24908123 N chr1 24908172 N DUP 11
SRR1766449.10873285 chr1 24907958 N chr1 24908184 N DEL 15
SRR1766442.29140521 chr1 24907783 N chr1 24908184 N DEL 15
SRR1766456.2379281 chr1 24908214 N chr1 24908263 N DUP 10
SRR1766442.28055915 chr1 24908214 N chr1 24908263 N DUP 15
SRR1766477.5304532 chr1 24908214 N chr1 24908263 N DUP 15
SRR1766452.9406567 chr1 24908214 N chr1 24908263 N DUP 10
SRR1766485.3604234 chr1 24908282 N chr1 24908333 N DEL 10
SRR1766447.6754007 chr1 24908199 N chr1 24908273 N DUP 10
SRR1766464.7141671 chr1 24908214 N chr1 24908263 N DUP 14
SRR1766469.4339725 chr1 24908251 N chr1 24908327 N DEL 15
SRR1766475.2712178 chr1 24908282 N chr1 24908333 N DEL 15
SRR1766477.6135919 chr1 24908208 N chr1 24908284 N DEL 10
SRR1766484.1858938 chr1 24908208 N chr1 24908284 N DEL 10
SRR1766442.24885332 chr1 24908282 N chr1 24908333 N DEL 11
SRR1766479.13071233 chr1 24908273 N chr1 24908349 N DEL 10
SRR1766457.5759551 chr1 24907808 N chr1 24908359 N DEL 10
SRR1766477.1740154 chr1 24907864 N chr1 24908440 N DEL 10
SRR1766460.10188705 chr1 24908241 N chr1 24908442 N DEL 10
SRR1766445.9655537 chr7 205405 N chr7 205496 N DUP 14
SRR1766451.5194082 chr1 125179352 N chr1 125179428 N DEL 12
SRR1766442.33367673 chr1 125179358 N chr1 125179434 N DEL 10
SRR1766469.2496600 chr17 44590386 N chr17 44591083 N DEL 10
SRR1766464.9138537 chr17 44590415 N chr17 44590930 N DEL 10
SRR1766454.1684115 chr17 44590385 N chr17 44590606 N DUP 15
SRR1766483.10037354 chr17 44590677 N chr17 44591092 N DEL 10
SRR1766445.3499027 chr17 44590620 N chr17 44591127 N DUP 14
SRR1766442.15969032 chr17 44590395 N chr17 44590740 N DUP 12
SRR1766443.8243244 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766473.2822904 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766484.3240924 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766475.9173113 chr17 44590740 N chr17 44591091 N DEL 13
SRR1766463.6044678 chr17 44590740 N chr17 44591091 N DEL 13
SRR1766449.7492892 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766471.6130177 chr17 44590761 N chr17 44590930 N DEL 18
SRR1766442.10353299 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766450.8761951 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766477.2407161 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766479.13315133 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766455.947410 chr17 44590389 N chr17 44590734 N DUP 11
SRR1766478.11726904 chr17 44590422 N chr17 44590765 N DEL 13
SRR1766471.213104 chr17 44590270 N chr17 44591057 N DEL 10
SRR1766450.1105841 chr16 88470628 N chr16 88470679 N DEL 10
SRR1766479.11691689 chr2 3171190 N chr2 3171244 N DUP 18
SRR1766460.3353206 chr2 3170821 N chr2 3171216 N DEL 10
SRR1766481.9609543 chr11 134759990 N chr11 134760197 N DUP 15
SRR1766443.5917413 chr11 134760031 N chr11 134760104 N DUP 18
SRR1766456.3078444 chr11 134760031 N chr11 134760104 N DUP 15
SRR1766466.4152538 chr11 134760031 N chr11 134760104 N DUP 14
SRR1766483.3873771 chr11 134760031 N chr11 134760104 N DUP 10
SRR1766485.517087 chr11 134760040 N chr11 134760395 N DUP 10
SRR1766442.7435638 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766482.6260456 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766474.9422298 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766457.7477206 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766443.35058 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766443.10428085 chr11 134760094 N chr11 134760301 N DUP 16
SRR1766462.1531734 chr11 134760143 N chr11 134760202 N DUP 11
SRR1766446.9018027 chr11 134760211 N chr11 134760286 N DEL 15
SRR1766447.10436602 chr11 134760143 N chr11 134760202 N DUP 11
SRR1766442.10088735 chr11 134760143 N chr11 134760202 N DUP 18
SRR1766475.6873438 chr11 134760144 N chr11 134760351 N DUP 10
SRR1766456.3047089 chr11 134760004 N chr11 134760285 N DUP 14
SRR1766468.7882697 chr11 134760104 N chr11 134760239 N DEL 10
SRR1766462.5882867 chr11 134760063 N chr11 134760344 N DUP 10
SRR1766445.8997835 chr1 241713498 N chr1 241713566 N DEL 14
SRR1766481.2768284 chr1 22227678 N chr1 22227733 N DUP 16
SRR1766469.9191209 chr22 18418066 N chr22 18418235 N DEL 13
SRR1766466.9481213 chr22 18418066 N chr22 18418235 N DEL 15
SRR1766450.1178376 chr22 18418212 N chr22 18418294 N DUP 17
SRR1766465.4943142 chr22 18418212 N chr22 18418294 N DUP 18
SRR1766485.10781574 chr22 18418212 N chr22 18418294 N DUP 19
SRR1766477.3328323 chr22 18418212 N chr22 18418294 N DUP 17
SRR1766465.5426755 chr22 18418189 N chr22 18418266 N DUP 15
SRR1766449.8824936 chr22 18418145 N chr22 18418209 N DEL 14
SRR1766459.10890299 chr22 18418060 N chr22 18418211 N DEL 10
SRR1766459.9571510 chr22 18418143 N chr22 18418391 N DUP 10
SRR1766442.22207367 chr22 18418140 N chr22 18418410 N DEL 19
SRR1766476.5808589 chr22 18418140 N chr22 18418410 N DEL 19
SRR1766457.4857609 chr22 18418144 N chr22 18418416 N DEL 10
SRR1766442.11542737 chr22 18418547 N chr22 18418729 N DUP 11
SRR1766478.10964601 chr22 18418547 N chr22 18418729 N DUP 14
SRR1766442.31499190 chr1 225833808 N chr1 225834419 N DEL 12
SRR1766479.295951 chr18 59233868 N chr18 59233988 N DEL 12
SRR1766483.3881660 chr18 59233868 N chr18 59233988 N DEL 12
SRR1766478.8731711 chr18 59233835 N chr18 59233932 N DUP 11
SRR1766475.9609132 chr18 59233810 N chr18 59233931 N DUP 15
SRR1766446.3165791 chr18 59233835 N chr18 59233932 N DUP 13
SRR1766466.3317853 chr18 59233852 N chr18 59233901 N DUP 14
SRR1766442.9341603 chr18 59233751 N chr18 59234005 N DUP 14
SRR1766461.10760957 chr18 59233823 N chr18 59234088 N DUP 12
SRR1766458.5704118 chr18 59234185 N chr18 59234258 N DEL 11
SRR1766448.6989772 chr18 59234185 N chr18 59234258 N DEL 13
SRR1766469.7383809 chr18 59234187 N chr18 59234260 N DEL 10
SRR1766481.1496601 chr18 59234187 N chr18 59234260 N DEL 10
SRR1766470.7982521 chrX 140768792 N chrX 140768849 N DEL 12
SRR1766481.10174862 chrX 140768792 N chrX 140768849 N DEL 13
SRR1766442.20578156 chr12 5928554 N chr12 5928618 N DEL 13
SRR1766442.20617090 chr12 5928554 N chr12 5928618 N DEL 13
SRR1766442.25710574 chr12 5928554 N chr12 5928618 N DEL 13
SRR1766452.7158607 chr12 5928554 N chr12 5928618 N DEL 18
SRR1766468.5479529 chr12 5928691 N chr12 5929724 N DEL 10
SRR1766461.10704418 chr12 5928691 N chr12 5929724 N DEL 15
SRR1766470.6906476 chr12 5928691 N chr12 5929724 N DEL 15
SRR1766442.35696168 chr12 5928691 N chr12 5929724 N DEL 15
SRR1766467.1280076 chr12 5928691 N chr12 5929724 N DEL 15
SRR1766446.3027580 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766459.2811676 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766477.9709290 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766449.9216613 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766471.12207763 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766452.6820522 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766469.4702599 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766446.7427157 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766459.898553 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766446.10526081 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766459.3715909 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766477.10938337 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766469.3814881 chr12 5929797 N chr12 5929868 N DEL 10
SRR1766475.4266602 chr12 5929797 N chr12 5929868 N DEL 10
SRR1766482.550243 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766454.5418474 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766475.5056492 chr12 5928663 N chr12 5928810 N DUP 10
SRR1766482.3930703 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766442.34141561 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766443.6187103 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766453.1126053 chr12 5928744 N chr12 5929263 N DEL 10
SRR1766470.6387460 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766486.11566260 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766467.8152235 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766470.3645154 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766470.3952904 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766456.2132819 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766458.2751128 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766477.4216808 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766478.1657900 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766464.8127649 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766477.4271506 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766484.809816 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766442.13385760 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766449.907380 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766442.16581484 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766475.961206 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766442.40349687 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766469.10298811 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766458.2911336 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766460.8653614 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766482.3930703 chr12 5928894 N chr12 5929337 N DUP 10
SRR1766456.2132819 chr12 5929511 N chr12 5929804 N DEL 15
SRR1766462.8068802 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766447.6487537 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766450.8794248 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766465.2393348 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766481.424250 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766481.6765539 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766471.3674475 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766481.7697176 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766484.9151315 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766474.7186199 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766442.13385760 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766455.9250164 chr12 5928894 N chr12 5929337 N DUP 10
SRR1766463.3562469 chr12 5929804 N chr12 5929877 N DUP 10
SRR1766459.4505908 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766473.3316822 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766446.6596242 chr12 5928894 N chr12 5929337 N DUP 10
SRR1766482.6561632 chr12 5928663 N chr12 5928958 N DUP 10
SRR1766463.2108008 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766442.13764130 chr12 5928892 N chr12 5929629 N DEL 10
SRR1766442.41978246 chr12 5929269 N chr12 5929782 N DUP 10
SRR1766454.5418474 chr12 5928744 N chr12 5929263 N DEL 10
SRR1766478.2533654 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766483.3214319 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766442.26905964 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766459.4629066 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766456.3939774 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766475.5056492 chr12 5929424 N chr12 5930087 N DEL 14
SRR1766473.529077 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766475.9371722 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766456.4130722 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766457.8425680 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766459.4629066 chr12 5929789 N chr12 5930082 N DEL 10
SRR1766471.7865627 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766477.4899102 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766454.4674653 chr12 5928681 N chr12 5929274 N DEL 10
SRR1766469.1265258 chr12 5929367 N chr12 5929804 N DEL 13
SRR1766442.14279952 chr12 5929422 N chr12 5930085 N DEL 10
SRR1766442.11314633 chr12 5929422 N chr12 5930085 N DEL 10
SRR1766459.10593179 chr12 5929422 N chr12 5930085 N DEL 11
SRR1766472.8895753 chr12 5929419 N chr12 5930082 N DEL 15
SRR1766452.3700988 chr12 5929422 N chr12 5930085 N DEL 15
SRR1766448.8597871 chr12 5928760 N chr12 5930085 N DEL 10
SRR1766458.7161007 chr12 5929487 N chr12 5929782 N DUP 10
SRR1766442.6809372 chr12 5928905 N chr12 5929492 N DUP 10
SRR1766477.2409670 chr12 5928905 N chr12 5929492 N DUP 10
SRR1766464.5984668 chr12 5929493 N chr12 5930082 N DEL 10
SRR1766447.8588736 chr12 5929511 N chr12 5929804 N DEL 11
SRR1766443.2697334 chr12 5929511 N chr12 5929804 N DEL 15
SRR1766478.2533654 chr12 5928744 N chr12 5929263 N DEL 10
SRR1766442.23668787 chr12 5929650 N chr12 5929867 N DUP 10
SRR1766465.696922 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766442.42200809 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766465.3969839 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766448.6711066 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766456.3939774 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766443.1801683 chr12 5929429 N chr12 5929652 N DEL 10
SRR1766466.621726 chr12 5929491 N chr12 5929786 N DUP 10
SRR1766448.6711066 chr12 5929337 N chr12 5929848 N DEL 10
SRR1766442.36126599 chr12 5928978 N chr12 5929715 N DEL 15
SRR1766456.2078241 chr12 5928905 N chr12 5929492 N DUP 10
SRR1766482.612998 chr12 5928663 N chr12 5930282 N DUP 10
SRR1766469.2484114 chr12 5928978 N chr12 5929715 N DEL 11
SRR1766448.10418503 chr12 5928756 N chr12 5929715 N DEL 10
SRR1766470.10141030 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766481.11343330 chr12 5928756 N chr12 5929715 N DEL 10
SRR1766442.46155632 chr12 5928756 N chr12 5929715 N DEL 10
SRR1766482.10295176 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766442.29850140 chr12 5928756 N chr12 5929715 N DEL 10
SRR1766473.4342316 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766454.2961043 chr12 5929642 N chr12 5930081 N DUP 10
SRR1766465.696922 chr12 5928687 N chr12 5929792 N DUP 13
SRR1766446.9972609 chr12 5928687 N chr12 5929792 N DUP 13
SRR1766479.10974705 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766474.2704687 chr12 5928687 N chr12 5929792 N DUP 14
SRR1766486.2490837 chr12 5929346 N chr12 5929804 N DEL 13
SRR1766453.7185109 chr12 5929346 N chr12 5929804 N DEL 13
SRR1766462.2937861 chr12 5928703 N chr12 5929806 N DEL 13
SRR1766442.32418744 chr12 5928927 N chr12 5929808 N DEL 10
SRR1766478.3802562 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766466.7490940 chr12 5929354 N chr12 5929865 N DEL 10
SRR1766472.7826794 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766455.408025 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766444.4841162 chr12 5929789 N chr12 5930082 N DEL 12
SRR1766463.1949630 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766469.9544908 chr12 5928668 N chr12 5928741 N DUP 10
SRR1766443.6694150 chr12 5929645 N chr12 5929792 N DUP 10
SRR1766465.9789340 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766485.11783333 chr12 5929932 N chr12 5930007 N DEL 10
SRR1766442.30731671 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766443.9452570 chr12 5928684 N chr12 5930009 N DEL 10
SRR1766473.4342316 chr12 5929337 N chr12 5929848 N DEL 10
SRR1766474.10714393 chr12 5928894 N chr12 5929337 N DUP 10
SRR1766478.5441170 chr12 5929525 N chr12 5929746 N DUP 10
SRR1766481.4209435 chr12 5929501 N chr12 5929650 N DEL 10
SRR1766466.1999136 chr12 5929777 N chr12 5930292 N DEL 10
SRR1766466.5373344 chr12 5929777 N chr12 5930292 N DEL 12
SRR1766485.6063647 chr12 5928686 N chr12 5930011 N DEL 10
SRR1766464.4366081 chr12 5929511 N chr12 5929804 N DEL 10
SRR1766442.17094521 chr12 5929511 N chr12 5929804 N DEL 10
SRR1766463.4931578 chr12 5928894 N chr12 5929777 N DUP 10
SRR1766442.30731671 chr12 5929548 N chr12 5929915 N DEL 10
SRR1766442.1774884 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766482.9718139 chr12 5928903 N chr12 5929786 N DUP 10
SRR1766442.14279952 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766444.4841162 chr12 5929269 N chr12 5929782 N DUP 10
SRR1766465.9789340 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766459.5087434 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766479.10974705 chr12 5929269 N chr12 5929782 N DUP 10
SRR1766454.6337178 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766486.2490837 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766464.1168502 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766465.3724642 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766470.2808913 chr12 5930143 N chr12 5930292 N DEL 15
SRR1766446.9972609 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766474.9457543 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766455.5300617 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766455.5652074 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766460.700694 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766456.998954 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766469.9006952 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766453.7185109 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766452.10252382 chr12 5929777 N chr12 5930292 N DEL 11
SRR1766469.1101461 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766477.7193919 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766482.9184375 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766460.2497917 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766467.4086271 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766474.3521928 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766474.2550569 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766465.3807061 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766474.11667806 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766462.3698742 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766460.10344977 chr12 5929341 N chr12 5930296 N DEL 10
SRR1766482.11871869 chr3 186874222 N chr3 186874348 N DUP 12
SRR1766483.7398782 chr3 186874415 N chr3 186874494 N DEL 18
SRR1766452.3029510 chr3 186874415 N chr3 186874494 N DEL 15
SRR1766468.84702 chr19 458138 N chr19 458244 N DEL 10
SRR1766447.1320653 chr19 458137 N chr19 458687 N DEL 13
SRR1766458.1639952 chr19 458758 N chr19 458907 N DEL 10
SRR1766466.7941485 chr19 458294 N chr19 458697 N DEL 10
SRR1766470.8196713 chr7 63204972 N chr7 63205169 N DEL 14
SRR1766477.3574256 chr15 71564790 N chr15 71564844 N DEL 10
SRR1766450.7543360 chr15 71564790 N chr15 71564844 N DEL 11
SRR1766449.6751310 chr15 71564790 N chr15 71564844 N DEL 12
SRR1766480.7910161 chr2 239101994 N chr2 239102247 N DEL 10
SRR1766456.654239 chr19 10187807 N chr19 10188081 N DEL 10
SRR1766466.4287147 chr21 44953585 N chr21 44953635 N DUP 17
SRR1766463.8860220 chr21 44953585 N chr21 44953635 N DUP 17
SRR1766442.29204173 chr21 44953585 N chr21 44953635 N DUP 19
SRR1766465.6000768 chr8 28882646 N chr8 28882702 N DUP 14
SRR1766485.7409267 chr8 28882640 N chr8 28882696 N DUP 14
SRR1766442.31660393 chr8 28882644 N chr8 28882696 N DUP 15
SRR1766486.11178811 chr12 122093068 N chr12 122093269 N DUP 10
SRR1766463.8847399 chr12 122093069 N chr12 122093270 N DUP 10
SRR1766452.1592492 chr16 13019916 N chr16 13020021 N DUP 15
SRR1766460.2282043 chr16 13019916 N chr16 13020021 N DUP 15
SRR1766484.3780150 chr16 6773320 N chr16 6773422 N DUP 13
SRR1766457.4703329 chr16 6773320 N chr16 6773424 N DUP 15
SRR1766452.9864072 chr21 5329582 N chr21 5329646 N DUP 14
SRR1766449.7799874 chr21 5329580 N chr21 5329812 N DUP 10
SRR1766453.6875770 chr21 5329767 N chr21 5329841 N DUP 15
SRR1766462.2752522 chr11 473723 N chr11 473858 N DUP 19
SRR1766442.16078834 chr11 473726 N chr11 473861 N DUP 12
SRR1766462.1490056 chr11 473788 N chr11 473855 N DUP 12
SRR1766452.4597343 chr9 9275208 N chr9 9275278 N DEL 10
SRR1766462.8462440 chr9 9275257 N chr9 9275359 N DEL 13
SRR1766446.8531159 chr9 9275243 N chr9 9275349 N DEL 18
SRR1766482.5720344 chr9 9275243 N chr9 9275349 N DEL 18
SRR1766461.5205440 chr1 228633475 N chr1 228633534 N DUP 12
SRR1766454.7963000 chr1 228633477 N chr1 228633530 N DUP 11
SRR1766456.5628066 chr1 163552239 N chr1 163552396 N DEL 15
SRR1766462.7106137 chr1 163552239 N chr1 163552357 N DEL 10
SRR1766442.44251767 chr2 90382996 N chr2 90383045 N DUP 10
SRR1766470.6503296 chr2 90382998 N chr2 90383096 N DUP 10
SRR1766480.2428879 chr10 83462788 N chr10 83462919 N DUP 15
SRR1766452.447774 chr10 83462829 N chr10 83462919 N DUP 12
SRR1766447.11314208 chr10 83462899 N chr10 83462964 N DUP 10
SRR1766457.8216012 chr10 83462899 N chr10 83462964 N DUP 10
SRR1766470.1476081 chr1 3176212 N chr1 3176430 N DUP 15
SRR1766474.10155820 chr1 3176110 N chr1 3176307 N DEL 10
SRR1766455.3959176 chr1 3176302 N chr1 3176428 N DUP 11
SRR1766479.12487080 chr1 3176306 N chr1 3176440 N DUP 15
SRR1766470.3357621 chr8 70935280 N chr8 70935363 N DEL 10
SRR1766473.7952460 chr8 70935279 N chr8 70935362 N DEL 11
SRR1766482.9816880 chr8 70935282 N chr8 70935363 N DEL 10
SRR1766442.7384271 chr6 54310807 N chr6 54310873 N DEL 18
SRR1766471.10140423 chr6 54310807 N chr6 54310873 N DEL 16
SRR1766462.6687958 chr6 54310796 N chr6 54311048 N DUP 10
SRR1766482.2157800 chrX 131138107 N chrX 131138174 N DEL 12
SRR1766476.8579295 chr3 98837019 N chr3 98837182 N DUP 13
SRR1766462.794707 chr3 98836932 N chr3 98837207 N DUP 10
SRR1766480.675749 chr3 98837064 N chr3 98837191 N DUP 11
SRR1766474.10223131 chr3 98836936 N chr3 98837211 N DUP 15
SRR1766458.7059989 chr3 98836967 N chr3 98837242 N DUP 10
SRR1766450.4800700 chr11 90155473 N chr11 90155553 N DEL 11
SRR1766451.2844129 chr2 231848993 N chr2 231849121 N DUP 10
SRR1766467.7577496 chr2 231849126 N chr2 231849256 N DEL 10
SRR1766478.3148213 chr2 231849126 N chr2 231849256 N DEL 10
SRR1766445.8053166 chr2 231848976 N chr2 231849233 N DUP 10
SRR1766484.3077561 chr7 74053816 N chr7 74053933 N DEL 10
SRR1766458.584918 chr10 57693307 N chr10 57693432 N DEL 11
SRR1766470.3343466 chr10 57693309 N chr10 57693476 N DEL 12
SRR1766442.38684814 chr10 57693309 N chr10 57693532 N DEL 12
SRR1766474.2405713 chr10 57693309 N chr10 57693532 N DEL 12
SRR1766481.12121069 chr10 57693309 N chr10 57693476 N DEL 19
SRR1766471.10267820 chr10 57693307 N chr10 57693432 N DEL 15
SRR1766466.8655538 chr10 57693307 N chr10 57693432 N DEL 15
SRR1766448.1181766 chr10 57693310 N chr10 57693465 N DUP 12
SRR1766445.8409272 chr10 57693310 N chr10 57693465 N DUP 13
SRR1766448.10139971 chr10 57693310 N chr10 57693465 N DUP 13
SRR1766456.139808 chr10 57693408 N chr10 57693521 N DUP 11
SRR1766444.4934318 chr10 57693403 N chr10 57693470 N DUP 19
SRR1766450.7308757 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766454.6116447 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766442.38955487 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766443.2421400 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766464.10894326 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766468.3716087 chr10 57693472 N chr10 57693624 N DUP 11
SRR1766446.10530166 chr10 57693472 N chr10 57693624 N DUP 17
SRR1766442.33924965 chr10 57693472 N chr10 57693555 N DUP 19
SRR1766474.3338522 chr10 57693472 N chr10 57693555 N DUP 15
SRR1766443.2564668 chr10 57693367 N chr10 57693741 N DEL 11
SRR1766475.2287867 chr10 57693365 N chr10 57693739 N DEL 13
SRR1766463.8745275 chr10 1232482 N chr10 1232758 N DUP 10
SRR1766448.10161218 chr12 415452 N chr12 415509 N DEL 11
SRR1766443.3688781 chr12 415452 N chr12 415509 N DEL 11
SRR1766446.4119324 chr12 415452 N chr12 415509 N DEL 11
SRR1766452.4670150 chr10 133028342 N chr10 133028715 N DEL 13
SRR1766454.6476065 chr10 133028562 N chr10 133028715 N DEL 16
SRR1766466.8830080 chr10 133028636 N chr10 133028721 N DEL 13
SRR1766444.5670414 chr19 19770126 N chr19 19770360 N DEL 11
SRR1766475.4962381 chr18 47982686 N chr18 47982961 N DUP 11
SRR1766448.2953746 chr18 47982879 N chr18 47982932 N DEL 10
SRR1766478.8680833 chrX 153382734 N chrX 153382897 N DUP 15
SRR1766459.430459 chr13 29492175 N chr13 29492300 N DEL 13
SRR1766479.849787 chr16 88503535 N chr16 88503612 N DEL 14
SRR1766447.1116039 chr16 88503418 N chr16 88503612 N DEL 11
SRR1766448.7453874 chr16 88503418 N chr16 88503612 N DEL 11
SRR1766454.10387899 chr17 513777 N chr17 514376 N DEL 10
SRR1766454.8905852 chr17 513750 N chr17 513841 N DUP 15
SRR1766452.5574745 chr17 514000 N chr17 514553 N DEL 15
SRR1766474.1411407 chr17 513816 N chr17 514553 N DEL 10
SRR1766482.6382862 chr17 514092 N chr17 514507 N DEL 19
SRR1766484.10769514 chr17 514099 N chr17 514560 N DEL 10
SRR1766463.984017 chr17 513872 N chr17 514331 N DUP 10
SRR1766459.5800291 chr17 513845 N chr17 514628 N DEL 15
SRR1766459.2743242 chr17 514413 N chr17 514598 N DEL 10
SRR1766458.6279268 chr17 514397 N chr17 514582 N DEL 15
SRR1766460.8809729 chr17 514000 N chr17 514507 N DEL 17
SRR1766483.5323667 chr17 514414 N chr17 514507 N DEL 10
SRR1766471.5622111 chr17 513777 N chr17 514422 N DEL 10
SRR1766484.5300104 chr17 513777 N chr17 514422 N DEL 10
SRR1766483.9072803 chr17 513823 N chr17 514468 N DEL 10
SRR1766481.13060514 chr17 513872 N chr17 514515 N DUP 10
SRR1766464.7266408 chr17 513862 N chr17 514507 N DEL 15
SRR1766459.2533852 chr17 513819 N chr17 514510 N DEL 10
SRR1766461.6691777 chr17 513815 N chr17 514506 N DEL 10
SRR1766449.6367200 chr17 513799 N chr17 514582 N DEL 13
SRR1766445.1350308 chr17 513954 N chr17 514599 N DEL 15
SRR1766445.10318933 chr17 514000 N chr17 514645 N DEL 10
SRR1766472.7532989 chr17 513845 N chr17 514628 N DEL 10
SRR1766447.9491750 chr17 513799 N chr17 514674 N DEL 10
SRR1766460.1183346 chr17 513823 N chr17 514698 N DEL 11
SRR1766486.3899436 chr7 44307133 N chr7 44307194 N DEL 13
SRR1766483.6994981 chr7 44307045 N chr7 44307377 N DEL 13
SRR1766470.6803338 chr7 44306887 N chr7 44307377 N DEL 15
SRR1766476.5876239 chr5 107848382 N chr5 107848486 N DEL 15
SRR1766469.3822872 chr5 107848382 N chr5 107848486 N DEL 19
SRR1766442.17515044 chr20 18010659 N chr20 18010740 N DUP 15
SRR1766463.10108778 chr8 19450247 N chr8 19450302 N DEL 12
SRR1766467.10414418 chr5 173285163 N chr5 173285315 N DEL 10
SRR1766465.6205749 chr17 7176591 N chr17 7176654 N DUP 10
SRR1766467.8649616 chr3 127155601 N chr3 127155752 N DUP 10
SRR1766461.1455748 chr3 127155623 N chr3 127155916 N DEL 15
SRR1766450.5495346 chr3 127155667 N chr3 127156008 N DUP 10
SRR1766471.3912925 chr1 203781660 N chr1 203781969 N DEL 19
SRR1766464.528150 chr4 3567123 N chr4 3567235 N DUP 10
SRR1766477.11461267 chr1 194303954 N chr1 194304032 N DUP 18
SRR1766485.7707537 chr1 194303954 N chr1 194304032 N DUP 16
SRR1766481.358894 chr1 194303954 N chr1 194304032 N DUP 14
SRR1766443.621635 chr1 194303954 N chr1 194304032 N DUP 10
SRR1766474.5845751 chr1 194303954 N chr1 194304032 N DUP 10
SRR1766480.4817582 chr1 194303954 N chr1 194304032 N DUP 10
SRR1766455.5540420 chr1 194303954 N chr1 194304032 N DUP 10
SRR1766483.2815842 chr1 194303979 N chr1 194304052 N DUP 12
SRR1766452.9978218 chr1 194303979 N chr1 194304085 N DUP 15
SRR1766454.3881683 chr1 194303979 N chr1 194304085 N DUP 17
SRR1766459.9659730 chr1 194303974 N chr1 194304084 N DUP 11
SRR1766467.8135243 chr1 194303979 N chr1 194304089 N DUP 10
SRR1766463.9385861 chr1 194303954 N chr1 194304069 N DUP 16
SRR1766445.2556709 chr1 194303979 N chr1 194304052 N DUP 14
SRR1766457.7419715 chr1 194303979 N chr1 194304052 N DUP 15
SRR1766472.5164348 chr1 194303979 N chr1 194304052 N DUP 11
SRR1766479.11822420 chr1 194303937 N chr1 194304098 N DEL 11
SRR1766454.9385242 chr1 194303938 N chr1 194304099 N DEL 10
SRR1766456.3353895 chr15 99538164 N chr15 99538229 N DUP 12
SRR1766471.7649534 chr15 99538217 N chr15 99538328 N DUP 17
SRR1766462.7051149 chr3 53220698 N chr3 53220773 N DUP 10
SRR1766450.2468939 chr3 53220693 N chr3 53220768 N DUP 11
SRR1766445.3229622 chr3 53220693 N chr3 53220768 N DUP 11
SRR1766473.10806054 chr3 53220693 N chr3 53220768 N DUP 17
SRR1766455.9494665 chr4 151732108 N chr4 151732201 N DUP 11
SRR1766483.8017323 chr4 151732125 N chr4 151732219 N DUP 14
SRR1766449.5351571 chr4 151732125 N chr4 151732219 N DUP 15
SRR1766473.7014302 chr14 41808350 N chr14 41808476 N DUP 10
SRR1766452.6164498 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766471.697922 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766479.11559321 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766476.222021 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766484.7408776 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766478.338504 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766463.2790873 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766480.7357442 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766485.12066027 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766485.10768909 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766457.6262873 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766458.9287330 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766481.3283283 chr3 60860671 N chr3 60860889 N DEL 10
SRR1766483.5993109 chr3 60860671 N chr3 60860889 N DEL 13
SRR1766448.1799644 chr3 60860671 N chr3 60860889 N DEL 14
SRR1766462.4903994 chr3 60860671 N chr3 60860889 N DEL 14
SRR1766471.11733694 chr3 60860671 N chr3 60860889 N DEL 15
SRR1766462.2354933 chr3 60860671 N chr3 60860889 N DEL 15
SRR1766442.15233988 chr3 60860671 N chr3 60860889 N DEL 15
SRR1766442.38204776 chr3 60860671 N chr3 60860889 N DEL 15
SRR1766471.7923542 chr3 60860888 N chr3 60861013 N DEL 16
SRR1766465.1580462 chr3 60860800 N chr3 60860861 N DUP 12
SRR1766463.4530372 chr3 60860819 N chr3 60860911 N DUP 18
SRR1766456.4561025 chr3 60860911 N chr3 60860976 N DEL 13
SRR1766445.3556066 chr3 60860911 N chr3 60860976 N DEL 12
SRR1766451.9911731 chr3 60860911 N chr3 60860976 N DEL 12
SRR1766473.817752 chr3 60860911 N chr3 60860976 N DEL 11
SRR1766442.29031690 chr3 60860976 N chr3 60861370 N DUP 11
SRR1766442.21664132 chr3 60860976 N chr3 60861370 N DUP 10
SRR1766483.12388682 chr3 60861325 N chr3 60861374 N DUP 19
SRR1766484.5797667 chr3 60861331 N chr3 60861397 N DUP 13
SRR1766460.997619 chr3 60861331 N chr3 60861397 N DUP 14
SRR1766466.5425960 chr3 60861331 N chr3 60861397 N DUP 15
SRR1766469.4226798 chr3 60861325 N chr3 60861374 N DUP 15
SRR1766479.12526102 chr8 92949831 N chr8 92949944 N DEL 17
SRR1766442.12497524 chr8 92949831 N chr8 92949940 N DEL 13
SRR1766456.15467 chr8 92949831 N chr8 92949940 N DEL 13
SRR1766471.7744362 chr8 92949831 N chr8 92949944 N DEL 17
SRR1766459.281501 chr8 92949831 N chr8 92949944 N DEL 17
SRR1766483.8249271 chr8 92949831 N chr8 92949940 N DEL 13
SRR1766442.1491400 chr8 92949831 N chr8 92949944 N DEL 17
SRR1766482.12930706 chr8 92949831 N chr8 92949940 N DEL 13
SRR1766442.26922800 chr8 92949950 N chr8 92950062 N DUP 12
SRR1766467.553454 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766454.3934622 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766452.5436474 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766470.2893510 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766462.3998730 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766464.709182 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766448.630881 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766442.44025291 chr9 137346675 N chr9 137346755 N DUP 12
SRR1766466.5871898 chr9 137346675 N chr9 137346755 N DUP 15
SRR1766442.9207384 chr9 137346675 N chr9 137346755 N DUP 15
SRR1766452.5061677 chr9 137346675 N chr9 137346755 N DUP 17
SRR1766459.11523964 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766465.485204 chr9 137346675 N chr9 137346755 N DUP 14
SRR1766465.8611863 chr9 137346675 N chr9 137346755 N DUP 16
SRR1766473.438832 chr9 137346675 N chr9 137346755 N DUP 18
SRR1766451.3158204 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766450.9886743 chr9 137346675 N chr9 137346755 N DUP 11
SRR1766486.1270104 chr9 137346675 N chr9 137346755 N DUP 17
SRR1766477.4644375 chr9 137346675 N chr9 137346755 N DUP 18
SRR1766455.4979907 chr16 89118096 N chr16 89118368 N DEL 10
SRR1766465.11264477 chr1 246783161 N chr1 246783272 N DEL 12
SRR1766461.4373721 chr1 246783161 N chr1 246783272 N DEL 12
SRR1766474.6356817 chr1 246783144 N chr1 246783255 N DEL 10
SRR1766469.2045721 chr1 246783161 N chr1 246783272 N DEL 12
SRR1766447.11089647 chr1 246783161 N chr1 246783272 N DEL 12
SRR1766479.11196940 chr1 246783658 N chr1 246783711 N DUP 10
SRR1766468.3913814 chr22 35343026 N chr22 35343145 N DEL 10
SRR1766480.607020 chr22 35343029 N chr22 35343148 N DEL 10
SRR1766483.4128890 chr22 35342943 N chr22 35343108 N DUP 10
SRR1766443.5069973 chr22 35343444 N chr22 35343562 N DUP 15
SRR1766475.1516000 chr22 35343444 N chr22 35343562 N DUP 18
SRR1766477.768154 chr22 35343353 N chr22 35343471 N DUP 19
SRR1766469.858437 chr22 35343444 N chr22 35343562 N DUP 13
SRR1766469.5288738 chr2 117643589 N chr2 117643669 N DEL 13
SRR1766467.4962233 chr2 117643589 N chr2 117643669 N DEL 14
SRR1766484.7938859 chr2 117643589 N chr2 117643669 N DEL 14
SRR1766450.4983810 chr2 117643600 N chr2 117643742 N DEL 15
SRR1766442.41170099 chr2 117643612 N chr2 117643669 N DEL 13
SRR1766447.7657057 chr2 117643581 N chr2 117643651 N DUP 14
SRR1766475.321428 chr2 117643581 N chr2 117643651 N DUP 14
SRR1766473.6403983 chr2 117643588 N chr2 117643663 N DUP 18
SRR1766443.6199221 chr2 117643583 N chr2 117643643 N DEL 10
SRR1766442.37490237 chr2 117643666 N chr2 117643743 N DEL 13
SRR1766459.7648564 chr7 98242710 N chr7 98242916 N DEL 10
SRR1766449.1934320 chr7 98242677 N chr7 98243204 N DUP 10
SRR1766450.10299331 chr7 98242740 N chr7 98242950 N DEL 16
SRR1766466.6080538 chr7 98242740 N chr7 98242950 N DEL 10
SRR1766451.8430121 chr7 98242722 N chr7 98242888 N DEL 10
SRR1766451.8963773 chr7 98242720 N chr7 98242882 N DEL 14
SRR1766483.2533620 chr7 98242585 N chr7 98242932 N DEL 10
SRR1766486.5729006 chr7 98242680 N chr7 98243069 N DUP 17
SRR1766445.3465306 chr7 98242680 N chr7 98243069 N DUP 17
SRR1766459.5195443 chr7 98242680 N chr7 98243069 N DUP 17
SRR1766445.3465306 chr7 98242710 N chr7 98243099 N DUP 16
SRR1766481.2920189 chr7 98242680 N chr7 98243069 N DUP 17
SRR1766472.319119 chr7 98242631 N chr7 98243010 N DEL 10
SRR1766483.4972764 chr7 98243151 N chr7 98243236 N DEL 13
SRR1766445.2933269 chr7 98242933 N chr7 98243125 N DUP 10
SRR1766460.7656836 chr7 98243143 N chr7 98243197 N DUP 13
SRR1766475.8964712 chr7 98242588 N chr7 98243186 N DEL 11
SRR1766461.4851364 chr7 98242859 N chr7 98243215 N DEL 10
SRR1766478.7636865 chr7 98242583 N chr7 98243245 N DEL 15
SRR1766442.34405836 chr14 105693685 N chr14 105693776 N DUP 13
SRR1766456.1765955 chr14 105693591 N chr14 105693682 N DEL 13
SRR1766469.1574397 chr14 105693724 N chr14 105693849 N DUP 13
SRR1766483.10386505 chr14 105693724 N chr14 105693849 N DUP 13
SRR1766482.6452191 chr14 105693685 N chr14 105693776 N DUP 18
SRR1766467.6138329 chr14 105693767 N chr14 105693898 N DEL 13
SRR1766456.1765955 chr14 105693767 N chr14 105693898 N DEL 13
SRR1766480.7451536 chr14 105693767 N chr14 105693898 N DEL 13
SRR1766470.5418221 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766453.1635179 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766461.3897103 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766482.7587429 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766447.6165974 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766460.2399364 chr14 105693624 N chr14 105693991 N DUP 15
SRR1766466.2330993 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766483.2379837 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766463.1477430 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766462.3769719 chr14 105694008 N chr14 105694175 N DEL 12
SRR1766474.1253906 chr14 105693764 N chr14 105693993 N DUP 14
SRR1766479.848576 chr14 105693636 N chr14 105693899 N DEL 13
SRR1766442.15504051 chr14 105693640 N chr14 105693903 N DEL 10
SRR1766474.3952943 chr14 105693488 N chr14 105693904 N DUP 11
SRR1766442.2051280 chr14 105694118 N chr14 105694245 N DEL 10
SRR1766456.5459490 chr14 105694201 N chr14 105694410 N DEL 15
SRR1766442.40990022 chr14 105693788 N chr14 105694750 N DUP 15
SRR1766446.2603995 chr14 105694158 N chr14 105694860 N DUP 10
SRR1766442.30736685 chr11 38147208 N chr11 38147263 N DUP 10
SRR1766458.8687225 chr1 2977522 N chr1 2978110 N DEL 11
SRR1766475.1560710 chr14 100546488 N chr14 100546608 N DEL 15
SRR1766453.128358 chr7 62441836 N chr7 62442285 N DEL 15
SRR1766447.3670339 chr7 62442456 N chr7 62442751 N DEL 15
SRR1766465.11230860 chr7 62441916 N chr7 62442590 N DEL 10
SRR1766478.191833 chr7 62441916 N chr7 62442590 N DEL 10
SRR1766442.698419 chr2 206372218 N chr2 206372321 N DEL 12
SRR1766453.5812362 chr2 206372218 N chr2 206372321 N DEL 12
SRR1766454.9060274 chr2 206372220 N chr2 206372323 N DEL 10
SRR1766453.5600855 chr2 206372218 N chr2 206372321 N DEL 12
SRR1766479.2594768 chr4 70516460 N chr4 70516561 N DEL 10
SRR1766462.776988 chr4 70516460 N chr4 70516561 N DEL 12
SRR1766473.10455670 chr4 70516460 N chr4 70516561 N DEL 13
SRR1766466.5291348 chr4 70516459 N chr4 70516538 N DEL 18
SRR1766464.1177064 chr4 70516455 N chr4 70516556 N DEL 13
SRR1766485.7186165 chr4 70516455 N chr4 70516556 N DEL 13
SRR1766473.808173 chr4 70516455 N chr4 70516564 N DEL 10
SRR1766442.8935067 chr2 64375803 N chr2 64375868 N DEL 13
SRR1766470.4626732 chr2 64375858 N chr2 64376377 N DEL 13
SRR1766456.6162646 chr2 64375868 N chr2 64375952 N DUP 19
SRR1766479.1785907 chr2 64375822 N chr2 64375950 N DUP 11
SRR1766478.3040180 chr2 64375800 N chr2 64376035 N DEL 19
SRR1766482.4175847 chr2 64375740 N chr2 64375815 N DUP 10
SRR1766443.8429926 chr2 64375748 N chr2 64375917 N DUP 17
SRR1766479.12516280 chr2 64375838 N chr2 64376193 N DEL 13
SRR1766476.2181495 chr2 64375766 N chr2 64376092 N DEL 18
SRR1766456.1368625 chr2 64375800 N chr2 64375880 N DEL 13
SRR1766447.7497881 chr2 64375897 N chr2 64376202 N DEL 11
SRR1766482.10989921 chr2 64375749 N chr2 64375876 N DEL 10
SRR1766469.1311668 chr2 64376173 N chr2 64376289 N DUP 13
SRR1766466.2982883 chr2 64375915 N chr2 64376221 N DUP 10
SRR1766467.11058203 chr2 64375918 N chr2 64376069 N DUP 11
SRR1766463.318073 chr2 64375874 N chr2 64376338 N DUP 13
SRR1766446.8520773 chr2 64375900 N chr2 64375975 N DUP 10
SRR1766447.4097105 chr2 64375735 N chr2 64375977 N DUP 18
SRR1766473.8323290 chr2 64375797 N chr2 64376187 N DEL 11
SRR1766483.6953215 chr2 64375747 N chr2 64375989 N DUP 11
SRR1766445.8500216 chr2 64375828 N chr2 64376345 N DUP 13
SRR1766476.9592672 chr2 64375874 N chr2 64375952 N DUP 13
SRR1766465.992677 chr2 64375874 N chr2 64375990 N DUP 16
SRR1766469.8584880 chr2 64375874 N chr2 64376338 N DUP 13
SRR1766478.10710367 chr2 64375944 N chr2 64376173 N DEL 13
SRR1766456.5515521 chr2 64375874 N chr2 64376069 N DUP 10
SRR1766453.3260526 chr2 64375824 N chr2 64376016 N DUP 11
SRR1766477.3223782 chr2 64375736 N chr2 64376086 N DUP 16
SRR1766480.3121727 chr2 64375825 N chr2 64376017 N DUP 10
SRR1766452.4615466 chr2 64375874 N chr2 64375990 N DUP 10
SRR1766476.6838937 chr2 64375874 N chr2 64376256 N DUP 14
SRR1766442.7354464 chr2 64375874 N chr2 64375987 N DUP 13
SRR1766478.9075524 chr2 64375886 N chr2 64376347 N DUP 10
SRR1766456.3795525 chr2 64375874 N chr2 64375990 N DUP 10
SRR1766453.3864471 chr2 64375874 N chr2 64375990 N DUP 10
SRR1766480.4931241 chr2 64375874 N chr2 64375987 N DUP 13
SRR1766446.5563350 chr2 64375868 N chr2 64375952 N DUP 11
SRR1766452.8880707 chr2 64375780 N chr2 64376208 N DEL 16
SRR1766481.3941539 chr2 64375737 N chr2 64376093 N DUP 13
SRR1766453.3880162 chr2 64375795 N chr2 64376145 N DUP 12
SRR1766455.3219840 chr2 64375944 N chr2 64376135 N DEL 11
SRR1766472.3668981 chr2 64375782 N chr2 64375874 N DEL 11
SRR1766469.11046682 chr2 64375747 N chr2 64375989 N DUP 18
SRR1766458.1451090 chr2 64375737 N chr2 64375856 N DUP 13
SRR1766481.9487105 chr2 64375791 N chr2 64375874 N DEL 13
SRR1766456.5934369 chr2 64375737 N chr2 64375979 N DUP 18
SRR1766479.3600612 chr2 64375884 N chr2 64376218 N DEL 15
SRR1766455.8841869 chr2 64376174 N chr2 64376290 N DUP 10
SRR1766457.4284435 chr2 64375737 N chr2 64375979 N DUP 15
SRR1766448.10928298 chr2 64375812 N chr2 64375975 N DUP 13
SRR1766469.6997753 chr2 64375737 N chr2 64375979 N DUP 17
SRR1766452.8798532 chr2 64375801 N chr2 64376344 N DUP 13
SRR1766472.5977698 chr2 64375807 N chr2 64376116 N DUP 11
SRR1766483.11075530 chr2 64375795 N chr2 64376069 N DUP 13
SRR1766485.7896807 chr2 64375944 N chr2 64376018 N DEL 16
SRR1766442.31898883 chr2 64375838 N chr2 64376231 N DEL 16
SRR1766445.9821722 chr2 64376005 N chr2 64376193 N DEL 10
SRR1766447.8266882 chr2 64375758 N chr2 64376310 N DUP 12
SRR1766484.31648 chr2 64375944 N chr2 64376018 N DEL 12
SRR1766447.8266882 chr2 64375759 N chr2 64376308 N DUP 14
SRR1766484.10428003 chr2 64375746 N chr2 64376295 N DUP 11
SRR1766450.8013720 chr2 64375862 N chr2 64376173 N DEL 10
SRR1766448.3886690 chr2 64375874 N chr2 64376297 N DUP 17
SRR1766479.4471343 chr2 64375874 N chr2 64376145 N DUP 18
SRR1766463.1685291 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766478.6116256 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766481.409521 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766463.2518470 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766445.4818764 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766449.5423178 chr2 94283690 N chr2 94283788 N DEL 10
SRR1766462.10448532 chrX 35692503 N chrX 35692560 N DUP 19
SRR1766479.9065739 chrX 35692503 N chrX 35692560 N DUP 16
SRR1766482.12448661 chrX 35692503 N chrX 35692610 N DUP 19
SRR1766442.25600171 chrX 35692503 N chrX 35692610 N DUP 19
SRR1766442.1184542 chrX 1472802 N chrX 1472960 N DUP 12
SRR1766451.9472057 chrX 1473000 N chrX 1473199 N DEL 13
SRR1766482.6957216 chrX 1472867 N chrX 1473034 N DUP 11
SRR1766445.4822830 chrX 1473013 N chrX 1473139 N DUP 15
SRR1766454.8447095 chr1 8301356 N chr1 8301441 N DEL 10
SRR1766452.5510176 chr1 8301356 N chr1 8301441 N DEL 12
SRR1766450.6225578 chr1 8301482 N chr1 8301931 N DEL 11
SRR1766474.4394840 chr1 8301462 N chr1 8301659 N DEL 10
SRR1766447.1099627 chr1 8301430 N chr1 8301851 N DEL 10
SRR1766457.5066481 chr1 8301505 N chr1 8301926 N DEL 11
SRR1766467.3794240 chr1 8301437 N chr1 8301548 N DUP 13
SRR1766480.2029925 chr1 8301505 N chr1 8301588 N DUP 10
SRR1766471.2724162 chr1 8301428 N chr1 8301567 N DUP 10
SRR1766454.847125 chr1 8301542 N chr1 8301961 N DUP 10
SRR1766466.9790793 chr1 8301634 N chr1 8301915 N DEL 10
SRR1766477.9827703 chr1 8301653 N chr1 8301960 N DUP 10
SRR1766485.4436147 chr1 8301393 N chr1 8301758 N DEL 10
SRR1766485.4460136 chr1 8301589 N chr1 8301758 N DEL 12
SRR1766442.4413872 chr1 8301781 N chr1 8301948 N DUP 15
SRR1766463.6086776 chr1 8301586 N chr1 8301783 N DEL 12
SRR1766486.8460964 chr1 8301502 N chr1 8301783 N DEL 10
SRR1766442.40547766 chr1 8301486 N chr1 8301851 N DEL 16
SRR1766454.5673377 chr1 8301486 N chr1 8301851 N DEL 16
SRR1766475.8036736 chr1 8301709 N chr1 8301878 N DEL 11
SRR1766474.8666197 chr1 8301541 N chr1 8301878 N DEL 10
SRR1766467.5122452 chr1 8301389 N chr1 8302033 N DEL 10
SRR1766458.3312228 chr8 132187932 N chr8 132188029 N DEL 10
SRR1766451.5424159 chr8 132187947 N chr8 132188000 N DUP 10
SRR1766485.4977296 chr8 132187791 N chr8 132188011 N DEL 14
SRR1766484.7598318 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766476.5880276 chr5 180615360 N chr5 180615464 N DEL 15
SRR1766456.6470003 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766452.7138667 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766472.2125366 chr5 180615386 N chr5 180615548 N DEL 10
SRR1766447.2809373 chr5 180615335 N chr5 180615437 N DUP 13
SRR1766442.9426009 chr5 180615317 N chr5 180615522 N DUP 15
SRR1766448.1807269 chr5 180615318 N chr5 180615420 N DUP 10
SRR1766442.3611502 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766454.4593470 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766465.5023132 chr5 180615372 N chr5 180615521 N DEL 10
SRR1766485.11657075 chr22 18370651 N chr22 18370706 N DEL 15
SRR1766480.6806500 chr22 18370628 N chr22 18370710 N DEL 10
SRR1766469.9155466 chr2 225783072 N chr2 225783687 N DUP 12
SRR1766475.4779788 chr12 48664595 N chr12 48664900 N DEL 16
SRR1766483.1458972 chr12 48664443 N chr12 48665032 N DEL 12
SRR1766476.1026075 chr10 49105183 N chr10 49105333 N DEL 12
SRR1766473.5023340 chr15 101763542 N chr15 101763634 N DEL 10
SRR1766471.4159492 chr15 101763538 N chr15 101763816 N DUP 10
SRR1766444.3613729 chr15 101763835 N chr15 101763990 N DUP 15
SRR1766457.8535198 chr15 101763708 N chr15 101764045 N DUP 15
SRR1766476.8083468 chr2 91411569 N chr2 91411720 N DEL 12
SRR1766457.6475972 chr2 91411569 N chr2 91411720 N DEL 14
SRR1766482.7385798 chr2 91411561 N chr2 91411637 N DEL 15
SRR1766442.9203551 chr2 91411561 N chr2 91411637 N DEL 16
SRR1766442.5604741 chr2 91411561 N chr2 91411637 N DEL 16
SRR1766442.8615401 chr2 91411589 N chr2 91411642 N DEL 14
SRR1766442.28051979 chr2 91411589 N chr2 91411642 N DEL 14
SRR1766442.45350726 chr2 91411600 N chr2 91411653 N DEL 10
SRR1766450.9897887 chr2 91411600 N chr2 91411653 N DEL 11
SRR1766456.5372149 chr2 91411600 N chr2 91411653 N DEL 12
SRR1766462.84490 chr2 91411600 N chr2 91411653 N DEL 12
SRR1766442.474109 chr13 99620946 N chr13 99620995 N DUP 10
SRR1766464.5004418 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766464.1312386 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766462.11166545 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766470.8699690 chr10 58708156 N chr10 58708299 N DEL 16
SRR1766454.8558581 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766472.11610492 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766443.4177231 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766449.3936321 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766483.2040401 chr6 36364101 N chr6 36364262 N DEL 10
SRR1766449.5793786 chr13 18468420 N chr13 18469084 N DEL 14
SRR1766479.7061399 chr10 83585215 N chr10 83585312 N DEL 13
SRR1766443.4056017 chr10 83585260 N chr10 83585312 N DEL 19
SRR1766465.9769986 chr10 83585215 N chr10 83585312 N DEL 12
SRR1766447.9802070 chr10 83585216 N chr10 83585313 N DEL 12
SRR1766472.9956458 chr10 83585264 N chr10 83585316 N DEL 11
SRR1766467.11122595 chr17 41123891 N chr17 41124132 N DEL 10
SRR1766469.5487914 chr17 41123891 N chr17 41124132 N DEL 10
SRR1766453.8800494 chr17 41123891 N chr17 41124132 N DEL 10
SRR1766454.218979 chr17 41123891 N chr17 41124132 N DEL 10
SRR1766474.9424075 chr17 10475742 N chr17 10475797 N DUP 19
SRR1766455.5567930 chr7 111539297 N chr7 111539354 N DEL 15
SRR1766463.1755430 chr19 53559050 N chr19 53559157 N DUP 17
SRR1766475.5827848 chr19 53559050 N chr19 53559157 N DUP 16
SRR1766482.11081530 chr19 53559050 N chr19 53559157 N DUP 16
SRR1766443.4797883 chr1 191828617 N chr1 191828736 N DEL 14
SRR1766452.8612104 chr1 191828611 N chr1 191828736 N DEL 14
SRR1766466.5250270 chr1 191828611 N chr1 191828738 N DEL 13
SRR1766461.3313195 chr22 32330694 N chr22 32330952 N DEL 10
SRR1766469.7646005 chr22 32330227 N chr22 32331116 N DUP 10
SRR1766484.3511511 chr22 32330744 N chr22 32331014 N DEL 11
SRR1766452.4833591 chr22 32329821 N chr22 32331337 N DEL 11
SRR1766471.10757781 chr13 84125790 N chr13 84125882 N DUP 10
SRR1766450.5530687 chr10 110411888 N chr10 110411961 N DUP 13
SRR1766451.9033452 chr9 89671689 N chr9 89671819 N DEL 18
SRR1766483.11646071 chr9 89671698 N chr9 89671748 N DUP 15
SRR1766442.15415282 chr9 89671740 N chr9 89671895 N DUP 15
SRR1766450.81952 chr9 89671770 N chr9 89671826 N DUP 19
SRR1766483.186203 chr9 89671770 N chr9 89671877 N DUP 17
SRR1766465.3894362 chr9 89671698 N chr9 89671808 N DUP 18
SRR1766442.43397043 chr9 89671656 N chr9 89671793 N DUP 13
SRR1766442.31375677 chr9 89671738 N chr9 89671923 N DUP 10
SRR1766442.34575855 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766453.6777803 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766442.3282057 chr9 89671713 N chr9 89671769 N DUP 17
SRR1766474.9109956 chr9 89671692 N chr9 89671802 N DUP 14
SRR1766468.7418887 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766462.6278994 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766467.648867 chr9 89671742 N chr9 89671945 N DUP 10
SRR1766460.2499286 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766482.10510174 chr9 89671701 N chr9 89671850 N DUP 15
SRR1766479.889896 chr9 89671755 N chr9 89671859 N DUP 12
SRR1766445.3147857 chr9 89671755 N chr9 89671859 N DUP 12
SRR1766472.10619239 chr9 89671713 N chr9 89671769 N DUP 17
SRR1766458.2726627 chr9 89671692 N chr9 89671802 N DUP 14
SRR1766468.6203617 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766453.4804902 chr9 89671692 N chr9 89671802 N DUP 19
SRR1766442.36499330 chr9 89671729 N chr9 89671833 N DUP 10
SRR1766460.6361669 chr9 89671729 N chr9 89671833 N DUP 15
SRR1766472.1245181 chr9 89671771 N chr9 89671878 N DUP 17
SRR1766470.5022487 chr9 89671692 N chr9 89671802 N DUP 19
SRR1766484.3901896 chr9 89671729 N chr9 89671782 N DUP 15
SRR1766471.11994022 chr9 89671701 N chr9 89671859 N DUP 17
SRR1766473.6578963 chr9 89671698 N chr9 89671775 N DUP 17
SRR1766466.9088531 chr9 89671701 N chr9 89671859 N DUP 19
SRR1766471.2137093 chr9 89671705 N chr9 89671812 N DUP 10
SRR1766447.2003579 chr9 89671692 N chr9 89671853 N DUP 11
SRR1766450.1914612 chr9 89671792 N chr9 89671878 N DUP 12
SRR1766483.8401693 chr9 89671818 N chr9 89671874 N DUP 19
SRR1766457.3867954 chr9 89671720 N chr9 89671793 N DEL 12
SRR1766447.10681820 chr9 89671690 N chr9 89671935 N DUP 17
SRR1766442.17130031 chr9 89671743 N chr9 89671841 N DUP 12
SRR1766456.5141629 chr9 89671829 N chr9 89671881 N DEL 10
SRR1766485.3052228 chr9 89671724 N chr9 89671884 N DEL 12
SRR1766444.4934578 chr6 89125933 N chr6 89126832 N DUP 11
SRR1766443.9191301 chr22 48858144 N chr22 48858243 N DUP 10
SRR1766463.7196809 chr22 36434243 N chr22 36434385 N DUP 12
SRR1766458.1222399 chr22 36434323 N chr22 36434386 N DUP 10
SRR1766442.4509105 chr22 36434260 N chr22 36434359 N DEL 10
SRR1766478.6579743 chr22 36434260 N chr22 36434359 N DEL 10
SRR1766477.7379421 chr1 96153244 N chr1 96153309 N DUP 12
SRR1766481.6612261 chr1 96153244 N chr1 96153309 N DUP 13
SRR1766442.24511617 chr1 96153244 N chr1 96153309 N DUP 19
SRR1766448.3634630 chr1 96153244 N chr1 96153309 N DUP 18
SRR1766463.3962757 chr1 96153244 N chr1 96153309 N DUP 18
SRR1766456.5549548 chrX 143492665 N chrX 143492759 N DEL 10
SRR1766445.3944385 chr11 82625239 N chr11 82625701 N DUP 11
SRR1766448.4917194 chr11 82625239 N chr11 82625701 N DUP 12
SRR1766450.2529431 chr11 82625268 N chr11 82625639 N DEL 15
SRR1766470.10170800 chr1 67930134 N chr1 67930185 N DEL 16
SRR1766442.28711279 chr1 67930132 N chr1 67930188 N DEL 12
SRR1766459.4334118 chr1 67930132 N chr1 67930188 N DEL 12
SRR1766442.36425228 chr1 67930133 N chr1 67930189 N DEL 11
SRR1766453.453629 chr6 64296679 N chr6 64296774 N DEL 13
SRR1766474.10119312 chr6 64296679 N chr6 64296774 N DEL 13
SRR1766442.31667097 chr18 79631143 N chr18 79631305 N DUP 10
SRR1766468.4850778 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766463.3065180 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766472.12030894 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766482.6565003 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766459.2999629 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766474.1018088 chr20 22378591 N chr20 22378658 N DEL 14
SRR1766442.4714973 chr20 22378591 N chr20 22378658 N DEL 15
SRR1766448.10370720 chr20 22378581 N chr20 22378638 N DEL 15
SRR1766463.7254966 chr20 22378615 N chr20 22378744 N DEL 12
SRR1766461.1932418 chr11 132162754 N chr11 132162869 N DUP 18
SRR1766459.2603290 chr2 5172401 N chr2 5172504 N DUP 10
SRR1766464.6095762 chr2 5172452 N chr2 5172521 N DUP 10
SRR1766451.2656153 chr2 5172441 N chr2 5172667 N DUP 14
SRR1766458.5366035 chr2 5172479 N chr2 5172548 N DUP 11
SRR1766464.5250533 chr2 5172442 N chr2 5172738 N DUP 13
SRR1766485.7867618 chr2 5172442 N chr2 5172738 N DUP 14
SRR1766482.7999140 chr2 5172442 N chr2 5172738 N DUP 15
SRR1766465.4066721 chr2 5172453 N chr2 5172819 N DUP 10
SRR1766478.6416402 chr4 1652212 N chr4 1652711 N DEL 15
SRR1766483.10468105 chr4 1652233 N chr4 1652733 N DEL 12
SRR1766444.3148256 chr4 1652332 N chr4 1652384 N DEL 10
SRR1766450.10170017 chr4 1652285 N chr4 1652595 N DUP 12
SRR1766442.32025554 chr4 1652385 N chr4 1652752 N DUP 11
SRR1766475.8193333 chr4 1652624 N chr4 1652788 N DUP 12
SRR1766442.20982458 chr4 1652791 N chr4 1652929 N DEL 11
SRR1766477.5301882 chr5 29743712 N chr5 29743790 N DUP 12
SRR1766465.9281932 chr10 17629553 N chr10 17629750 N DEL 10
SRR1766462.7797835 chr6 104424368 N chr6 104424501 N DEL 11
SRR1766442.967555 chr6 104424329 N chr6 104424462 N DEL 18
SRR1766473.4522759 chr6 104424329 N chr6 104424462 N DEL 18
SRR1766445.8931811 chr6 104424329 N chr6 104424462 N DEL 18
SRR1766444.532132 chr6 104424448 N chr6 104424549 N DEL 16
SRR1766464.8385957 chr6 104424385 N chr6 104424566 N DEL 13
SRR1766485.9612350 chr6 104424385 N chr6 104424566 N DEL 13
SRR1766483.517225 chr6 104424385 N chr6 104424566 N DEL 13
SRR1766457.1495452 chr3 122780252 N chr3 122780351 N DEL 10
SRR1766486.4183173 chr3 122780546 N chr3 122780721 N DEL 10
SRR1766483.6427839 chr3 122780546 N chr3 122780721 N DEL 15
SRR1766477.6589296 chr3 181743074 N chr3 181743217 N DEL 16
SRR1766482.795057 chr3 181743062 N chr3 181743157 N DEL 15
SRR1766466.1381218 chr15 84672895 N chr15 84673012 N DEL 13
SRR1766461.475316 chrY 10750602 N chrY 10750701 N DUP 10
SRR1766447.5041538 chr19 108019 N chr19 108076 N DUP 12
SRR1766477.4433814 chr19 108019 N chr19 108076 N DUP 14
SRR1766458.3282239 chr19 108015 N chr19 108082 N DUP 10
SRR1766478.10914553 chr19 108120 N chr19 108206 N DEL 12
SRR1766465.7444298 chr19 108043 N chr19 108100 N DEL 18
SRR1766442.26622570 chr19 108120 N chr19 108206 N DEL 12
SRR1766442.24412388 chr19 108120 N chr19 108206 N DEL 12
SRR1766442.18570184 chr19 108076 N chr19 108245 N DUP 17
SRR1766482.10962747 chr19 108014 N chr19 108167 N DUP 19
SRR1766451.2923848 chr19 108014 N chr19 108167 N DUP 19
SRR1766453.3918307 chr19 108014 N chr19 108167 N DUP 19
SRR1766453.3911643 chr19 107913 N chr19 108087 N DEL 11
SRR1766453.10539642 chr19 108118 N chr19 108200 N DUP 10
SRR1766449.10487788 chr6 38103619 N chr6 38103674 N DEL 13
SRR1766474.6505441 chr6 38103619 N chr6 38103674 N DEL 13
SRR1766473.1415475 chr6 38103619 N chr6 38103674 N DEL 14
SRR1766444.4120140 chr7 47736367 N chr7 47736539 N DUP 15
SRR1766473.8540541 chrX 30602965 N chrX 30603420 N DUP 10
SRR1766448.8688647 chrX 30603179 N chrX 30603404 N DUP 12
SRR1766456.1890393 chrX 30602889 N chrX 30603245 N DUP 10
SRR1766462.7762510 chrX 30602984 N chrX 30603391 N DEL 11
SRR1766451.858048 chr6 25206655 N chr6 25206732 N DUP 13
SRR1766466.4973155 chr6 25206655 N chr6 25206732 N DUP 15
SRR1766476.4947481 chr6 25206644 N chr6 25206699 N DUP 13
SRR1766442.47090403 chr6 25206702 N chr6 25206775 N DUP 17
SRR1766447.8831279 chr6 25206659 N chr6 25206737 N DEL 11
SRR1766465.4195719 chr6 25206657 N chr6 25206767 N DEL 16
SRR1766483.11930667 chr6 25206657 N chr6 25206767 N DEL 16
SRR1766442.46609057 chrX 114387100 N chrX 114387232 N DEL 11
SRR1766462.3490905 chrX 114387100 N chrX 114387232 N DEL 11
SRR1766473.11346133 chrX 114387100 N chrX 114387232 N DEL 13
SRR1766442.31322311 chrX 114387100 N chrX 114387232 N DEL 18
SRR1766467.11197680 chrX 114387100 N chrX 114387232 N DEL 19
SRR1766481.10066704 chrX 114387100 N chrX 114387232 N DEL 12
SRR1766471.10706270 chrX 114387100 N chrX 114387232 N DEL 19
SRR1766482.10018456 chrX 114387045 N chrX 114387176 N DUP 10
SRR1766462.10247388 chrX 114387129 N chrX 114387595 N DEL 11
SRR1766442.45939718 chrX 114387042 N chrX 114387195 N DUP 11
SRR1766442.43858060 chrX 114387075 N chrX 114387475 N DEL 10
SRR1766479.2283950 chrX 114387120 N chrX 114387406 N DEL 19
SRR1766485.943342 chrX 114387063 N chrX 114387387 N DUP 18
SRR1766470.1011863 chrX 114387178 N chrX 114387241 N DEL 11
SRR1766482.8774494 chrX 114387178 N chrX 114387241 N DEL 11
SRR1766453.9217813 chrX 114387182 N chrX 114387266 N DUP 17
SRR1766462.3490905 chrX 114387198 N chrX 114387299 N DEL 14
SRR1766460.6309865 chrX 114387244 N chrX 114387566 N DUP 18
SRR1766472.10854182 chrX 114387221 N chrX 114387385 N DUP 19
SRR1766454.2139521 chrX 114387265 N chrX 114387320 N DUP 12
SRR1766442.5682528 chrX 114387261 N chrX 114387336 N DUP 19
SRR1766481.9076653 chrX 114387221 N chrX 114387385 N DUP 13
SRR1766442.44913756 chrX 114387315 N chrX 114387541 N DEL 17
SRR1766447.1511369 chrX 114387258 N chrX 114387323 N DEL 13
SRR1766472.8561265 chrX 114387175 N chrX 114387342 N DEL 14
SRR1766462.10247388 chrX 114387053 N chrX 114387357 N DUP 14
SRR1766443.7709385 chrX 114387321 N chrX 114387505 N DEL 17
SRR1766443.992595 chrX 114387199 N chrX 114387385 N DUP 12
SRR1766442.12813109 chrX 114387199 N chrX 114387385 N DUP 13
SRR1766461.10309545 chrX 114387324 N chrX 114387503 N DEL 12
SRR1766486.1008721 chrX 114387199 N chrX 114387385 N DUP 13
SRR1766442.22025397 chrX 114387063 N chrX 114387366 N DUP 10
SRR1766460.4809186 chrX 114387199 N chrX 114387385 N DUP 13
SRR1766454.5525715 chrX 114387199 N chrX 114387385 N DUP 16
SRR1766465.10827398 chrX 114387199 N chrX 114387385 N DUP 17
SRR1766467.864445 chrX 114387178 N chrX 114387299 N DEL 11
SRR1766477.8918353 chrX 114387080 N chrX 114387323 N DEL 16
SRR1766459.6544722 chrX 114387281 N chrX 114387376 N DUP 16
SRR1766455.4469180 chrX 114387089 N chrX 114387297 N DEL 11
SRR1766473.7390007 chrX 114387258 N chrX 114387341 N DEL 15
SRR1766486.1274959 chrX 114387247 N chrX 114387403 N DUP 17
SRR1766473.9805277 chrX 114387339 N chrX 114387392 N DUP 10
SRR1766443.10125434 chrX 114387120 N chrX 114387406 N DEL 19
SRR1766450.6363542 chrX 114387221 N chrX 114387385 N DUP 11
SRR1766467.9461684 chrX 114387115 N chrX 114387497 N DUP 11
SRR1766469.1993856 chrX 114387221 N chrX 114387385 N DUP 19
SRR1766480.3075486 chrX 114387378 N chrX 114387533 N DEL 16
SRR1766445.8908361 chrX 114387352 N chrX 114387576 N DEL 17
SRR1766482.4114782 chr8 140120705 N chr8 140120870 N DEL 12
SRR1766477.6411351 chr22 11330112 N chr22 11330207 N DUP 10
SRR1766461.1126524 chr22 11330112 N chr22 11330207 N DUP 10
SRR1766442.10339754 chr22 11330119 N chr22 11330214 N DUP 14
SRR1766442.46585745 chr22 11330120 N chr22 11330215 N DUP 12
SRR1766453.3022385 chr22 11330119 N chr22 11330214 N DUP 14
SRR1766455.2889090 chr22 11330122 N chr22 11330217 N DUP 10
SRR1766465.9343204 chr22 11330119 N chr22 11330214 N DUP 13
SRR1766482.8128168 chr22 11330119 N chr22 11330214 N DUP 14
SRR1766454.6074728 chr22 11330119 N chr22 11330214 N DUP 14
SRR1766471.9921091 chr22 11330074 N chr22 11330258 N DUP 14
SRR1766446.1583450 chr22 11330127 N chr22 11330224 N DEL 10
SRR1766477.9859847 chr6 139308115 N chr6 139308166 N DEL 11
SRR1766478.979686 chr6 139308121 N chr6 139308173 N DEL 14
SRR1766462.3627008 chr6 139308114 N chr6 139308165 N DEL 19
SRR1766473.10807103 chr4 127417316 N chr4 127417375 N DEL 12
SRR1766476.9377565 chr4 127417316 N chr4 127417375 N DEL 10
SRR1766464.4648920 chr4 127417350 N chr4 127417451 N DUP 17
SRR1766447.6353005 chr10 33028397 N chr10 33028456 N DEL 12
SRR1766452.1366004 chr10 33028397 N chr10 33028456 N DEL 12
SRR1766465.6949820 chr10 33028393 N chr10 33028456 N DEL 12
SRR1766448.2835657 chr10 33028347 N chr10 33028455 N DEL 12
SRR1766461.8582858 chr2 871439 N chr2 871549 N DUP 10
SRR1766472.6523051 chr13 19779565 N chr13 19779743 N DEL 10
SRR1766477.8344625 chr13 19779565 N chr13 19779743 N DEL 14
SRR1766443.219929 chr13 19779673 N chr13 19779801 N DEL 10
SRR1766479.349534 chr13 19779673 N chr13 19779801 N DEL 10
SRR1766473.6766822 chr13 19779565 N chr13 19779743 N DEL 12
SRR1766470.5637666 chr8 138865753 N chr8 138865864 N DEL 13
SRR1766454.6765661 chr8 138865768 N chr8 138865861 N DEL 10
SRR1766486.11242618 chr12 132621012 N chr12 132621074 N DEL 10
SRR1766483.9079138 chr12 132621012 N chr12 132621074 N DEL 10
SRR1766444.871769 chr12 132621012 N chr12 132621074 N DEL 12
SRR1766454.1314268 chr12 132621012 N chr12 132621074 N DEL 15
SRR1766456.5769056 chr4 19288874 N chr4 19288965 N DUP 13
SRR1766442.10979661 chr5 69515568 N chr5 69515745 N DUP 12
SRR1766452.6884391 chr5 69515690 N chr5 69515739 N DUP 12
SRR1766477.7031888 chr5 69515689 N chr5 69515738 N DUP 15
SRR1766463.5740455 chr5 69515678 N chr5 69515776 N DUP 16
SRR1766442.21952003 chr3 127155225 N chr3 127155469 N DEL 12
SRR1766485.7810432 chr3 127155310 N chr3 127155555 N DUP 12
SRR1766480.981493 chr3 127155047 N chr3 127155597 N DEL 11
SRR1766467.8649616 chr3 127155255 N chr3 127155601 N DEL 10
SRR1766463.10639667 chr19 480778 N chr19 481549 N DEL 18
SRR1766483.4152223 chr19 480691 N chr19 480818 N DEL 14
SRR1766475.3744517 chr19 480929 N chr19 481158 N DEL 10
SRR1766472.6534139 chr19 481005 N chr19 481057 N DEL 13
SRR1766479.4817102 chr19 480992 N chr19 481586 N DEL 17
SRR1766443.6832162 chr19 481022 N chr19 481588 N DUP 15
SRR1766460.7260932 chr19 480631 N chr19 481516 N DEL 10
SRR1766486.4514432 chr19 481591 N chr19 481665 N DUP 17
SRR1766459.11167873 chr19 480653 N chr19 481649 N DUP 11
SRR1766475.3884818 chr19 481321 N chr19 481648 N DEL 18
SRR1766484.10780905 chr19 481725 N chr19 481823 N DEL 10
SRR1766457.1057925 chr11 131680982 N chr11 131681073 N DUP 14
SRR1766467.6577654 chr11 131680936 N chr11 131681081 N DUP 15
SRR1766444.700229 chr11 131681184 N chr11 131681311 N DEL 14
SRR1766465.1142782 chr11 131681142 N chr11 131681311 N DEL 19
SRR1766462.8258259 chr11 131680938 N chr11 131681267 N DUP 12
SRR1766454.2824306 chr11 131680952 N chr11 131681185 N DEL 11
SRR1766484.5088782 chr11 131680938 N chr11 131681395 N DUP 14
SRR1766482.5509295 chr11 131681134 N chr11 131681345 N DEL 10
SRR1766447.7790093 chr11 131680952 N chr11 131681319 N DEL 12
SRR1766471.2917280 chr11 131680937 N chr11 131681450 N DUP 13
SRR1766486.9741504 chr11 131681574 N chr11 131681745 N DEL 11
SRR1766480.4244510 chr11 131681024 N chr11 131681581 N DUP 14
SRR1766442.22272196 chr11 131680956 N chr11 131681431 N DEL 11
SRR1766472.5422475 chr11 131681127 N chr11 131681464 N DEL 13
SRR1766485.9659235 chr11 131680954 N chr11 131681449 N DEL 13
SRR1766475.10705296 chr11 131681127 N chr11 131681464 N DEL 13
SRR1766452.3067670 chr11 131681127 N chr11 131681464 N DEL 13
SRR1766443.7504084 chr11 131681691 N chr11 131681958 N DUP 13
SRR1766485.9168166 chr11 131681704 N chr11 131681881 N DEL 11
SRR1766482.4839095 chr11 131681398 N chr11 131681743 N DUP 10
SRR1766445.2478786 chr11 131681391 N chr11 131681478 N DEL 16
SRR1766480.4230284 chr11 131680951 N chr11 131681746 N DEL 14
SRR1766446.106277 chr11 131680971 N chr11 131681836 N DUP 11
SRR1766460.11013096 chr9 125780243 N chr9 125780420 N DEL 10
SRR1766457.6876832 chr9 125780243 N chr9 125780420 N DEL 15
SRR1766463.1836404 chr9 125780243 N chr9 125780420 N DEL 15
SRR1766466.8953459 chr9 125779983 N chr9 125780284 N DUP 15
SRR1766463.3716772 chr10 133121487 N chr10 133121775 N DUP 10
SRR1766462.10970962 chr20 62452080 N chr20 62452262 N DUP 10
SRR1766460.11014805 chr20 18022266 N chr20 18022702 N DEL 10
SRR1766479.9930182 chr20 18022337 N chr20 18022394 N DEL 10
SRR1766483.1002366 chr20 18022498 N chr20 18022859 N DEL 10
SRR1766444.7293689 chr20 18022169 N chr20 18022473 N DUP 11
SRR1766442.1739994 chr20 18022232 N chr20 18022610 N DEL 19
SRR1766458.8738183 chr20 18022224 N chr20 18022602 N DEL 19
SRR1766475.5806936 chr20 18022233 N chr20 18022611 N DEL 19
SRR1766452.2423012 chr20 18022166 N chr20 18022602 N DEL 17
SRR1766449.3501766 chr20 18022721 N chr20 18022836 N DEL 10
SRR1766473.2436685 chr20 18022230 N chr20 18022896 N DEL 10
SRR1766465.8939666 chr20 18022781 N chr20 18022897 N DEL 11
SRR1766457.4923504 chr20 18022213 N chr20 18023039 N DEL 10
SRR1766464.10273931 chr20 18022721 N chr20 18023068 N DEL 14
SRR1766473.10484335 chr20 18023340 N chr20 18023487 N DEL 13
SRR1766470.1795646 chr20 18022317 N chr20 18023334 N DEL 10
SRR1766442.34298947 chr6 9163024 N chr6 9163077 N DUP 10
SRR1766460.11236143 chr11 17764211 N chr11 17764341 N DUP 13
SRR1766468.742747 chrX 82073193 N chrX 82073286 N DEL 12
SRR1766479.13149448 chr19 16379964 N chr19 16380370 N DEL 10
SRR1766444.4134240 chr19 16379926 N chr19 16380036 N DEL 18
SRR1766460.7979433 chr19 16380399 N chr19 16380620 N DUP 10
SRR1766466.6781506 chr3 134701429 N chr3 134701482 N DUP 19
SRR1766462.793001 chr3 134701368 N chr3 134701427 N DEL 18
SRR1766482.12756642 chr3 134701446 N chr3 134701521 N DUP 14
SRR1766485.5117594 chr3 134701351 N chr3 134701552 N DUP 10
SRR1766448.2380883 chr3 134701351 N chr3 134701552 N DUP 10
SRR1766480.2346701 chr1 4939626 N chr1 4939729 N DUP 15
SRR1766481.2051429 chr1 4939626 N chr1 4939729 N DUP 14
SRR1766457.8085612 chr1 4939626 N chr1 4939729 N DUP 13
SRR1766460.878317 chr20 60500735 N chr20 60501080 N DEL 15
SRR1766460.8051837 chr20 60500396 N chr20 60500846 N DEL 10
SRR1766483.547354 chr20 60500395 N chr20 60501189 N DEL 10
SRR1766446.5126123 chr20 60500445 N chr20 60501452 N DEL 15
SRR1766446.5579418 chr20 60500426 N chr20 60501533 N DEL 14
SRR1766462.5804078 chr15 28105152 N chr15 28105998 N DEL 10
SRR1766447.8968805 chr3 88436022 N chr3 88436081 N DEL 14
