SRR1766466.1404632 chr7 57927474 N chr7 57927815 N DEL 44
SRR1766455.337821 chr10 36190353 N chr10 36190404 N DEL 52
SRR1766461.10304192 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766442.7404353 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766442.15088056 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766463.2954081 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766448.1187225 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766455.9479418 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766460.8068078 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766468.6580840 chr15 21776993 N chr15 21777343 N DEL 53
SRR1766457.2160821 chr8 121201731 N chr8 121201814 N DUP 43
SRR1766485.5863073 chr8 121201731 N chr8 121201814 N DUP 40
SRR1766454.9742568 chr8 121201731 N chr8 121201814 N DUP 43
SRR1766459.384090 chr8 121201731 N chr8 121201814 N DUP 40
SRR1766459.183775 chr8 121201731 N chr8 121201814 N DUP 40
SRR1766486.4938184 chr8 121201731 N chr8 121201814 N DUP 41
SRR1766458.1283414 chr8 121201731 N chr8 121201814 N DUP 43
SRR1766457.8514731 chr7 157994662 N chr7 157995435 N DEL 41
SRR1766468.1900450 chr5 40697200 N chr5 40697301 N DEL 50
SRR1766460.5875149 chr5 40697200 N chr5 40697301 N DEL 50
SRR1766474.2218712 chr18 22740454 N chr18 22740521 N DUP 46
SRR1766472.2340108 chr18 22740454 N chr18 22740521 N DUP 46
SRR1766467.9015539 chr18 22740454 N chr18 22740521 N DUP 46
SRR1766443.10189656 chr13 87990186 N chr13 87990243 N DEL 56
SRR1766469.7932559 chr13 87990186 N chr13 87990243 N DEL 57
SRR1766457.5232709 chr13 87990186 N chr13 87990243 N DEL 60
SRR1766463.7962679 chr13 87990186 N chr13 87990243 N DEL 53
SRR1766455.7092090 chr13 87990186 N chr13 87990243 N DEL 42
SRR1766445.812646 chr13 87990186 N chr13 87990243 N DEL 41
SRR1766442.46781775 chr4 117740001 N chr4 117740063 N DUP 41
SRR1766448.9274559 chr16 89342136 N chr16 89342227 N DEL 48
SRR1766477.4580543 chr16 89342136 N chr16 89342227 N DEL 44
SRR1766471.8788883 chr12 39712527 N chr12 39712642 N DEL 46
SRR1766446.2492785 chr10 92393323 N chr10 92393556 N DEL 42
SRR1766445.1971641 chr9 9845167 N chr9 9845230 N DEL 53
SRR1766468.6985064 chr9 135261811 N chr9 135261926 N DEL 53
SRR1766442.8095465 chr12 78626252 N chr12 78626307 N DUP 41
SRR1766442.12445560 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766450.3138475 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766472.1700060 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766442.8815642 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766445.9892531 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766462.8181061 chr16 73349787 N chr16 73349847 N DEL 40
SRR1766480.7124154 chr10 47500918 N chr10 47501079 N DEL 50
SRR1766445.7827924 chr4 180390615 N chr4 180391224 N DEL 42
SRR1766454.5424402 chr4 180390615 N chr4 180391224 N DEL 41
SRR1766442.25714311 chr6 162011471 N chr6 162011656 N DEL 51
SRR1766444.6190508 chr6 162011471 N chr6 162011656 N DEL 51
SRR1766482.136209 chr13 62019547 N chr13 62019606 N DEL 63
SRR1766468.6325797 chr8 140120705 N chr8 140120870 N DEL 41
SRR1766483.6629982 chr3 184414763 N chr3 184414888 N DEL 43
SRR1766476.10462932 chr13 27999196 N chr13 27999260 N DUP 42
SRR1766472.11328600 chr19 39153429 N chr19 39153611 N DUP 46
SRR1766444.4837942 chr7 132647014 N chr7 132647345 N DEL 55
SRR1766468.2074319 chr2 206104325 N chr2 206104473 N DEL 44
SRR1766486.9950591 chr7 40377351 N chr7 40377404 N DEL 46
SRR1766478.7707663 chr7 40377351 N chr7 40377404 N DEL 46
SRR1766458.9347111 chr7 40377326 N chr7 40377404 N DEL 42
SRR1766442.35734643 chr5 175050945 N chr5 175051029 N DUP 46
SRR1766445.504216 chr5 175050945 N chr5 175051029 N DUP 45
SRR1766455.553817 chr5 175050953 N chr5 175051008 N DUP 42
SRR1766463.148498 chr5 175050945 N chr5 175051029 N DUP 43
SRR1766471.6238285 chr5 175050945 N chr5 175051029 N DUP 40
SRR1766483.8909131 chr5 175050944 N chr5 175051028 N DUP 41
SRR1766463.602383 chr5 175050945 N chr5 175051029 N DUP 41
SRR1766466.2065916 chr5 175050945 N chr5 175051029 N DUP 45
SRR1766469.4497478 chr5 175050945 N chr5 175051029 N DUP 46
SRR1766471.6698630 chr5 175050945 N chr5 175051029 N DUP 46
SRR1766466.9559969 chr5 175050953 N chr5 175051008 N DUP 48
SRR1766465.10918318 chr5 175050945 N chr5 175051029 N DUP 47
SRR1766474.3466537 chr5 175050945 N chr5 175051029 N DUP 47
SRR1766461.2177190 chr5 175050945 N chr5 175051029 N DUP 48
SRR1766475.5285578 chr5 175050945 N chr5 175051029 N DUP 48
SRR1766484.7853826 chr5 175050944 N chr5 175051028 N DUP 48
SRR1766486.8999378 chr5 175050945 N chr5 175051029 N DUP 48
SRR1766474.3490832 chr5 175050953 N chr5 175051008 N DUP 48
SRR1766457.579844 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766457.9467093 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766466.11002212 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766461.3594756 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766476.2840754 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766482.5844 chr5 175050953 N chr5 175051008 N DUP 41
SRR1766463.4045534 chr2 57548108 N chr2 57548161 N DEL 51
SRR1766463.2018673 chr14 86443460 N chr14 86443552 N DUP 41
SRR1766442.21800567 chr14 86443460 N chr14 86443584 N DUP 45
SRR1766452.10667945 chr14 86443460 N chr14 86443584 N DUP 41
SRR1766474.2676307 chr14 86443460 N chr14 86443513 N DUP 48
SRR1766473.9157197 chr14 86443753 N chr14 86443833 N DUP 40
SRR1766473.5821116 chr14 86443753 N chr14 86443833 N DUP 40
SRR1766453.2768409 chr3 93470409 N chr3 93470458 N DUP 43
SRR1766443.9825298 chr7 112391885 N chr7 112392302 N DEL 65
SRR1766444.374611 chr1 152910560 N chr1 152910891 N DEL 45
SRR1766453.5121668 chr4 43451137 N chr4 43451231 N DEL 42
SRR1766466.2585089 chr4 43451137 N chr4 43451231 N DEL 46
SRR1766481.4666068 chr4 43451137 N chr4 43451231 N DEL 46
SRR1766444.5700040 chr6 169924033 N chr6 169924140 N DUP 46
SRR1766457.772081 chr5 162906168 N chr5 162906219 N DEL 42
SRR1766447.3101985 chr4 157544042 N chr4 157544095 N DEL 57
SRR1766456.861808 chr11 71362439 N chr11 71363109 N DUP 45
SRR1766442.28055915 chr1 24907838 N chr1 24908214 N DEL 46
SRR1766481.10385244 chr1 125179351 N chr1 125179404 N DEL 57
SRR1766442.2578512 chr18 2222995 N chr18 2223048 N DEL 57
SRR1766448.4489752 chr2 90383062 N chr2 90383135 N DEL 43
SRR1766477.5099405 chr2 90383062 N chr2 90383135 N DEL 40
SRR1766485.3592883 chr2 90383062 N chr2 90383135 N DEL 42
SRR1766471.6817426 chr2 90383062 N chr2 90383135 N DEL 40
SRR1766442.26017437 chr6 54310807 N chr6 54310873 N DEL 40
SRR1766484.5243983 chr6 54310807 N chr6 54310873 N DEL 43
SRR1766443.5192120 chr6 54310807 N chr6 54310873 N DEL 45
SRR1766442.17971201 chr6 54310807 N chr6 54310873 N DEL 46
SRR1766446.5989979 chr6 54310807 N chr6 54310873 N DEL 49
SRR1766467.6641138 chr10 57693565 N chr10 57693737 N DEL 41
SRR1766444.253104 chr17 2226520 N chr17 2226837 N DEL 43
SRR1766449.1972374 chr3 60861363 N chr3 60861418 N DUP 45
SRR1766454.867446 chr3 60861363 N chr3 60861418 N DUP 49
SRR1766442.31422660 chr3 60861363 N chr3 60861418 N DUP 50
SRR1766464.1820646 chr3 60861363 N chr3 60861418 N DUP 50
SRR1766476.518582 chr3 60861363 N chr3 60861418 N DUP 43
SRR1766447.3730770 chrX 35692492 N chrX 35692559 N DUP 41
SRR1766461.9713008 chrX 35692492 N chrX 35692559 N DUP 41
SRR1766460.3099710 chrX 35692492 N chrX 35692559 N DUP 40
SRR1766476.5571681 chr5 138143756 N chr5 138143823 N DEL 58
SRR1766461.4433608 chr10 2871852 N chr10 2871910 N DEL 49
SRR1766476.3675767 chr6 38103619 N chr6 38103674 N DEL 57
SRR1766484.7238743 chr6 38103619 N chr6 38103674 N DEL 43
SRR1766449.2476763 chr6 38103619 N chr6 38103674 N DEL 43
SRR1766459.2346732 chr6 38103619 N chr6 38103674 N DEL 46
SRR1766468.6325797 chr8 140120705 N chr8 140120870 N DEL 41
SRR1766486.3719446 chr3 134701427 N chr3 134701504 N DUP 41
SRR1766447.5094949 chr3 134701427 N chr3 134701504 N DUP 44
