SRR1766474.5265723 chrX 146812286 N chrX 146812377 N DEL 9
SRR1766474.68894 chrX 146812286 N chrX 146812377 N DEL 7
SRR1766449.1087981 chrX 146812304 N chrX 146812395 N DUP 7
SRR1766443.607980 chr6 161746956 N chr6 161747005 N DUP 5
SRR1766480.5833704 chr6 161746788 N chr6 161747013 N DUP 5
SRR1766442.13839240 chr6 40209132 N chr6 40209689 N DEL 5
SRR1766469.2711675 chr6 40209132 N chr6 40209689 N DEL 5
SRR1766477.3216402 chr6 40209132 N chr6 40209689 N DEL 5
SRR1766453.7868313 chr6 40209142 N chr6 40209887 N DEL 6
SRR1766483.6750295 chr6 40209142 N chr6 40209887 N DEL 7
SRR1766466.5890291 chr6 40209142 N chr6 40209647 N DEL 7
SRR1766454.8474156 chr6 40209142 N chr6 40209647 N DEL 9
SRR1766473.9568686 chr6 40209174 N chr6 40209625 N DEL 10
SRR1766462.670452 chr6 40209145 N chr6 40209198 N DUP 14
SRR1766473.4075371 chr6 40209145 N chr6 40209198 N DUP 14
SRR1766477.890951 chr6 40209145 N chr6 40209198 N DUP 14
SRR1766457.549986 chr6 40209145 N chr6 40209198 N DUP 14
SRR1766442.4751937 chr6 40209147 N chr6 40209234 N DUP 5
SRR1766472.5819937 chr6 40209147 N chr6 40209234 N DUP 6
SRR1766447.3435014 chr6 40209145 N chr6 40209198 N DUP 10
SRR1766446.7051739 chr6 40209154 N chr6 40209913 N DUP 18
SRR1766442.42445526 chr6 40209513 N chr6 40209764 N DUP 22
SRR1766469.1573710 chr6 40209513 N chr6 40209764 N DUP 22
SRR1766447.9882624 chr6 40209134 N chr6 40209197 N DUP 14
SRR1766457.4275394 chr6 40209138 N chr6 40209275 N DUP 11
SRR1766460.3882408 chr6 40209227 N chr6 40209914 N DUP 17
SRR1766456.5530273 chr6 40209275 N chr6 40209364 N DEL 17
SRR1766486.8209297 chr6 40209227 N chr6 40209606 N DUP 14
SRR1766457.4145131 chr6 40209161 N chr6 40209718 N DUP 10
SRR1766462.7242706 chr6 40209314 N chr6 40209409 N DEL 16
SRR1766469.2711675 chr6 40209267 N chr6 40209776 N DEL 21
SRR1766444.5330388 chr6 40209267 N chr6 40209812 N DEL 23
SRR1766472.1493340 chr6 40209267 N chr6 40209812 N DEL 23
SRR1766485.9634000 chr6 40209227 N chr6 40209606 N DUP 11
SRR1766450.2073233 chr6 40209343 N chr6 40209416 N DEL 23
SRR1766475.10669225 chr6 40209327 N chr6 40209528 N DEL 28
SRR1766478.7536017 chr6 40209309 N chr6 40209422 N DEL 13
SRR1766447.9326736 chr6 40209275 N chr6 40209364 N DEL 17
SRR1766463.815128 chr6 40209192 N chr6 40209273 N DEL 15
SRR1766449.5984102 chr6 40209267 N chr6 40209704 N DEL 22
SRR1766464.7652180 chr6 40209267 N chr6 40209704 N DEL 22
SRR1766442.26017208 chr6 40209267 N chr6 40209740 N DEL 24
SRR1766472.4368075 chr6 40209267 N chr6 40209740 N DEL 24
SRR1766454.1184692 chr6 40209226 N chr6 40209693 N DEL 11
SRR1766453.3507462 chr6 40209389 N chr6 40209866 N DEL 19
SRR1766459.619374 chr6 40209389 N chr6 40209812 N DEL 21
SRR1766466.2830877 chr6 40209389 N chr6 40209812 N DEL 21
SRR1766473.7390458 chr6 40209309 N chr6 40209422 N DEL 20
SRR1766462.2079898 chr6 40209327 N chr6 40209792 N DEL 29
SRR1766455.914097 chr6 40209327 N chr6 40209792 N DEL 28
SRR1766478.7660085 chr6 40209309 N chr6 40209422 N DEL 20
SRR1766464.6163263 chr6 40209693 N chr6 40209762 N DUP 5
SRR1766472.8450164 chr6 40209322 N chr6 40209805 N DEL 23
SRR1766460.7211391 chr6 40209322 N chr6 40209805 N DEL 24
SRR1766451.1403969 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766481.6328673 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766477.7553933 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766442.33120376 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766450.3168715 chr6 40209322 N chr6 40209805 N DEL 29
SRR1766445.9878414 chr6 40209470 N chr6 40209805 N DEL 25
SRR1766457.3977199 chr6 40209292 N chr6 40209805 N DEL 36
SRR1766462.2718922 chr6 40209297 N chr6 40209792 N DEL 31
SRR1766456.4428090 chr6 40209509 N chr6 40209570 N DUP 7
SRR1766453.1306798 chr6 40209557 N chr6 40209782 N DUP 17
SRR1766479.11915969 chr6 40209557 N chr6 40209782 N DUP 17
SRR1766469.6318633 chr6 40209535 N chr6 40209850 N DUP 21
SRR1766485.4396315 chr6 40209471 N chr6 40209550 N DUP 9
SRR1766482.13049617 chr6 40209435 N chr6 40209568 N DUP 11
SRR1766462.670452 chr6 40209327 N chr6 40209528 N DEL 24
SRR1766486.9317420 chr6 40209219 N chr6 40209446 N DUP 7
SRR1766447.9305880 chr6 40209172 N chr6 40209646 N DEL 14
SRR1766446.10490628 chr6 40209435 N chr6 40209642 N DEL 9
SRR1766446.6025057 chr6 40209597 N chr6 40209828 N DEL 23
SRR1766447.8376972 chr6 40209597 N chr6 40209828 N DEL 21
SRR1766485.5998535 chr6 40209605 N chr6 40209864 N DEL 31
SRR1766482.12819399 chr6 40209605 N chr6 40209864 N DEL 28
SRR1766455.1378690 chr6 40209699 N chr6 40209910 N DUP 17
SRR1766468.5053632 chr6 40209605 N chr6 40209864 N DEL 22
SRR1766455.7600844 chr6 40209710 N chr6 40209933 N DUP 17
SRR1766461.225301 chr6 40209766 N chr6 40209863 N DUP 19
SRR1766473.9568686 chr6 40209766 N chr6 40209863 N DUP 19
SRR1766454.7893747 chr6 40209767 N chr6 40209864 N DUP 17
SRR1766454.2849246 chr6 40209810 N chr6 40209905 N DUP 12
SRR1766460.7018530 chr6 40209521 N chr6 40209914 N DUP 17
SRR1766482.5377961 chr6 40209566 N chr6 40209751 N DEL 16
SRR1766457.8845115 chr6 40209789 N chr6 40209910 N DUP 28
SRR1766471.5915735 chr6 40209710 N chr6 40209933 N DUP 27
SRR1766447.4273536 chr6 40209710 N chr6 40209933 N DUP 28
SRR1766466.1461148 chr6 40209513 N chr6 40209900 N DUP 14
SRR1766455.7104459 chr6 40209476 N chr6 40209871 N DUP 7
SRR1766448.7464201 chr6 40209594 N chr6 40209789 N DEL 22
SRR1766444.1954797 chr6 40209576 N chr6 40209771 N DEL 26
SRR1766443.8549389 chr6 40209602 N chr6 40209789 N DEL 25
SRR1766450.6976269 chr6 40209710 N chr6 40209933 N DUP 35
SRR1766454.7416014 chr6 40209710 N chr6 40209933 N DUP 33
SRR1766442.38069493 chr6 40209710 N chr6 40209933 N DUP 32
SRR1766451.3569801 chr6 40209440 N chr6 40209555 N DUP 17
SRR1766474.4657954 chr6 40209710 N chr6 40209933 N DUP 29
SRR1766476.4536931 chr6 40209710 N chr6 40209933 N DUP 28
SRR1766470.642355 chr6 40209792 N chr6 40209845 N DUP 3
SRR1766450.929104 chr6 40209792 N chr6 40209845 N DUP 4
SRR1766481.7621377 chr6 40209792 N chr6 40209845 N DUP 5
SRR1766461.10258966 chr6 40209699 N chr6 40209910 N DUP 22
SRR1766462.11185331 chr6 40209446 N chr6 40209799 N DEL 24
SRR1766453.1324498 chr6 40209446 N chr6 40209799 N DEL 24
SRR1766443.5327830 chr6 40209446 N chr6 40209799 N DEL 23
SRR1766443.2709190 chr6 40209581 N chr6 40209792 N DEL 27
SRR1766467.10408201 chr6 40209439 N chr6 40209792 N DEL 23
SRR1766449.601789 chr6 40209545 N chr6 40209792 N DEL 10
SRR1766482.5377961 chr6 40209297 N chr6 40209792 N DEL 25
SRR1766451.3864695 chr6 40209512 N chr6 40209899 N DUP 11
SRR1766476.2995335 chr6 40209512 N chr6 40209899 N DUP 11
SRR1766485.2258795 chr6 40209679 N chr6 40209884 N DUP 9
SRR1766472.10092431 chr6 40209486 N chr6 40209883 N DUP 17
SRR1766467.2602274 chr6 40209520 N chr6 40209921 N DUP 11
SRR1766484.202117 chr6 40209545 N chr6 40209792 N DEL 10
SRR1766486.4930575 chr6 40209164 N chr6 40209713 N DEL 1
SRR1766442.26986129 chr6 40209710 N chr6 40209933 N DUP 31
SRR1766442.25191808 chr6 40209521 N chr6 40209914 N DUP 17
SRR1766467.3039022 chr6 40209434 N chr6 40209805 N DEL 9
SRR1766444.2847076 chr6 40209789 N chr6 40209910 N DUP 27
SRR1766447.7717411 chr6 40209436 N chr6 40209927 N DUP 4
SRR1766469.2973266 chr6 40209561 N chr6 40209810 N DEL 9
SRR1766445.4999125 chr6 40209512 N chr6 40209899 N DUP 16
SRR1766442.27163626 chr6 40209563 N chr6 40209800 N DEL 22
SRR1766463.2468135 chr6 40209605 N chr6 40209864 N DEL 28
SRR1766458.1050790 chr6 40209513 N chr6 40209900 N DUP 12
SRR1766484.3925706 chr6 40209513 N chr6 40209900 N DUP 13
SRR1766442.12541431 chr6 40209810 N chr6 40209913 N DUP 19
SRR1766473.6636659 chr6 40209605 N chr6 40209864 N DEL 18
SRR1766450.8524 chr6 40209605 N chr6 40209864 N DEL 18
SRR1766442.20536606 chr6 40209605 N chr6 40209864 N DEL 17
SRR1766471.2270222 chr6 40209161 N chr6 40209864 N DEL 14
SRR1766442.27668881 chr6 40209535 N chr6 40209864 N DEL 12
SRR1766443.296974 chr6 40209787 N chr6 40209912 N DEL 13
SRR1766473.9221763 chr6 40209554 N chr6 40209889 N DEL 11
SRR1766476.9406087 chr6 40209554 N chr6 40209889 N DEL 9
SRR1766442.37302361 chr6 40209744 N chr6 40209903 N DEL 19
SRR1766460.3882408 chr6 40209744 N chr6 40209903 N DEL 18
SRR1766455.1329637 chr6 40209744 N chr6 40209903 N DEL 18
SRR1766475.10669225 chr6 40209765 N chr6 40209908 N DEL 16
SRR1766442.26017208 chr6 40209744 N chr6 40209903 N DEL 18
SRR1766473.680692 chr6 40209744 N chr6 40209903 N DEL 18
SRR1766470.8625940 chr6 40209491 N chr6 40209896 N DEL 14
SRR1766444.2979777 chr6 40209154 N chr6 40209913 N DEL 18
SRR1766482.2261671 chr6 40209154 N chr6 40209913 N DEL 18
SRR1766467.5781574 chr6 40209144 N chr6 40209913 N DEL 15
SRR1766442.21006621 chr6 40209144 N chr6 40209913 N DEL 12
SRR1766442.45028464 chr6 40209144 N chr6 40209915 N DEL 3
SRR1766486.6464121 chr6 40209147 N chr6 40209916 N DEL 9
SRR1766449.1627369 chr6 40209153 N chr6 40209922 N DEL 6
SRR1766457.4582181 chr10 1409649 N chr10 1409734 N DEL 5
SRR1766453.4064964 chr10 1409628 N chr10 1409861 N DUP 5
SRR1766453.537775 chr10 1409618 N chr10 1409851 N DUP 5
SRR1766454.1072266 chr10 1409628 N chr10 1409861 N DUP 10
SRR1766473.9695147 chr10 1409618 N chr10 1409935 N DUP 2
SRR1766474.518223 chr10 1409618 N chr10 1409935 N DUP 7
SRR1766484.1873160 chr10 1409637 N chr10 1409954 N DUP 5
SRR1766482.6415157 chr10 1409638 N chr10 1409955 N DUP 5
SRR1766480.2458580 chr7 57927384 N chr7 57928234 N DUP 14
SRR1766484.4095234 chr7 57927506 N chr7 57927676 N DEL 3
SRR1766467.5869904 chr7 57927523 N chr7 57928204 N DEL 3
SRR1766466.1404632 chr7 57927474 N chr7 57927815 N DEL 44
SRR1766469.4500409 chr7 57927287 N chr7 57927968 N DEL 9
SRR1766443.2053383 chr7 57927344 N chr7 57928025 N DEL 8
SRR1766485.3726830 chr7 57928293 N chr7 57928807 N DEL 17
SRR1766473.11750216 chr7 57928532 N chr7 57928704 N DEL 5
SRR1766482.11358115 chr7 57927963 N chr7 57928474 N DEL 8
SRR1766448.11045315 chr7 57928109 N chr7 57928618 N DUP 7
SRR1766442.35470626 chr7 57927759 N chr7 57928608 N DUP 2
SRR1766472.10424680 chr7 57927521 N chr7 57928541 N DEL 11
SRR1766458.1129689 chr7 57927457 N chr7 57928646 N DUP 13
SRR1766444.6967693 chr7 57928565 N chr7 57928735 N DUP 1
SRR1766454.9642876 chr7 57928584 N chr7 57928756 N DEL 15
SRR1766461.10244698 chr7 57928741 N chr7 57928913 N DEL 13
SRR1766444.5162074 chr2 10015464 N chr2 10015521 N DUP 5
SRR1766448.3577138 chr2 10015482 N chr2 10015812 N DUP 2
SRR1766486.11951114 chr2 10015504 N chr2 10016131 N DUP 5
SRR1766443.5158616 chr2 10015574 N chr2 10015631 N DUP 10
SRR1766442.3545447 chr2 10015535 N chr2 10016022 N DUP 6
SRR1766462.4603369 chr2 10015918 N chr2 10016004 N DUP 34
SRR1766471.380841 chr2 10015572 N chr2 10016199 N DUP 5
SRR1766476.5927099 chr2 10015563 N chr2 10015622 N DEL 5
SRR1766445.7480971 chr2 10015566 N chr2 10015681 N DUP 5
SRR1766468.5914649 chr2 10015615 N chr2 10016015 N DUP 5
SRR1766442.39674558 chr2 10015560 N chr2 10015648 N DEL 10
SRR1766482.2468977 chr2 10015560 N chr2 10015648 N DEL 5
SRR1766462.3249282 chr2 10015519 N chr2 10015665 N DEL 5
SRR1766482.10143995 chr2 10015689 N chr2 10016171 N DUP 2
SRR1766453.1367953 chr2 10015493 N chr2 10015697 N DEL 2
SRR1766442.22180632 chr2 10015549 N chr2 10015724 N DEL 10
SRR1766444.5811458 chr2 10015461 N chr2 10015820 N DUP 14
SRR1766453.2312095 chr2 10015549 N chr2 10015724 N DEL 10
SRR1766461.7945951 chr2 10015650 N chr2 10015767 N DEL 2
SRR1766482.3981777 chr2 10015503 N chr2 10015874 N DUP 10
SRR1766445.6450227 chr2 10015479 N chr2 10015770 N DEL 5
SRR1766461.3630218 chr2 10015560 N chr2 10015834 N DEL 10
SRR1766455.6460420 chr2 10015856 N chr2 10016256 N DUP 10
SRR1766463.10068212 chr2 10015695 N chr2 10015865 N DEL 5
SRR1766442.6929645 chr2 10015632 N chr2 10015918 N DEL 20
SRR1766447.5536306 chr2 10015522 N chr2 10015866 N DEL 5
SRR1766450.387849 chr2 10015545 N chr2 10015889 N DEL 12
SRR1766472.2917252 chr2 10015538 N chr2 10015911 N DEL 10
SRR1766483.12509417 chr2 10015665 N chr2 10015893 N DEL 11
SRR1766461.5928700 chr2 10015545 N chr2 10015918 N DEL 32
SRR1766448.3180146 chr2 10015562 N chr2 10015935 N DEL 10
SRR1766450.7506182 chr2 10015632 N chr2 10015918 N DEL 18
SRR1766461.10190401 chr2 10015480 N chr2 10015940 N DEL 12
SRR1766443.799642 chr2 10015544 N chr2 10015975 N DEL 1
SRR1766469.1792511 chr2 10015570 N chr2 10016139 N DUP 5
SRR1766448.41819 chr2 10015585 N chr2 10016127 N DEL 5
SRR1766442.25280663 chr2 10016168 N chr2 10016225 N DUP 1
SRR1766446.162094 chr2 10015475 N chr2 10016191 N DEL 5
SRR1766454.6729304 chr2 10015488 N chr2 10016262 N DEL 5
SRR1766444.5811458 chr2 10016098 N chr2 10016354 N DEL 22
SRR1766484.4623757 chr5 92251214 N chr5 92251265 N DUP 13
SRR1766442.10696079 chr5 92251214 N chr5 92251265 N DUP 13
SRR1766485.4612852 chr5 92251214 N chr5 92251265 N DUP 13
SRR1766449.1832322 chr5 92251215 N chr5 92251326 N DUP 21
SRR1766467.1739391 chr5 92251231 N chr5 92251312 N DEL 8
SRR1766442.36759277 chr5 92251454 N chr5 92251513 N DUP 12
SRR1766482.6350970 chr5 92251454 N chr5 92251513 N DUP 13
SRR1766450.10885329 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766484.8893486 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766447.9303687 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766477.6271903 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766476.4404715 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766472.6831349 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766470.6645822 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766443.2272923 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766471.11106732 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766475.9824406 chr5 92251454 N chr5 92251513 N DUP 18
SRR1766461.7556522 chr5 92251207 N chr5 92251454 N DEL 9
SRR1766481.9077045 chr5 92251211 N chr5 92251458 N DEL 9
SRR1766459.7837757 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766473.6477462 chr5 92251502 N chr5 92251635 N DUP 7
SRR1766454.5150949 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766442.39144130 chr5 92251472 N chr5 92251567 N DUP 11
SRR1766481.7325313 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766476.166040 chr5 92251472 N chr5 92251567 N DUP 11
SRR1766447.4120250 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766484.2954826 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766479.9735463 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766477.9224121 chr5 92251472 N chr5 92251601 N DUP 11
SRR1766471.3081370 chr5 92251472 N chr5 92251567 N DUP 11
SRR1766442.15349372 chr5 92251472 N chr5 92251533 N DUP 11
SRR1766482.8105708 chr5 92251477 N chr5 92251576 N DEL 1
SRR1766443.5229751 chr10 36190353 N chr10 36190404 N DEL 9
SRR1766458.8518665 chr10 36190353 N chr10 36190404 N DEL 11
SRR1766455.337821 chr10 36190353 N chr10 36190404 N DEL 52
SRR1766461.10304192 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766442.7404353 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766442.15088056 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766463.2954081 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766448.1187225 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766455.9479418 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766460.8068078 chr10 36190353 N chr10 36190404 N DEL 55
SRR1766470.8866232 chr10 36190358 N chr10 36190409 N DEL 10
SRR1766476.7031268 chr15 21777101 N chr15 21777450 N DEL 5
SRR1766472.9719126 chr15 21777066 N chr15 21777415 N DEL 5
SRR1766451.4329725 chr15 21777066 N chr15 21777415 N DEL 25
SRR1766458.9133773 chr15 21777133 N chr15 21777482 N DEL 10
SRR1766464.10702561 chr15 21777136 N chr15 21777485 N DEL 15
SRR1766451.9012934 chr15 21777254 N chr15 21777605 N DEL 1
SRR1766468.6580840 chr15 21776993 N chr15 21777343 N DEL 53
SRR1766473.10090113 chr15 21777161 N chr15 21777510 N DEL 5
SRR1766481.5992998 chr17 81432869 N chr17 81432992 N DEL 8
SRR1766482.9682475 chr2 208177113 N chr2 208177164 N DEL 27
SRR1766461.1182085 chr2 208177089 N chr2 208177164 N DEL 19
SRR1766469.7791650 chr2 208177089 N chr2 208177164 N DEL 21
SRR1766472.3314723 chr2 208177089 N chr2 208177164 N DEL 19
SRR1766477.8871954 chr4 5842753 N chr4 5842834 N DEL 7
SRR1766444.4229060 chr19 40349878 N chr19 40350181 N DEL 8
SRR1766473.7750635 chr19 40349984 N chr19 40350287 N DEL 6
SRR1766443.212780 chr19 40350033 N chr19 40350336 N DEL 15
SRR1766467.4685206 chr19 40349851 N chr19 40350154 N DEL 5
SRR1766476.1051098 chr19 40349859 N chr19 40350162 N DEL 1
SRR1766484.2812032 chr19 40349896 N chr19 40350199 N DEL 10
SRR1766460.2912233 chr19 40349941 N chr19 40350244 N DEL 5
SRR1766462.5698135 chr19 40350057 N chr19 40350358 N DUP 3
SRR1766442.2128103 chr19 40349976 N chr19 40350279 N DEL 20
SRR1766442.17693725 chr19 40349973 N chr19 40350276 N DEL 10
SRR1766473.7750635 chr19 40349984 N chr19 40350287 N DEL 19
SRR1766461.9059112 chr4 95191954 N chr4 95192079 N DEL 3
SRR1766484.11270634 chr4 95192117 N chr4 95192452 N DUP 2
SRR1766445.7894087 chr4 95192460 N chr4 95192556 N DEL 10
SRR1766469.552333 chr4 95192523 N chr4 95192684 N DUP 5
SRR1766481.10261924 chr2 129895076 N chr2 129895281 N DEL 1
SRR1766442.41231614 chr2 129895151 N chr2 129895325 N DUP 5
SRR1766455.636635 chr2 129895049 N chr2 129895324 N DEL 5
SRR1766471.6046448 chr19 36796431 N chr19 36796482 N DEL 11
SRR1766456.1922052 chr9 65398366 N chr9 65398565 N DEL 12
SRR1766457.6043521 chr2 216226166 N chr2 216226736 N DUP 5
SRR1766442.17666671 chr2 216226366 N chr2 216226541 N DUP 5
SRR1766442.1556793 chr2 216226436 N chr2 216226632 N DUP 3
SRR1766475.8026983 chr2 216226465 N chr2 216226563 N DUP 12
SRR1766481.2976672 chr2 216226492 N chr2 216226541 N DUP 2
SRR1766480.6672806 chr2 216226480 N chr2 216226578 N DUP 5
SRR1766453.8194295 chr2 216226136 N chr2 216226488 N DEL 5
SRR1766469.6259942 chr2 216226332 N chr2 216226559 N DEL 5
SRR1766460.1221891 chr2 216226573 N chr2 216226742 N DUP 8
SRR1766477.231572 chr2 216226162 N chr2 216226689 N DUP 1
SRR1766459.122153 chr2 216226162 N chr2 216226689 N DUP 2
SRR1766481.1869062 chr2 216226288 N chr2 216226689 N DUP 8
SRR1766444.728493 chrX 21731630 N chrX 21731720 N DEL 16
SRR1766479.6363057 chrX 21731583 N chrX 21731636 N DUP 2
SRR1766443.3870587 chrX 21731583 N chrX 21731636 N DUP 2
SRR1766477.3338487 chrX 21731583 N chrX 21731636 N DUP 4
SRR1766475.2277589 chrX 21731583 N chrX 21731663 N DUP 2
SRR1766480.7780946 chrX 21731615 N chrX 21731670 N DEL 4
SRR1766452.9674882 chrX 21731713 N chrX 21731848 N DUP 5
SRR1766461.2215129 chrX 21731713 N chrX 21731848 N DUP 6
SRR1766477.1686589 chrX 21731713 N chrX 21731848 N DUP 8
SRR1766442.8330757 chrX 21731713 N chrX 21731848 N DUP 11
SRR1766479.957156 chrX 21731713 N chrX 21731848 N DUP 14
SRR1766446.6764419 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766472.4613969 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766458.3116698 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766466.1567353 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766476.854244 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766453.110206 chrX 21731713 N chrX 21731848 N DUP 21
SRR1766466.1548001 chrX 21731730 N chrX 21731859 N DEL 5
SRR1766478.3694025 chrX 21731762 N chrX 21731855 N DEL 9
SRR1766478.4823949 chr9 43335788 N chr9 43335865 N DUP 6
SRR1766481.4382009 chr9 43335699 N chr9 43335824 N DEL 15
SRR1766475.7535635 chr9 43335699 N chr9 43335824 N DEL 15
SRR1766486.1965635 chr9 43335699 N chr9 43335824 N DEL 15
SRR1766466.1359692 chr9 43335699 N chr9 43335902 N DEL 5
SRR1766470.1585931 chr9 43335703 N chr9 43335906 N DEL 5
SRR1766461.7813620 chr9 43335703 N chr9 43335906 N DEL 5
SRR1766443.4410980 chr8 82371371 N chr8 82371445 N DUP 1
SRR1766460.2664958 chr8 82371371 N chr8 82371445 N DUP 2
SRR1766468.7577578 chr3 111167155 N chr3 111167254 N DEL 24
SRR1766483.1620268 chr8 121201478 N chr8 121201629 N DEL 7
SRR1766473.9949580 chr8 121201478 N chr8 121201629 N DEL 7
SRR1766458.8963091 chr8 121201478 N chr8 121201629 N DEL 7
SRR1766451.1209638 chr8 121201478 N chr8 121201629 N DEL 7
SRR1766470.10134647 chr8 121201380 N chr8 121201459 N DUP 10
SRR1766456.643668 chr8 121201378 N chr8 121201457 N DUP 15
SRR1766442.42071246 chr8 121201360 N chr8 121201425 N DEL 5
SRR1766474.4601276 chr8 121201426 N chr8 121201769 N DUP 4
SRR1766472.5290621 chr8 121201652 N chr8 121201729 N DEL 4
SRR1766448.8348723 chr8 121201479 N chr8 121201666 N DUP 10
SRR1766443.1768199 chr8 121201535 N chr8 121201722 N DUP 1
SRR1766442.5720328 chr8 121201531 N chr8 121201644 N DEL 4
SRR1766453.10457893 chr8 121201534 N chr8 121201647 N DEL 1
SRR1766448.514375 chr8 121201495 N chr8 121201720 N DEL 2
SRR1766453.7906072 chr8 121201742 N chr8 121201797 N DUP 27
SRR1766466.5978198 chr8 121201742 N chr8 121201797 N DUP 31
SRR1766457.2160821 chr8 121201731 N chr8 121201814 N DUP 43
SRR1766461.9745147 chr8 121201743 N chr8 121201798 N DUP 36
SRR1766473.10430545 chr8 121201731 N chr8 121201814 N DUP 37
SRR1766482.12682478 chr8 121201731 N chr8 121201814 N DUP 37
SRR1766442.30384333 chr8 121201731 N chr8 121201814 N DUP 36
SRR1766472.4290844 chr8 121201742 N chr8 121201797 N DUP 36
SRR1766479.7782704 chr8 121201731 N chr8 121201814 N DUP 38
SRR1766485.5863073 chr8 121201731 N chr8 121201814 N DUP 40
SRR1766454.9742568 chr8 121201731 N chr8 121201814 N DUP 43
SRR1766459.384090 chr8 121201731 N chr8 121201814 N DUP 40
SRR1766476.1120260 chr8 121201731 N chr8 121201814 N DUP 36
SRR1766442.10320318 chr8 121201731 N chr8 121201814 N DUP 36
SRR1766479.12075917 chr8 121201731 N chr8 121201814 N DUP 36
SRR1766484.3570631 chr8 121201742 N chr8 121201797 N DUP 23
SRR1766445.6162180 chr8 121201760 N chr8 121201851 N DUP 21
SRR1766442.32155005 chr8 121201742 N chr8 121201797 N DUP 23
SRR1766451.288703 chr8 121201731 N chr8 121201814 N DUP 34
SRR1766454.3139006 chr8 121201731 N chr8 121201814 N DUP 34
SRR1766459.183775 chr8 121201731 N chr8 121201814 N DUP 40
SRR1766486.4938184 chr8 121201731 N chr8 121201814 N DUP 41
SRR1766464.1264448 chr8 121201742 N chr8 121201797 N DUP 36
SRR1766458.1283414 chr8 121201731 N chr8 121201814 N DUP 43
SRR1766444.450563 chr8 121201916 N chr8 121201977 N DEL 5
SRR1766474.2896056 chr8 121201769 N chr8 121201834 N DEL 18
SRR1766479.3003673 chr8 121201769 N chr8 121201834 N DEL 15
SRR1766460.3454021 chr8 121201770 N chr8 121201835 N DEL 14
SRR1766469.10075970 chr8 121201777 N chr8 121201842 N DEL 7
SRR1766453.7944451 chr8 121201770 N chr8 121201835 N DEL 14
SRR1766480.96935 chr8 121201775 N chr8 121201840 N DEL 9
SRR1766482.1825687 chr8 121201776 N chr8 121201841 N DEL 8
SRR1766459.390752 chr2 205380379 N chr2 205380509 N DEL 6
SRR1766478.80759 chr2 205380379 N chr2 205380509 N DEL 9
SRR1766463.3220717 chr2 205380379 N chr2 205380509 N DEL 9
SRR1766472.1960259 chr2 205380379 N chr2 205380509 N DEL 9
SRR1766442.14458877 chr2 205380379 N chr2 205380509 N DEL 9
SRR1766453.5941322 chr2 205380379 N chr2 205380509 N DEL 9
SRR1766472.9535453 chr2 205380379 N chr2 205380509 N DEL 9
SRR1766442.21275634 chr2 205380379 N chr2 205380612 N DEL 13
SRR1766470.1516395 chr2 205380379 N chr2 205380612 N DEL 13
SRR1766464.9212812 chr2 205380379 N chr2 205380612 N DEL 17
SRR1766474.8397851 chr2 205380379 N chr2 205380612 N DEL 18
SRR1766474.10150232 chr2 205380461 N chr2 205381219 N DEL 5
SRR1766444.6049303 chr2 205380379 N chr2 205380612 N DEL 18
SRR1766453.9676631 chr2 205380305 N chr2 205380501 N DEL 9
SRR1766451.2545851 chr2 205380454 N chr2 205380633 N DUP 7
SRR1766483.5358359 chr2 205380533 N chr2 205380633 N DUP 12
SRR1766484.6104771 chr2 205380453 N chr2 205380688 N DUP 8
SRR1766442.37992016 chr2 205380411 N chr2 205380619 N DEL 7
SRR1766446.8883970 chr2 205380406 N chr2 205380612 N DEL 2
SRR1766448.3783836 chr2 205380387 N chr2 205380751 N DUP 10
SRR1766451.9007298 chr2 205380453 N chr2 205380661 N DUP 7
SRR1766462.1118952 chr2 205380619 N chr2 205380697 N DUP 9
SRR1766479.611816 chr2 205380453 N chr2 205380688 N DUP 9
SRR1766465.2096849 chr2 205380489 N chr2 205380622 N DEL 15
SRR1766474.4326775 chr2 205380379 N chr2 205380612 N DEL 17
SRR1766484.291650 chr2 205380384 N chr2 205380617 N DEL 10
SRR1766479.4309612 chr2 205380453 N chr2 205380531 N DUP 7
SRR1766455.9590767 chr2 205380548 N chr2 205380600 N DEL 7
SRR1766471.4982973 chr2 205380453 N chr2 205380688 N DUP 7
SRR1766472.3022630 chr2 205380379 N chr2 205380612 N DEL 17
SRR1766460.6134476 chr2 205380496 N chr2 205380600 N DEL 7
SRR1766466.170331 chr2 205380453 N chr2 205380558 N DUP 7
SRR1766453.4539720 chr2 205380343 N chr2 205380599 N DEL 1
SRR1766467.2110545 chr2 205380343 N chr2 205380599 N DEL 1
SRR1766484.10565014 chr2 205380419 N chr2 205380600 N DEL 7
SRR1766470.4027341 chr2 205380453 N chr2 205380688 N DUP 7
SRR1766463.10809476 chr2 205380453 N chr2 205380715 N DUP 5
SRR1766466.7675469 chr2 205380453 N chr2 205380715 N DUP 8
SRR1766469.5152683 chr2 205380453 N chr2 205380688 N DUP 10
SRR1766460.5693910 chr2 205381058 N chr2 205381115 N DEL 9
SRR1766457.1764423 chr2 205381058 N chr2 205381115 N DEL 12
SRR1766471.4466941 chr2 205380388 N chr2 205381064 N DUP 14
SRR1766459.1387881 chr2 205380418 N chr2 205381046 N DEL 15
SRR1766455.7206234 chr2 205380406 N chr2 205381059 N DEL 2
SRR1766453.8585299 chr2 205380299 N chr2 205381296 N DEL 7
SRR1766447.9707278 chr2 205380503 N chr2 205381303 N DEL 7
SRR1766463.4679538 chr2 205380503 N chr2 205381303 N DEL 7
SRR1766454.7246248 chrX 899611 N chrX 899673 N DUP 2
SRR1766485.9084489 chrX 899434 N chrX 899696 N DEL 5
SRR1766476.1303951 chr16 1067918 N chr16 1067994 N DUP 3
SRR1766461.3065168 chr2 201283099 N chr2 201283548 N DEL 12
SRR1766465.11167067 chr2 201283147 N chr2 201283841 N DEL 5
SRR1766452.6971304 chr2 201283091 N chr2 201283539 N DUP 5
SRR1766452.6232413 chr2 201283115 N chr2 201283262 N DUP 5
SRR1766486.7962145 chr2 201283139 N chr2 201283188 N DUP 7
SRR1766484.8460363 chr2 201283100 N chr2 201283198 N DUP 5
SRR1766452.7383575 chr2 201283199 N chr2 201283373 N DUP 5
SRR1766470.2244457 chr2 201283502 N chr2 201283678 N DEL 5
SRR1766465.5738202 chr2 201283241 N chr2 201283417 N DEL 3
SRR1766479.878678 chr2 201283422 N chr2 201283598 N DEL 5
SRR1766453.3676431 chr2 201283502 N chr2 201283678 N DEL 6
SRR1766458.8789487 chr2 201283099 N chr2 201283548 N DEL 12
SRR1766482.12502555 chr2 201283555 N chr2 201283729 N DUP 5
SRR1766479.6378661 chr2 201283099 N chr2 201283548 N DEL 12
SRR1766459.7854680 chr2 201283270 N chr2 201283618 N DUP 5
SRR1766479.4487844 chr2 201283124 N chr2 201283525 N DEL 1
SRR1766461.3065168 chr2 201283100 N chr2 201283549 N DEL 11
SRR1766481.1235923 chr2 201283148 N chr2 201283596 N DEL 7
SRR1766449.6084280 chr2 201283081 N chr2 201283579 N DEL 5
SRR1766452.7658996 chr2 201283208 N chr2 201283683 N DUP 5
SRR1766455.6700331 chr2 201283198 N chr2 201283725 N DUP 2
SRR1766469.1270350 chr2 201283722 N chr2 201283842 N DEL 1
SRR1766485.9133509 chr2 201283053 N chr2 201283678 N DEL 5
SRR1766471.9960290 chr2 201283066 N chr2 201283691 N DEL 5
SRR1766454.1719378 chr2 201283193 N chr2 201283768 N DEL 4
SRR1766474.8011988 chr7 157994667 N chr7 157995319 N DEL 6
SRR1766457.8514731 chr7 157994662 N chr7 157995435 N DEL 41
SRR1766463.1769967 chr7 157994701 N chr7 157994819 N DEL 29
SRR1766481.5622972 chr7 157994701 N chr7 157994819 N DEL 30
SRR1766463.10420251 chr7 157994701 N chr7 157994819 N DEL 30
SRR1766459.8791744 chr7 157994652 N chr7 157994733 N DUP 9
SRR1766468.1303758 chr7 157994657 N chr7 157994738 N DUP 24
SRR1766475.7774262 chr7 157994720 N chr7 157995450 N DUP 12
SRR1766442.35192898 chr7 157994652 N chr7 157994733 N DUP 25
SRR1766462.881771 chr7 157994652 N chr7 157994733 N DUP 32
SRR1766478.1854747 chr7 157994652 N chr7 157994733 N DUP 24
SRR1766477.517048 chr7 157994647 N chr7 157994809 N DUP 6
SRR1766442.45589070 chr7 157994720 N chr7 157995450 N DUP 6
SRR1766460.4180092 chr7 157994717 N chr7 157995447 N DUP 9
SRR1766454.6011466 chr7 157994771 N chr7 157994852 N DUP 18
SRR1766464.5066659 chr7 157994771 N chr7 157994852 N DUP 20
SRR1766483.9778397 chr7 157994771 N chr7 157994852 N DUP 25
SRR1766462.1996092 chr7 157994867 N chr7 157995235 N DEL 10
SRR1766468.6902912 chr7 157994720 N chr7 157994802 N DEL 4
SRR1766479.7647386 chr7 157994706 N chr7 157994908 N DUP 5
SRR1766458.626563 chr7 157994701 N chr7 157994819 N DEL 30
SRR1766442.11428825 chr7 157994833 N chr7 157995441 N DUP 5
SRR1766468.143507 chr7 157994953 N chr7 157995401 N DEL 5
SRR1766462.1921776 chr7 157994819 N chr7 157994939 N DUP 5
SRR1766453.10766090 chr7 157994806 N chr7 157995129 N DUP 5
SRR1766452.6302503 chr7 157994706 N chr7 157994908 N DUP 5
SRR1766444.1025321 chr7 157994860 N chr7 157994939 N DUP 5
SRR1766450.2211671 chr7 157994953 N chr7 157995401 N DEL 5
SRR1766471.10616074 chr7 157995142 N chr7 157995307 N DEL 5
SRR1766470.8900673 chr7 157994749 N chr7 157994951 N DUP 5
SRR1766442.24421643 chr7 157994832 N chr7 157995155 N DUP 6
SRR1766468.143507 chr7 157994771 N chr7 157995176 N DUP 6
SRR1766462.1921776 chr7 157994771 N chr7 157995176 N DUP 9
SRR1766447.2652367 chr7 157994832 N chr7 157995155 N DUP 9
SRR1766479.10692806 chr7 157994850 N chr7 157995218 N DEL 7
SRR1766470.3759027 chr7 157994850 N chr7 157995218 N DEL 7
SRR1766456.4570169 chr7 157994892 N chr7 157995219 N DEL 12
SRR1766464.1898583 chr7 157994927 N chr7 157995253 N DUP 4
SRR1766467.727192 chr7 157994850 N chr7 157995218 N DEL 7
SRR1766461.10448449 chr7 157994850 N chr7 157995218 N DEL 7
SRR1766466.4874667 chr7 157994850 N chr7 157995218 N DEL 12
SRR1766473.11356491 chr7 157994660 N chr7 157995190 N DEL 6
SRR1766466.7139180 chr7 157994661 N chr7 157995191 N DEL 6
SRR1766461.5777529 chr7 157994809 N chr7 157995218 N DEL 12
SRR1766478.1115482 chr7 157994858 N chr7 157995226 N DEL 12
SRR1766460.8932977 chr7 157994874 N chr7 157995240 N DUP 9
SRR1766479.12727241 chr7 157994809 N chr7 157995218 N DEL 6
SRR1766476.6885246 chr7 157994850 N chr7 157995218 N DEL 11
SRR1766445.3981511 chr7 157994809 N chr7 157995218 N DEL 6
SRR1766478.6885597 chr7 157994835 N chr7 157995244 N DEL 11
SRR1766442.12778434 chr7 157994870 N chr7 157995278 N DEL 10
SRR1766476.1377314 chr7 157994659 N chr7 157995231 N DEL 2
SRR1766475.10165586 chr7 157995243 N chr7 157995322 N DUP 5
SRR1766442.13603770 chr7 157995311 N chr7 157995430 N DUP 5
SRR1766452.6302503 chr7 157994853 N chr7 157995342 N DEL 6
SRR1766442.45589070 chr7 157994951 N chr7 157995319 N DEL 5
SRR1766450.1773276 chr7 157994871 N chr7 157995480 N DEL 9
SRR1766477.3405814 chr7 157994834 N chr7 157995484 N DEL 4
SRR1766464.5803569 chr7 157994907 N chr7 157995476 N DEL 5
SRR1766460.1621464 chr7 157994755 N chr7 157995487 N DEL 5
SRR1766463.7774461 chr2 36182096 N chr2 36182155 N DUP 1
SRR1766471.8406063 chr2 36182096 N chr2 36182155 N DUP 6
SRR1766442.16096874 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766443.6334765 chr2 36182198 N chr2 36182379 N DEL 6
SRR1766447.1575509 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766453.8522873 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766445.1310117 chr2 36182114 N chr2 36182199 N DEL 8
SRR1766445.9125244 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766471.1777261 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766482.11346965 chr2 36182150 N chr2 36182205 N DEL 3
SRR1766442.45549660 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766455.2898692 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766462.4787455 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766459.2785444 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766451.2213510 chr2 36182228 N chr2 36182301 N DEL 10
SRR1766470.4532228 chr2 36182231 N chr2 36182304 N DEL 10
SRR1766449.1846243 chr2 36182257 N chr2 36182400 N DUP 10
SRR1766442.5578821 chr2 36182235 N chr2 36182308 N DEL 8
SRR1766470.946016 chr2 36182240 N chr2 36182313 N DEL 3
SRR1766467.665054 chr2 36182229 N chr2 36182302 N DEL 10
SRR1766478.4081387 chr2 36182309 N chr2 36182414 N DUP 12
SRR1766447.1916193 chr2 36182257 N chr2 36182400 N DUP 10
SRR1766442.27504393 chr12 97249742 N chr12 97249793 N DEL 5
SRR1766446.335026 chr12 97249742 N chr12 97249793 N DEL 5
SRR1766462.966500 chr12 97249742 N chr12 97249793 N DEL 5
SRR1766465.2797079 chr22 47647661 N chr22 47647900 N DUP 4
SRR1766452.8877926 chrX 738778 N chrX 738858 N DUP 5
SRR1766467.7387588 chrX 738954 N chrX 739063 N DEL 10
SRR1766442.34995685 chrX 738839 N chrX 739067 N DEL 1
SRR1766448.10505436 chrX 738839 N chrX 739067 N DEL 1
SRR1766477.8673389 chrX 738848 N chrX 739076 N DEL 6
SRR1766452.9190140 chr21 5891865 N chr21 5892138 N DEL 2
SRR1766444.610448 chr21 45452872 N chr21 45453134 N DUP 12
SRR1766467.3745615 chr21 45452872 N chr21 45453134 N DUP 12
SRR1766443.313535 chr21 45452904 N chr21 45452959 N DEL 1
SRR1766478.7693287 chr22 35754187 N chr22 35754496 N DEL 6
SRR1766462.7819178 chr20 53837892 N chr20 53837947 N DUP 18
SRR1766451.2412593 chr20 53837892 N chr20 53837947 N DUP 13
SRR1766463.9996456 chr1 42324194 N chr1 42324285 N DEL 15
SRR1766481.9989619 chr1 42324217 N chr1 42324308 N DEL 10
SRR1766459.4770473 chr1 42324194 N chr1 42324285 N DEL 27
SRR1766481.12724776 chr1 42324208 N chr1 42324297 N DUP 5
SRR1766448.19336 chr1 42324204 N chr1 42324293 N DUP 18
SRR1766485.648402 chr1 42324204 N chr1 42324293 N DUP 18
SRR1766455.5763460 chr1 42324204 N chr1 42324293 N DUP 10
SRR1766444.5503561 chr1 42324204 N chr1 42324293 N DUP 12
SRR1766458.8745256 chr1 42324207 N chr1 42324296 N DUP 8
SRR1766457.2180570 chr1 42324225 N chr1 42324292 N DEL 9
SRR1766486.496162 chr1 42324391 N chr1 42324446 N DUP 2
SRR1766478.243561 chr6 65443284 N chr6 65443347 N DUP 9
SRR1766442.5989375 chr6 65443284 N chr6 65443347 N DUP 11
SRR1766462.1760252 chr6 65443405 N chr6 65443470 N DEL 1
SRR1766462.9209368 chr6 65443405 N chr6 65443470 N DEL 2
SRR1766446.4756085 chr6 65443281 N chr6 65443332 N DEL 7
SRR1766442.3554828 chr6 65443311 N chr6 65443378 N DEL 11
SRR1766443.6485012 chr6 65443311 N chr6 65443378 N DEL 11
SRR1766442.31688981 chr6 65443311 N chr6 65443378 N DEL 11
SRR1766457.2957956 chr6 65443311 N chr6 65443378 N DEL 10
SRR1766453.7950980 chr6 65443311 N chr6 65443378 N DEL 10
SRR1766481.6748158 chr2 238769470 N chr2 238769574 N DEL 1
SRR1766455.6205566 chr2 238769437 N chr2 238769550 N DEL 13
SRR1766481.11335399 chrX 118709201 N chrX 118709638 N DEL 5
SRR1766449.3599290 chrX 118709201 N chrX 118709638 N DEL 5
SRR1766463.4458631 chrX 118709224 N chrX 118709661 N DUP 6
SRR1766486.692995 chr2 122274144 N chr2 122274269 N DEL 21
SRR1766450.1531917 chr4 3919303 N chr4 3919454 N DEL 8
SRR1766455.1407251 chr4 3919303 N chr4 3919454 N DEL 9
SRR1766450.7920914 chr4 3919305 N chr4 3919454 N DEL 11
SRR1766474.5937043 chr4 3919299 N chr4 3919449 N DUP 7
SRR1766482.3859369 chr4 160510962 N chr4 160511078 N DEL 2
SRR1766486.4488070 chr4 160510961 N chr4 160511083 N DEL 3
SRR1766480.6247684 chr3 103072314 N chr3 103072379 N DUP 7
SRR1766464.10344375 chr3 103072314 N chr3 103072379 N DUP 9
SRR1766480.1997618 chr3 103072314 N chr3 103072379 N DUP 9
SRR1766469.3236365 chr3 103072314 N chr3 103072379 N DUP 9
SRR1766466.6797563 chr3 103072314 N chr3 103072379 N DUP 9
SRR1766483.10920300 chr3 103072314 N chr3 103072379 N DUP 9
SRR1766458.8587764 chr3 103072314 N chr3 103072379 N DUP 9
SRR1766448.8700463 chr3 103072314 N chr3 103072379 N DUP 9
SRR1766443.6572958 chr3 103072314 N chr3 103072379 N DUP 9
SRR1766442.47061987 chr3 103072362 N chr3 103072427 N DEL 9
SRR1766448.6407016 chr3 103072362 N chr3 103072427 N DEL 9
SRR1766479.5627308 chr3 103072362 N chr3 103072427 N DEL 9
SRR1766482.8026115 chr3 103072362 N chr3 103072427 N DEL 9
SRR1766454.5769396 chr3 103072362 N chr3 103072427 N DEL 9
SRR1766452.1273220 chr3 103072362 N chr3 103072427 N DEL 9
SRR1766442.37997981 chr3 103072362 N chr3 103072427 N DEL 9
SRR1766443.11110433 chr3 103072296 N chr3 103072427 N DEL 9
SRR1766448.3136072 chr3 103072296 N chr3 103072427 N DEL 9
SRR1766486.7199176 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766466.7073609 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766455.4791355 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766475.10743860 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766465.8455944 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766471.8115941 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766457.2160918 chr12 6399412 N chr12 6399789 N DEL 3
SRR1766463.10901242 chr12 6399368 N chr12 6399555 N DUP 5
SRR1766447.757403 chr12 6399379 N chr12 6399566 N DUP 2
SRR1766483.4589219 chr12 6399380 N chr12 6399567 N DUP 1
SRR1766463.3888570 chr12 6399376 N chr12 6399563 N DUP 5
SRR1766445.3441349 chr12 6399473 N chr12 6399848 N DUP 5
SRR1766461.3036370 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766458.335083 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766451.3969012 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766457.9248681 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766442.20429786 chr12 6399361 N chr12 6399550 N DEL 5
SRR1766461.10397281 chr12 6399366 N chr12 6399553 N DUP 1
SRR1766460.7835548 chr12 6399366 N chr12 6399553 N DUP 5
SRR1766466.7078893 chr12 6399366 N chr12 6399553 N DUP 5
SRR1766481.4644535 chr12 6399366 N chr12 6399553 N DUP 5
SRR1766446.3146874 chr12 6399366 N chr12 6399553 N DUP 5
SRR1766457.4541576 chr12 6399367 N chr12 6399554 N DUP 5
SRR1766477.9327118 chr12 6399368 N chr12 6399555 N DUP 5
SRR1766473.6360937 chr12 6399369 N chr12 6399556 N DUP 5
SRR1766452.3530878 chr12 6399371 N chr12 6399558 N DUP 5
SRR1766475.2615503 chr12 6399484 N chr12 6399673 N DEL 5
SRR1766476.9173809 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766442.18002623 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766467.7837058 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766444.5653331 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766458.2786256 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766481.11479095 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766484.3319637 chr12 6399483 N chr12 6399672 N DEL 5
SRR1766459.8405718 chr12 6399484 N chr12 6399673 N DEL 5
SRR1766456.2472339 chr12 6399485 N chr12 6399674 N DEL 5
SRR1766442.1987578 chr12 6399361 N chr12 6399738 N DEL 5
SRR1766449.10808301 chr1 23173465 N chr1 23173521 N DEL 5
SRR1766460.8351104 chr1 23173465 N chr1 23173521 N DEL 5
SRR1766485.10823155 chr5 158582790 N chr5 158583061 N DEL 7
SRR1766480.7368196 chr5 158582707 N chr5 158583006 N DUP 10
SRR1766475.6662371 chr5 158582832 N chr5 158583332 N DEL 5
SRR1766462.11019012 chr5 158582812 N chr5 158583082 N DUP 5
SRR1766445.1993163 chr5 158582961 N chr5 158583285 N DEL 8
SRR1766452.72925 chr5 158582999 N chr5 158583323 N DEL 10
SRR1766450.2095519 chr5 158582904 N chr5 158583030 N DUP 3
SRR1766475.4422922 chr5 158582879 N chr5 158583005 N DUP 5
SRR1766467.8364024 chr5 158583032 N chr5 158583454 N DEL 5
SRR1766467.977255 chr5 158583079 N chr5 158583501 N DEL 5
SRR1766474.1888789 chr5 158582841 N chr5 158583114 N DUP 5
SRR1766465.6983568 chr5 158582935 N chr5 158583063 N DEL 7
SRR1766460.2405654 chr5 158582895 N chr5 158583119 N DUP 5
SRR1766485.12076664 chr5 158582858 N chr5 158583084 N DEL 1
SRR1766451.3819984 chr5 158583104 N chr5 158583426 N DUP 5
SRR1766474.3017455 chr5 158582953 N chr5 158583130 N DEL 5
SRR1766456.6188695 chr5 158583151 N chr5 158583375 N DUP 15
SRR1766442.10595909 chr5 158583249 N chr5 158583328 N DEL 6
SRR1766483.5891433 chr5 158583252 N chr5 158583331 N DEL 1
SRR1766472.7987703 chr5 158582863 N chr5 158583187 N DEL 1
SRR1766482.7901179 chr5 158583270 N chr5 158583545 N DEL 1
SRR1766452.441225 chr5 158582950 N chr5 158583225 N DEL 2
SRR1766442.8780358 chr5 158582935 N chr5 158583259 N DEL 5
SRR1766476.1186937 chr5 158583328 N chr5 158583601 N DUP 5
SRR1766486.2165560 chr5 158583323 N chr5 158583596 N DUP 5
SRR1766460.2250089 chr5 158583323 N chr5 158583596 N DUP 5
SRR1766450.10172292 chr5 158583330 N chr5 158583603 N DUP 5
SRR1766449.5175158 chr5 158583011 N chr5 158583335 N DEL 1
SRR1766478.2484870 chr5 158583382 N chr5 158583528 N DUP 5
SRR1766472.930962 chr5 158582986 N chr5 158583582 N DUP 10
SRR1766457.1309895 chrX 62523280 N chrX 62523790 N DEL 9
SRR1766485.5102688 chrX 62523394 N chrX 62523731 N DUP 1
SRR1766442.35815738 chrX 62523363 N chrX 62523533 N DUP 5
SRR1766452.5630979 chrX 62523676 N chrX 62524186 N DEL 5
SRR1766449.8637137 chrX 62523322 N chrX 62523832 N DEL 10
SRR1766485.6609093 chrX 62523940 N chrX 62524112 N DEL 10
SRR1766480.1648543 chrX 62523355 N chrX 62523525 N DUP 10
SRR1766478.11978237 chrX 62523591 N chrX 62524101 N DEL 5
SRR1766467.1461203 chrX 62523742 N chrX 62524252 N DEL 25
SRR1766464.2484636 chrX 62523414 N chrX 62524767 N DEL 5
SRR1766472.6811732 chr15 78373784 N chr15 78373875 N DUP 1
SRR1766460.3028012 chr15 78373872 N chr15 78373925 N DUP 10
SRR1766450.1400025 chr15 78373799 N chr15 78373888 N DEL 2
SRR1766478.9147209 chr7 100970811 N chr7 100970936 N DEL 2
SRR1766442.18635948 chr5 145742265 N chr5 145742354 N DEL 12
SRR1766461.4868162 chr5 145742264 N chr5 145742353 N DEL 13
SRR1766485.3981109 chr6 168044283 N chr6 168044533 N DEL 4
SRR1766459.5657206 chr6 168044285 N chr6 168044407 N DUP 5
SRR1766470.2789417 chr6 168044293 N chr6 168044415 N DUP 5
SRR1766442.31986657 chr6 168044452 N chr6 168044534 N DUP 5
SRR1766456.5364479 chr6 168044308 N chr6 168044475 N DEL 6
SRR1766456.4979845 chr6 168044326 N chr6 168044533 N DEL 5
SRR1766484.7608245 chr6 168044620 N chr6 168044788 N DUP 5
SRR1766463.450881 chr6 168044543 N chr6 168044673 N DEL 5
SRR1766476.4714898 chr6 168044533 N chr6 168044744 N DUP 5
SRR1766470.3183711 chr6 168044327 N chr6 168044789 N DEL 23
SRR1766465.6295866 chr6 168044332 N chr6 168044794 N DEL 5
SRR1766475.9077804 chr17 21235992 N chr17 21236722 N DEL 8
SRR1766469.6388566 chr17 21235999 N chr17 21236725 N DEL 5
SRR1766457.583913 chr17 21236030 N chr17 21236295 N DEL 5
SRR1766476.9709638 chr17 21236030 N chr17 21236295 N DEL 6
SRR1766477.2671457 chr17 21236030 N chr17 21236309 N DUP 3
SRR1766464.1589747 chr17 21236171 N chr17 21236723 N DEL 7
SRR1766479.5459461 chr17 21236168 N chr17 21236720 N DEL 8
SRR1766473.10051906 chr17 21236107 N chr17 21236178 N DUP 1
SRR1766465.5923299 chr17 21236038 N chr17 21236185 N DEL 1
SRR1766445.3523783 chr17 21236038 N chr17 21236213 N DEL 6
SRR1766457.6281789 chr17 21236243 N chr17 21236380 N DUP 5
SRR1766479.6146588 chr17 21236149 N chr17 21236254 N DEL 5
SRR1766455.1913097 chr17 21236262 N chr17 21236736 N DUP 6
SRR1766455.8371815 chr17 21235981 N chr17 21236406 N DUP 5
SRR1766466.9191287 chr17 21236281 N chr17 21236422 N DUP 1
SRR1766478.6204976 chr17 21236631 N chr17 21236710 N DUP 5
SRR1766466.7102673 chr17 21236631 N chr17 21236710 N DUP 5
SRR1766475.4691188 chr17 21236631 N chr17 21236710 N DUP 5
SRR1766474.5706260 chr17 21236631 N chr17 21236710 N DUP 5
SRR1766457.5094193 chr7 155932809 N chr7 155933018 N DEL 13
SRR1766467.402072 chr7 155932809 N chr7 155933018 N DEL 19
SRR1766482.5016453 chr7 155932809 N chr7 155933018 N DEL 16
SRR1766463.1642958 chr3 179032608 N chr3 179032725 N DEL 6
SRR1766454.2465506 chr3 179032687 N chr3 179032921 N DEL 5
SRR1766478.10092968 chr3 179032803 N chr3 179032921 N DEL 5
SRR1766469.10628306 chr3 179032622 N chr3 179032739 N DEL 1
SRR1766460.6080464 chr3 179032643 N chr3 179032797 N DEL 5
SRR1766462.5972052 chr21 42348741 N chr21 42348838 N DUP 5
SRR1766445.201821 chr21 42348756 N chr21 42348855 N DEL 6
SRR1766485.5808584 chr21 42349017 N chr21 42349206 N DUP 5
SRR1766477.6075710 chr21 42349171 N chr21 42349248 N DUP 3
SRR1766452.7597640 chr21 42349171 N chr21 42349322 N DUP 5
SRR1766481.12504452 chr21 42348766 N chr21 42349236 N DEL 8
SRR1766479.4235537 chr21 42349289 N chr21 42349366 N DUP 5
SRR1766483.10025292 chr21 42349289 N chr21 42349366 N DUP 5
SRR1766483.7209969 chr21 42349289 N chr21 42349366 N DUP 5
SRR1766451.7273075 chr21 42349289 N chr21 42349366 N DUP 10
SRR1766461.5423633 chr21 42349016 N chr21 42349460 N DUP 1
SRR1766484.1086883 chr21 42349027 N chr21 42349471 N DUP 5
SRR1766475.6046822 chr5 117993527 N chr5 117993580 N DEL 9
SRR1766480.219519 chr5 117993527 N chr5 117993580 N DEL 12
SRR1766446.1599666 chr5 117993527 N chr5 117993580 N DEL 13
SRR1766442.11850697 chr5 117993528 N chr5 117993579 N DUP 5
SRR1766482.11208196 chr5 117993528 N chr5 117993579 N DUP 5
SRR1766474.1092769 chr5 117993518 N chr5 117993589 N DUP 5
SRR1766475.10193603 chr5 117993542 N chr5 117993595 N DEL 5
SRR1766467.3757217 chr5 117993545 N chr5 117993598 N DEL 5
SRR1766452.4998773 chr5 117993533 N chr5 117993606 N DEL 2
SRR1766448.10222591 chr5 117993534 N chr5 117993607 N DEL 1
SRR1766446.4916002 chr1 154714107 N chr1 154714760 N DEL 6
SRR1766442.28923231 chr1 154714107 N chr1 154714760 N DEL 9
SRR1766485.7620708 chr1 154714107 N chr1 154714760 N DEL 22
SRR1766484.6011862 chr1 154714107 N chr1 154714760 N DEL 22
SRR1766460.8417822 chr1 154714117 N chr1 154714693 N DEL 25
SRR1766447.2360655 chr1 154714147 N chr1 154714321 N DEL 5
SRR1766457.2030254 chr1 154714109 N chr1 154714339 N DUP 14
SRR1766461.8880584 chr1 154714216 N chr1 154714778 N DUP 1
SRR1766442.22327055 chr1 154714220 N chr1 154714709 N DUP 1
SRR1766469.3833488 chr1 154714159 N chr1 154714239 N DEL 5
SRR1766457.8843065 chr1 154714164 N chr1 154714379 N DUP 9
SRR1766442.11661224 chr1 154714167 N chr1 154714268 N DEL 6
SRR1766448.849667 chr1 154714288 N chr1 154714343 N DUP 4
SRR1766475.8181005 chr1 154714167 N chr1 154714303 N DEL 5
SRR1766442.19833827 chr1 154714274 N chr1 154714331 N DEL 23
SRR1766477.749271 chr1 154714331 N chr1 154714762 N DUP 17
SRR1766455.3191781 chr1 154714297 N chr1 154714354 N DEL 29
SRR1766478.8201486 chr1 154714192 N chr1 154714328 N DEL 2
SRR1766455.3191781 chr1 154714319 N chr1 154714691 N DUP 10
SRR1766444.1959785 chr1 154714375 N chr1 154714618 N DUP 10
SRR1766478.1726538 chr1 154714354 N chr1 154714716 N DUP 7
SRR1766459.3707523 chr1 154714163 N chr1 154714340 N DEL 8
SRR1766453.5342074 chr1 154714326 N chr1 154714486 N DUP 5
SRR1766469.2821435 chr1 154714381 N chr1 154714432 N DUP 11
SRR1766442.40563046 chr1 154714349 N chr1 154714427 N DEL 10
SRR1766486.2104134 chr1 154714468 N chr1 154714535 N DUP 15
SRR1766468.2370654 chr1 154714451 N chr1 154714631 N DUP 16
SRR1766453.2898949 chr1 154714526 N chr1 154714703 N DUP 11
SRR1766475.6450498 chr1 154714290 N chr1 154714532 N DEL 11
SRR1766442.21178965 chr1 154714141 N chr1 154714587 N DUP 26
SRR1766446.6990697 chr1 154714457 N chr1 154714607 N DEL 27
SRR1766481.10293459 chr1 154714139 N chr1 154714587 N DUP 24
SRR1766456.140230 chr1 154714457 N chr1 154714607 N DEL 35
SRR1766463.2151502 chr1 154714595 N chr1 154714734 N DUP 8
SRR1766485.75103 chr1 154714183 N chr1 154714580 N DEL 13
SRR1766467.10907432 chr1 154714134 N chr1 154714687 N DUP 26
SRR1766448.9273968 chr1 154714195 N chr1 154714762 N DEL 11
SRR1766470.2783005 chr1 154714599 N chr1 154714784 N DEL 12
SRR1766478.504357 chr1 154714352 N chr1 154714749 N DEL 10
SRR1766461.6421249 chr1 154714131 N chr1 154714762 N DEL 6
SRR1766460.126957 chr1 154714655 N chr1 154714786 N DEL 27
SRR1766462.8055582 chr16 34696431 N chr16 34696482 N DUP 10
SRR1766442.12016444 chr16 34696431 N chr16 34696482 N DUP 12
SRR1766465.2750913 chr16 34696431 N chr16 34696482 N DUP 16
SRR1766456.5369754 chr16 34696424 N chr16 34696524 N DUP 3
SRR1766442.28192804 chr16 34696417 N chr16 34696566 N DUP 8
SRR1766442.28153173 chr5 2594850 N chr5 2594909 N DUP 5
SRR1766453.528881 chr18 78753331 N chr18 78753577 N DEL 5
SRR1766483.11619175 chr18 78753462 N chr18 78753559 N DUP 5
SRR1766479.8402732 chr18 78753265 N chr18 78753462 N DEL 5
SRR1766443.684211 chr18 78753404 N chr18 78753503 N DEL 6
SRR1766443.6815422 chr18 78753264 N chr18 78753510 N DEL 3
SRR1766469.3162155 chr18 78753385 N chr18 78753533 N DEL 5
SRR1766478.1978258 chr5 345605 N chr5 345766 N DEL 5
SRR1766442.13854475 chr18 76587085 N chr18 76587307 N DEL 3
SRR1766479.2708796 chr18 76587105 N chr18 76587412 N DEL 33
SRR1766442.28804863 chr18 76587337 N chr18 76587389 N DEL 2
SRR1766470.2287325 chr18 76587337 N chr18 76587389 N DEL 5
SRR1766455.5916173 chr18 76587139 N chr18 76587293 N DEL 33
SRR1766480.2862494 chr18 76587059 N chr18 76587281 N DEL 15
SRR1766442.29225713 chr18 76587139 N chr18 76587293 N DEL 10
SRR1766447.73621 chr18 76587183 N chr18 76587303 N DEL 2
SRR1766467.3619138 chr18 76587029 N chr18 76587319 N DEL 11
SRR1766481.4038627 chr18 76587178 N chr18 76587332 N DEL 20
SRR1766456.3999652 chr18 76587048 N chr18 76587338 N DEL 30
SRR1766479.6528123 chr18 76587107 N chr18 76587329 N DEL 1
SRR1766480.6543590 chr18 76587176 N chr18 76587330 N DEL 5
SRR1766449.7258227 chr18 76587038 N chr18 76587396 N DEL 9
SRR1766450.7519023 chr18 76587089 N chr18 76587447 N DEL 5
SRR1766472.11008716 chr18 76587343 N chr18 76587480 N DEL 8
SRR1766458.9558801 chr18 76587262 N chr18 76587484 N DEL 5
SRR1766479.2930650 chr18 76587051 N chr18 76587528 N DEL 2
SRR1766458.1976028 chr9 72841809 N chr9 72841887 N DEL 8
SRR1766446.9074980 chr9 72841549 N chr9 72841920 N DUP 6
SRR1766475.2959095 chr9 72841562 N chr9 72842091 N DEL 7
SRR1766471.7479747 chr4 56780935 N chr4 56781246 N DEL 3
SRR1766476.445555 chr4 56781379 N chr4 56781512 N DUP 5
SRR1766480.4473228 chr16 89995321 N chr16 89995562 N DUP 5
SRR1766446.1731880 chr16 89995295 N chr16 89995441 N DUP 10
SRR1766465.9690040 chr16 89995446 N chr16 89995648 N DEL 5
SRR1766466.3150333 chr16 89995371 N chr16 89995506 N DUP 2
SRR1766442.42932604 chr16 89995549 N chr16 89995751 N DEL 5
SRR1766451.998448 chr16 89995453 N chr16 89995588 N DUP 1
SRR1766486.7319728 chr16 89995563 N chr16 89995765 N DEL 4
SRR1766442.14038791 chr16 89995492 N chr16 89995692 N DUP 2
SRR1766442.37976682 chr16 89995492 N chr16 89995692 N DUP 5
SRR1766478.9729536 chr16 89995492 N chr16 89995692 N DUP 5
SRR1766481.7847116 chr16 89995549 N chr16 89995751 N DEL 5
SRR1766445.7818242 chr16 89995549 N chr16 89995751 N DEL 5
SRR1766442.13071150 chr16 89995549 N chr16 89995751 N DEL 5
SRR1766480.4876650 chr16 89995413 N chr16 89995751 N DEL 5
SRR1766481.4371635 chr16 89995413 N chr16 89995751 N DEL 5
SRR1766470.3431046 chr16 89995413 N chr16 89995751 N DEL 5
SRR1766467.1758082 chr16 89995413 N chr16 89995751 N DEL 5
SRR1766481.7847116 chr16 89995413 N chr16 89995751 N DEL 5
SRR1766484.5355982 chr16 89995420 N chr16 89995758 N DEL 5
SRR1766457.7057130 chr16 89995413 N chr16 89995751 N DEL 5
SRR1766446.8819600 chr16 89995413 N chr16 89995751 N DEL 5
SRR1766470.6744108 chr5 32158113 N chr5 32158227 N DEL 8
SRR1766473.6594944 chr5 32158113 N chr5 32158227 N DEL 9
SRR1766457.5207991 chr5 32158113 N chr5 32158227 N DEL 9
SRR1766461.3207899 chr5 32158173 N chr5 32158287 N DUP 24
SRR1766462.5485256 chr5 32158136 N chr5 32158240 N DUP 6
SRR1766456.6140935 chr14 67193288 N chr14 67193341 N DEL 2
SRR1766442.15357695 chr14 67193288 N chr14 67193341 N DEL 4
SRR1766448.5628682 chr14 67193288 N chr14 67193341 N DEL 4
SRR1766466.11219754 chr14 67193291 N chr14 67193344 N DEL 9
SRR1766466.2206216 chr14 67193293 N chr14 67193346 N DEL 9
SRR1766445.1962853 chr11 42130724 N chr11 42130821 N DUP 2
SRR1766453.3121693 chr13 108258351 N chr13 108258400 N DUP 2
SRR1766467.11887624 chr13 108258351 N chr13 108258400 N DUP 4
SRR1766442.13571049 chr13 108258351 N chr13 108258400 N DUP 10
SRR1766478.8389258 chr13 108258351 N chr13 108258400 N DUP 10
SRR1766482.3535483 chr13 108258351 N chr13 108258400 N DUP 11
SRR1766476.11208833 chr13 108258351 N chr13 108258400 N DUP 12
SRR1766482.2054380 chr13 108258351 N chr13 108258400 N DUP 14
SRR1766483.5987532 chr13 108258355 N chr13 108258404 N DUP 25
SRR1766486.7066633 chr13 108258351 N chr13 108258400 N DUP 25
SRR1766465.4632427 chr13 108258351 N chr13 108258400 N DUP 25
SRR1766442.22260542 chr13 108258351 N chr13 108258400 N DUP 25
SRR1766469.18885 chr13 108258351 N chr13 108258400 N DUP 25
SRR1766455.1415730 chr13 108258351 N chr13 108258400 N DUP 27
SRR1766458.3779198 chr13 108258351 N chr13 108258400 N DUP 38
SRR1766459.1118596 chr13 108258351 N chr13 108258400 N DUP 20
SRR1766457.626318 chr13 108258351 N chr13 108258400 N DUP 24
SRR1766462.6406353 chr13 108258355 N chr13 108258404 N DUP 11
SRR1766454.1694565 chr13 108258363 N chr13 108258412 N DUP 3
SRR1766486.5008663 chr13 108258358 N chr13 108258407 N DUP 8
SRR1766476.5562289 chr2 183354507 N chr2 183354582 N DEL 9
SRR1766484.4674193 chr2 183354509 N chr2 183354582 N DEL 7
SRR1766472.3017673 chr2 183354507 N chr2 183354582 N DEL 9
SRR1766474.2672440 chr2 183354509 N chr2 183354582 N DEL 7
SRR1766465.11329254 chr2 183354509 N chr2 183354582 N DEL 7
SRR1766467.5727611 chr2 183354496 N chr2 183354587 N DEL 7
SRR1766483.4548854 chr2 183354506 N chr2 183354597 N DEL 1
SRR1766471.11447794 chr6 87128693 N chr6 87128744 N DUP 5
SRR1766470.827127 chr6 87128747 N chr6 87129270 N DEL 5
SRR1766445.7686164 chr6 87128747 N chr6 87129270 N DEL 5
SRR1766461.10317996 chr6 87128747 N chr6 87129270 N DEL 5
SRR1766477.5453663 chr6 87128747 N chr6 87129270 N DEL 5
SRR1766484.9283612 chr6 87128747 N chr6 87129270 N DEL 5
SRR1766450.4028698 chr6 87128765 N chr6 87129286 N DUP 5
SRR1766452.1040527 chr6 87128766 N chr6 87129287 N DUP 4
SRR1766486.11586897 chr6 87128835 N chr6 87128893 N DEL 6
SRR1766464.2253457 chr6 87128836 N chr6 87128894 N DEL 5
SRR1766462.7163229 chr6 87128940 N chr6 87129013 N DEL 10
SRR1766463.9171038 chr6 87128940 N chr6 87129013 N DEL 10
SRR1766481.4629916 chr6 87128940 N chr6 87129013 N DEL 9
SRR1766445.5011150 chr6 87128940 N chr6 87129013 N DEL 5
SRR1766442.14631556 chr6 87128940 N chr6 87129013 N DEL 5
SRR1766470.7655035 chr6 87128940 N chr6 87129013 N DEL 5
SRR1766455.7416900 chr6 87128940 N chr6 87129013 N DEL 5
SRR1766471.6435097 chr6 87129128 N chr6 87129267 N DEL 2
SRR1766475.8137547 chr6 87128696 N chr6 87129131 N DUP 9
SRR1766472.11713734 chr6 87129128 N chr6 87129267 N DEL 5
SRR1766464.4581255 chr6 87129128 N chr6 87129195 N DEL 1
SRR1766459.10130850 chr6 87129128 N chr6 87129195 N DEL 2
SRR1766452.5666579 chr6 87129128 N chr6 87129195 N DEL 7
SRR1766473.6069674 chr6 87129128 N chr6 87129195 N DEL 7
SRR1766479.13839151 chr6 87129128 N chr6 87129195 N DEL 8
SRR1766483.10743055 chr6 87129128 N chr6 87129195 N DEL 11
SRR1766443.3975051 chr6 87129128 N chr6 87129195 N DEL 13
SRR1766460.1351232 chr6 87129132 N chr6 87129195 N DUP 7
SRR1766486.447320 chr6 87129198 N chr6 87129265 N DUP 14
SRR1766455.6589869 chr6 87129166 N chr6 87129281 N DEL 5
SRR1766446.3787980 chr6 87129166 N chr6 87129281 N DEL 5
SRR1766474.10607700 chr6 87129166 N chr6 87129281 N DEL 5
SRR1766457.4107451 chr6 87129166 N chr6 87129281 N DEL 5
SRR1766450.4028698 chr6 87129143 N chr6 87129282 N DEL 5
SRR1766442.26665241 chr6 87129149 N chr6 87129288 N DEL 5
SRR1766447.6596045 chr6 87129160 N chr6 87129299 N DEL 5
SRR1766450.1746966 chr6 87129112 N chr6 87129299 N DEL 2
SRR1766453.8379490 chr17 79709755 N chr17 79710018 N DEL 4
SRR1766485.6501083 chr17 79710185 N chr17 79710272 N DUP 5
SRR1766475.95061 chr17 79709798 N chr17 79710193 N DEL 5
SRR1766463.10901475 chr17 79709877 N chr17 79710228 N DEL 1
SRR1766456.3004998 chr17 79710017 N chr17 79710368 N DEL 7
SRR1766482.4066739 chr17 79710018 N chr17 79710369 N DEL 6
SRR1766453.10238915 chr17 79710326 N chr17 79710414 N DEL 5
SRR1766449.1395501 chr17 79709889 N chr17 79710414 N DEL 17
SRR1766464.3869662 chr17 79709801 N chr17 79710414 N DEL 10
SRR1766471.8083702 chr17 79709821 N chr17 79710434 N DEL 8
SRR1766444.1493031 chr1 3502169 N chr1 3502247 N DUP 5
SRR1766474.11674704 chr1 3502172 N chr1 3502250 N DUP 25
SRR1766484.9346968 chr1 3502173 N chr1 3502251 N DUP 17
SRR1766445.7114706 chr1 243480506 N chr1 243480659 N DEL 3
SRR1766452.744684 chr1 243480510 N chr1 243480676 N DEL 2
SRR1766466.10579947 chr1 243480673 N chr1 243480751 N DUP 1
SRR1766454.8844611 chr1 243480544 N chr1 243480982 N DUP 19
SRR1766442.3456664 chr1 243480494 N chr1 243480948 N DUP 5
SRR1766483.6288009 chr1 243480793 N chr1 243481044 N DUP 18
SRR1766470.6972473 chr1 243480740 N chr1 243480906 N DEL 14
SRR1766462.7343981 chr1 243480580 N chr1 243480923 N DEL 10
SRR1766448.10728698 chr1 243480839 N chr1 243481059 N DEL 12
SRR1766485.10566962 chr2 89805048 N chr2 89805489 N DUP 5
SRR1766472.3168133 chr9 24739245 N chr9 24739363 N DUP 10
SRR1766476.10574619 chr6 116511255 N chr6 116511334 N DEL 2
SRR1766455.8863854 chr17 68001819 N chr17 68002124 N DEL 5
SRR1766467.321575 chr17 68001923 N chr17 68002228 N DEL 10
SRR1766448.4928990 chr17 68001933 N chr17 68003211 N DEL 5
SRR1766460.2710532 chr17 68001933 N chr17 68002238 N DEL 1
SRR1766460.9412751 chr17 68001953 N chr17 68002256 N DUP 3
SRR1766474.4290743 chr17 68002099 N chr17 68002400 N DEL 11
SRR1766442.25779218 chr17 68002245 N chr17 68002555 N DEL 10
SRR1766472.4209483 chr17 68001843 N chr17 68002148 N DEL 5
SRR1766482.2177939 chr17 68002260 N chr17 68002570 N DEL 7
SRR1766466.6402297 chr17 68001902 N chr17 68002207 N DEL 5
SRR1766442.5445257 chr17 68001906 N chr17 68002211 N DEL 5
SRR1766470.5701292 chr17 68001906 N chr17 68002211 N DEL 4
SRR1766461.6679482 chr17 68002263 N chr17 68002571 N DUP 5
SRR1766462.9456503 chr17 68002388 N chr17 68002699 N DEL 8
SRR1766475.2754809 chr17 68002113 N chr17 68002411 N DEL 4
SRR1766471.6344186 chr17 68002451 N chr17 68003116 N DEL 10
SRR1766472.11611706 chr17 68001848 N chr17 68002462 N DEL 4
SRR1766448.4928990 chr17 68001852 N chr17 68002466 N DEL 8
SRR1766461.3991952 chr17 68002098 N chr17 68002746 N DUP 5
SRR1766452.1606936 chr17 68001812 N chr17 68002764 N DEL 2
SRR1766450.2039784 chr17 68002335 N chr17 68002981 N DUP 1
SRR1766479.4092345 chr17 68002232 N chr17 68003204 N DUP 10
SRR1766485.10355801 chr17 68002634 N chr17 68003297 N DUP 1
SRR1766455.8001013 chr1 1192538 N chr1 1192707 N DEL 5
SRR1766470.8696700 chr1 1192538 N chr1 1192755 N DEL 10
SRR1766479.13223392 chr1 1192538 N chr1 1192926 N DEL 10
SRR1766450.3461519 chr1 1192564 N chr1 1192928 N DEL 1
SRR1766442.6204395 chr1 1192511 N chr1 1192678 N DUP 5
SRR1766466.8376865 chr1 1192631 N chr1 1192726 N DUP 5
SRR1766443.1267782 chr1 1192725 N chr1 1192921 N DEL 10
SRR1766480.5765364 chr1 1192565 N chr1 1192756 N DUP 5
SRR1766447.8577169 chr1 1192530 N chr1 1192723 N DEL 5
SRR1766457.3500556 chr1 1192776 N chr1 1192919 N DUP 5
SRR1766473.9500448 chr1 1192617 N chr1 1192834 N DEL 5
SRR1766469.2894144 chr1 1192610 N chr1 1192827 N DEL 10
SRR1766447.8631782 chr1 1192605 N chr1 1192822 N DEL 5
SRR1766471.1972827 chr1 1192617 N chr1 1192834 N DEL 15
SRR1766449.8500478 chr1 1192593 N chr1 1192834 N DEL 15
SRR1766462.4778579 chr1 1192617 N chr1 1192858 N DEL 11
SRR1766461.9957839 chr1 1192522 N chr1 1192958 N DEL 3
SRR1766442.13628522 chr10 132605310 N chr10 132605568 N DUP 10
SRR1766442.4591318 chr16 89074437 N chr16 89074673 N DEL 5
SRR1766469.8593948 chr16 89074450 N chr16 89074686 N DEL 5
SRR1766483.5560985 chr16 89074172 N chr16 89074437 N DEL 5
SRR1766455.1166976 chr16 89074536 N chr16 89074770 N DUP 5
SRR1766451.326249 chr16 89074496 N chr16 89074583 N DUP 4
SRR1766481.8762153 chr16 89074522 N chr16 89074858 N DUP 5
SRR1766456.4023159 chr16 89074320 N chr16 89074555 N DEL 16
SRR1766451.10215156 chr16 89074175 N chr16 89074528 N DEL 5
SRR1766485.9799571 chr16 89074281 N chr16 89074531 N DEL 5
SRR1766450.3307004 chr16 89074290 N chr16 89074555 N DEL 10
SRR1766456.2098082 chr16 89074207 N chr16 89074545 N DEL 5
SRR1766455.748114 chr16 89074657 N chr16 89074773 N DUP 5
SRR1766464.4832032 chr16 89074517 N chr16 89074665 N DEL 7
SRR1766473.1820778 chr16 89074752 N chr16 89074900 N DEL 5
SRR1766467.9624119 chr16 89074899 N chr16 89075119 N DEL 4
SRR1766469.8593948 chr16 89074369 N chr16 89074868 N DEL 5
SRR1766460.5125643 chr16 89074390 N chr16 89075005 N DUP 5
SRR1766442.44321818 chr16 89074390 N chr16 89075005 N DUP 5
SRR1766442.23745286 chr16 89074282 N chr16 89074973 N DEL 2
SRR1766475.7925597 chr16 89074858 N chr16 89075021 N DEL 5
SRR1766460.3361399 chr16 89074858 N chr16 89075021 N DEL 5
SRR1766486.8710236 chr16 89075081 N chr16 89075182 N DUP 1
SRR1766452.6858549 chr16 29197810 N chr16 29197984 N DUP 5
SRR1766442.29339462 chr10 132965341 N chr10 132965854 N DEL 10
SRR1766458.998726 chr10 132965277 N chr10 132965515 N DEL 5
SRR1766481.6927545 chr10 132965287 N chr10 132965525 N DEL 5
SRR1766446.5448719 chr10 132965434 N chr10 132965537 N DEL 5
SRR1766472.7492583 chr10 132965506 N chr10 132965710 N DEL 5
SRR1766452.9452001 chr10 132965332 N chr10 132965537 N DEL 5
SRR1766483.2854918 chr10 132965342 N chr10 132965545 N DUP 4
SRR1766458.4112546 chr13 58176973 N chr13 58177057 N DEL 6
SRR1766442.14699963 chr13 58176973 N chr13 58177057 N DEL 6
SRR1766485.7688781 chr13 58176977 N chr13 58177057 N DEL 9
SRR1766463.1494801 chr13 58176976 N chr13 58177048 N DUP 2
SRR1766466.2426217 chr13 58176976 N chr13 58177042 N DUP 12
SRR1766444.3076545 chr13 58177024 N chr13 58177088 N DEL 5
SRR1766462.10163603 chr17 2034659 N chr17 2034891 N DEL 10
SRR1766448.97907 chr19 52554530 N chr19 52555035 N DEL 30
SRR1766481.13234930 chr19 52554561 N chr19 52555318 N DEL 10
SRR1766453.9014228 chr19 52554082 N chr19 52554669 N DUP 5
SRR1766459.11038634 chr19 52554116 N chr19 52554787 N DUP 1
SRR1766446.2265413 chr19 52554136 N chr19 52554809 N DEL 12
SRR1766456.2387469 chr19 52555013 N chr19 52555182 N DEL 25
SRR1766458.46167 chr19 52554544 N chr19 52555049 N DEL 30
SRR1766449.4634801 chr19 52554235 N chr19 52555242 N DUP 5
SRR1766442.18587917 chr19 52554836 N chr19 52555341 N DEL 5
SRR1766471.1843198 chr19 52554578 N chr19 52555419 N DEL 1
SRR1766442.5276965 chr19 52554156 N chr19 52555583 N DUP 5
SRR1766471.11844205 chr22 47159175 N chr22 47159479 N DUP 7
SRR1766459.2164937 chr10 2374441 N chr10 2374574 N DUP 2
SRR1766442.31280042 chr5 40697200 N chr5 40697301 N DEL 2
SRR1766459.8336534 chr5 40697200 N chr5 40697301 N DEL 12
SRR1766479.99536 chr5 40697251 N chr5 40697306 N DUP 10
SRR1766443.9554326 chr5 40697251 N chr5 40697306 N DUP 10
SRR1766442.31258665 chr5 40697251 N chr5 40697306 N DUP 10
SRR1766467.8179777 chr5 40697251 N chr5 40697306 N DUP 10
SRR1766468.1900450 chr5 40697200 N chr5 40697301 N DEL 50
SRR1766460.5875149 chr5 40697200 N chr5 40697301 N DEL 50
SRR1766477.8398286 chr5 40697252 N chr5 40697307 N DUP 10
SRR1766472.9836874 chr5 40697278 N chr5 40697416 N DEL 3
SRR1766443.7104018 chr5 40697222 N chr5 40697420 N DEL 3
SRR1766484.11099372 chr5 169613851 N chr5 169613938 N DEL 1
SRR1766443.9356434 chr5 169613851 N chr5 169613934 N DEL 5
SRR1766472.3453397 chr5 169613850 N chr5 169613935 N DEL 4
SRR1766477.3311831 chr5 169613850 N chr5 169613937 N DEL 2
SRR1766481.3959264 chr10 26811885 N chr10 26811940 N DEL 7
SRR1766451.8094159 chr10 26811885 N chr10 26811940 N DEL 9
SRR1766442.25115702 chr10 26811885 N chr10 26811940 N DEL 9
SRR1766478.870281 chr10 26811898 N chr10 26811953 N DEL 2
SRR1766459.4474013 chr10 26811890 N chr10 26811945 N DEL 10
SRR1766460.9439543 chr10 26811890 N chr10 26811945 N DEL 10
SRR1766446.2690642 chr16 5488832 N chr16 5488951 N DUP 5
SRR1766472.8613193 chr16 5488875 N chr16 5488994 N DUP 5
SRR1766466.4984554 chr16 5488875 N chr16 5488994 N DUP 5
SRR1766480.2494670 chr16 5488879 N chr16 5488998 N DUP 5
SRR1766442.27210841 chr16 5488884 N chr16 5489003 N DUP 5
SRR1766478.10921560 chr16 5488771 N chr16 5488888 N DEL 2
SRR1766461.10189136 chr16 5488839 N chr16 5488960 N DEL 7
SRR1766448.4905658 chr9 43326680 N chr9 43327112 N DUP 1
SRR1766465.7092193 chr9 43326829 N chr9 43326903 N DUP 5
SRR1766480.2163447 chr9 43326669 N chr9 43326949 N DUP 3
SRR1766475.7417461 chr9 43326702 N chr9 43326951 N DEL 11
SRR1766462.6094011 chr19 37527331 N chr19 37527439 N DEL 7
SRR1766482.12406343 chr22 45291682 N chr22 45291834 N DUP 5
SRR1766461.1174252 chr22 45291462 N chr22 45291824 N DUP 6
SRR1766472.75379 chr22 45291815 N chr22 45292039 N DEL 5
SRR1766461.9062330 chr22 45291815 N chr22 45292039 N DEL 5
SRR1766475.5334340 chr22 45291480 N chr22 45291803 N DEL 5
SRR1766449.7864286 chr22 45291480 N chr22 45291900 N DEL 5
SRR1766450.790767 chr22 45291605 N chr22 45291944 N DEL 5
SRR1766455.3193400 chr22 45291743 N chr22 45292015 N DEL 6
SRR1766462.3222562 chr22 45291780 N chr22 45292052 N DEL 6
SRR1766457.1457189 chr22 45291824 N chr22 45292096 N DEL 5
SRR1766451.9390055 chr6 1054136 N chr6 1054188 N DUP 16
SRR1766453.750168 chr6 1054124 N chr6 1054177 N DUP 23
SRR1766476.11291175 chr17 15166151 N chr17 15166215 N DUP 8
SRR1766450.4982321 chr17 15166166 N chr17 15166232 N DEL 4
SRR1766484.2791278 chr17 15166167 N chr17 15166233 N DEL 3
SRR1766485.8927584 chr22 48757288 N chr22 48757406 N DEL 5
SRR1766451.5238599 chr22 48757307 N chr22 48757461 N DEL 2
SRR1766442.32708715 chr22 48757409 N chr22 48757482 N DEL 1
SRR1766460.8742278 chr22 48757389 N chr22 48757530 N DEL 5
SRR1766442.8735881 chr22 48757304 N chr22 48757589 N DUP 31
SRR1766479.10879454 chr22 48757389 N chr22 48757530 N DEL 5
SRR1766448.7457421 chr22 48757389 N chr22 48757528 N DUP 8
SRR1766453.9027704 chr22 48757290 N chr22 48757507 N DUP 12
SRR1766485.7566056 chr22 48757461 N chr22 48757593 N DUP 32
SRR1766445.9601123 chr22 48757462 N chr22 48757594 N DUP 32
SRR1766470.9224590 chr22 48757461 N chr22 48757593 N DUP 32
SRR1766482.9063439 chr22 48757314 N chr22 48757380 N DEL 8
SRR1766450.387174 chr22 48757463 N chr22 48757566 N DUP 17
SRR1766463.9759456 chr22 48757461 N chr22 48757593 N DUP 27
SRR1766447.6359185 chr22 48757423 N chr22 48757562 N DUP 5
SRR1766458.6284656 chr22 48757304 N chr22 48757482 N DUP 10
SRR1766468.3496635 chr22 48757314 N chr22 48757432 N DEL 5
SRR1766450.234388 chr22 48757304 N chr22 48757508 N DUP 21
SRR1766476.3236244 chr22 48757482 N chr22 48757549 N DUP 15
SRR1766451.7704511 chr22 48757482 N chr22 48757549 N DUP 15
SRR1766478.11778193 chr22 48757304 N chr22 48757446 N DUP 23
SRR1766483.9939486 chr22 48757482 N chr22 48757588 N DUP 10
SRR1766464.5258628 chr13 97949752 N chr13 97949887 N DEL 4
SRR1766479.12313687 chr13 97949770 N chr13 97949905 N DEL 5
SRR1766442.12723009 chr1 55662714 N chr1 55662790 N DUP 10
SRR1766482.8429665 chr1 55662714 N chr1 55662790 N DUP 11
SRR1766467.9973048 chr1 55662714 N chr1 55662790 N DUP 17
SRR1766462.4756125 chr1 55662693 N chr1 55662814 N DUP 9
SRR1766463.7141646 chr1 55662693 N chr1 55662814 N DUP 9
SRR1766484.12197963 chr1 55662693 N chr1 55662814 N DUP 9
SRR1766445.11000 chr8 93833401 N chr8 93833555 N DEL 1
SRR1766481.11856407 chr8 93833413 N chr8 93834274 N DEL 5
SRR1766471.415555 chr8 93833420 N chr8 93833802 N DEL 10
SRR1766483.8067136 chr8 93833434 N chr8 93834000 N DEL 9
SRR1766461.2663755 chr8 93833450 N chr8 93834016 N DEL 8
SRR1766476.11267475 chr8 93833416 N chr8 93833798 N DEL 19
SRR1766479.9870115 chr8 93833430 N chr8 93834628 N DEL 5
SRR1766467.1453960 chr8 93833460 N chr8 93833655 N DEL 4
SRR1766469.4498363 chr8 93833457 N chr8 93833802 N DEL 11
SRR1766442.31761761 chr8 93833474 N chr8 93833743 N DEL 1
SRR1766467.1500862 chr8 93833647 N chr8 93834531 N DEL 5
SRR1766454.9765982 chr8 93833623 N chr8 93834032 N DEL 5
SRR1766454.10964289 chr8 93833648 N chr8 93834241 N DEL 5
SRR1766454.10260786 chr8 93833694 N chr8 93833808 N DEL 10
SRR1766457.2251652 chr8 93833486 N chr8 93833605 N DEL 3
SRR1766457.6028421 chr8 93833486 N chr8 93833605 N DEL 3
SRR1766446.9710512 chr8 93833664 N chr8 93833999 N DEL 20
SRR1766454.6077255 chr8 93833697 N chr8 93833774 N DEL 5
SRR1766473.194906 chr8 93833772 N chr8 93833918 N DEL 5
SRR1766457.2120505 chr8 93833788 N chr8 93834010 N DEL 15
SRR1766457.5092573 chr8 93833797 N chr8 93834019 N DEL 5
SRR1766442.12588855 chr8 93833857 N chr8 93834409 N DEL 10
SRR1766465.795812 chr8 93833864 N chr8 93834416 N DEL 5
SRR1766447.5158641 chr8 93833866 N chr8 93834164 N DEL 5
SRR1766449.2446602 chr8 93833526 N chr8 93833794 N DEL 5
SRR1766451.983111 chr8 93833578 N chr8 93833807 N DEL 1
SRR1766485.3591504 chr8 93833820 N chr8 93834040 N DUP 5
SRR1766451.7106615 chr8 93833820 N chr8 93834040 N DUP 5
SRR1766466.10890946 chr8 93833820 N chr8 93834040 N DUP 5
SRR1766462.3975082 chr8 93833820 N chr8 93834040 N DUP 5
SRR1766482.137107 chr8 93833827 N chr8 93834047 N DUP 5
SRR1766475.2863457 chr8 93833976 N chr8 93834127 N DEL 3
SRR1766448.393606 chr8 93833981 N chr8 93834494 N DEL 5
SRR1766476.5263881 chr8 93833673 N chr8 93834008 N DEL 5
SRR1766444.4475118 chr8 93833718 N chr8 93834053 N DEL 17
SRR1766465.7612498 chr8 93834172 N chr8 93834498 N DEL 1
SRR1766462.3975082 chr8 93833417 N chr8 93834133 N DEL 5
SRR1766454.6077255 chr8 93833481 N chr8 93834160 N DEL 5
SRR1766466.5276754 chr8 93833894 N chr8 93834298 N DUP 5
SRR1766486.1994123 chr8 93833484 N chr8 93834234 N DEL 5
SRR1766475.11039084 chr8 93834128 N chr8 93834237 N DEL 2
SRR1766455.9077632 chr8 93833770 N chr8 93834252 N DEL 9
SRR1766460.4721376 chr8 93833890 N chr8 93834367 N DUP 1
SRR1766455.8497392 chr8 93834003 N chr8 93834370 N DUP 5
SRR1766463.5269019 chr8 93834284 N chr8 93834537 N DUP 5
SRR1766443.570601 chr8 93834031 N chr8 93834290 N DEL 8
SRR1766486.3691980 chr8 93833815 N chr8 93834295 N DEL 5
SRR1766485.2070842 chr8 93833481 N chr8 93834378 N DEL 3
SRR1766481.6907198 chr8 93833466 N chr8 93834505 N DUP 2
SRR1766465.1330118 chr8 93833900 N chr8 93834415 N DEL 4
SRR1766463.9926302 chr8 93834036 N chr8 93834441 N DEL 6
SRR1766478.7566217 chr8 93834418 N chr8 93834525 N DUP 11
SRR1766442.20731211 chr8 93834552 N chr8 93834670 N DEL 5
SRR1766452.4334828 chr8 93834033 N chr8 93834587 N DUP 5
SRR1766475.9845028 chr8 93834161 N chr8 93834524 N DEL 5
SRR1766471.8097515 chr8 93834171 N chr8 93834534 N DEL 5
SRR1766445.2625664 chr8 93834566 N chr8 93834645 N DUP 10
SRR1766468.6068525 chr8 93834558 N chr8 93834637 N DUP 5
SRR1766450.294347 chr8 93834558 N chr8 93834637 N DUP 5
SRR1766475.6150782 chr8 93834558 N chr8 93834637 N DUP 5
SRR1766445.7694183 chr8 93834558 N chr8 93834637 N DUP 5
SRR1766465.5009357 chr8 93834558 N chr8 93834637 N DUP 5
SRR1766446.2111625 chr8 93834558 N chr8 93834637 N DUP 5
SRR1766471.3274525 chr8 93834558 N chr8 93834637 N DUP 5
SRR1766471.6076670 chr8 93833445 N chr8 93834563 N DEL 5
SRR1766478.6747538 chr8 93834691 N chr8 93834883 N DEL 10
SRR1766442.13569260 chr8 93834718 N chr8 93834833 N DEL 16
SRR1766444.5612100 chr8 93833458 N chr8 93834768 N DUP 5
SRR1766467.11908307 chr8 93834432 N chr8 93834698 N DEL 9
SRR1766466.7674599 chr8 93833765 N chr8 93834883 N DEL 5
SRR1766479.11995470 chr8 93833420 N chr8 93834920 N DEL 5
SRR1766486.3006690 chr8 93834270 N chr8 93834949 N DEL 5
SRR1766474.1756665 chr19 50371787 N chr19 50371950 N DUP 9
SRR1766467.157147 chr18 29511747 N chr18 29511837 N DUP 5
SRR1766458.652419 chr18 29511747 N chr18 29511837 N DUP 5
SRR1766477.4940416 chr18 29511747 N chr18 29511837 N DUP 5
SRR1766474.2693825 chr18 29511747 N chr18 29511837 N DUP 5
SRR1766442.41957640 chr18 29511747 N chr18 29511837 N DUP 5
SRR1766478.5352112 chr18 29511747 N chr18 29511837 N DUP 5
SRR1766478.11142125 chr18 29511662 N chr18 29511838 N DEL 15
SRR1766476.7549764 chr18 29511662 N chr18 29511838 N DEL 12
SRR1766461.6612637 chr18 29511763 N chr18 29511881 N DEL 5
SRR1766442.27394378 chr18 29511893 N chr18 29511946 N DEL 22
SRR1766443.10079627 chr18 29511893 N chr18 29511946 N DEL 21
SRR1766464.7102646 chr18 29512113 N chr18 29512280 N DEL 1
SRR1766450.9517795 chr18 29512113 N chr18 29512280 N DEL 2
SRR1766449.2930437 chr18 29512100 N chr18 29512173 N DUP 7
SRR1766479.6730721 chr18 29512100 N chr18 29512173 N DUP 7
SRR1766458.8548974 chr18 29511918 N chr18 29512186 N DUP 5
SRR1766484.5172379 chr18 29511787 N chr18 29512116 N DEL 12
SRR1766476.2134445 chr18 29511761 N chr18 29512116 N DEL 12
SRR1766447.730327 chr18 29512116 N chr18 29512199 N DUP 22
SRR1766442.3639045 chr18 29511761 N chr18 29512116 N DEL 11
SRR1766484.3325011 chr18 29511761 N chr18 29512116 N DEL 8
SRR1766486.6897880 chr18 29512102 N chr18 29512175 N DUP 20
SRR1766451.10200674 chr18 29512116 N chr18 29512199 N DUP 29
SRR1766455.7116177 chr18 29512204 N chr18 29512344 N DUP 13
SRR1766467.292615 chr18 29512204 N chr18 29512344 N DUP 14
SRR1766476.1767158 chr18 29512133 N chr18 29512346 N DUP 21
SRR1766481.2297823 chr18 29512133 N chr18 29512346 N DUP 21
SRR1766442.28760933 chr18 29512204 N chr18 29512344 N DUP 27
SRR1766486.4476584 chr18 29512230 N chr18 29512344 N DUP 25
SRR1766450.1116268 chr18 29511666 N chr18 29512230 N DEL 20
SRR1766479.9912839 chr18 29511666 N chr18 29512230 N DEL 20
SRR1766450.9692300 chr18 29511751 N chr18 29512205 N DEL 12
SRR1766466.1942525 chr18 29511666 N chr18 29512204 N DEL 14
SRR1766475.5918332 chr18 29511666 N chr18 29512204 N DEL 18
SRR1766442.8245711 chr18 29511666 N chr18 29512230 N DEL 20
SRR1766469.3902827 chr18 29511666 N chr18 29512230 N DEL 20
SRR1766443.10089516 chr18 29511662 N chr18 29511838 N DEL 5
SRR1766485.12004081 chr18 29511666 N chr18 29512230 N DEL 14
SRR1766448.7994307 chr18 29511608 N chr18 29512243 N DEL 2
SRR1766481.11859953 chr18 29512199 N chr18 29512282 N DEL 26
SRR1766442.44756759 chr18 29512163 N chr18 29512282 N DEL 28
SRR1766454.325548 chr18 29512230 N chr18 29512344 N DUP 27
SRR1766464.10293517 chr12 53385186 N chr12 53385807 N DEL 4
SRR1766476.3860179 chr12 53385175 N chr12 53385794 N DUP 7
SRR1766457.5715172 chr12 53385561 N chr12 53385881 N DEL 5
SRR1766442.40295938 chr12 53385730 N chr12 53386049 N DEL 1
SRR1766470.1182425 chr12 53385171 N chr12 53385790 N DUP 1
SRR1766461.3529355 chr12 53385293 N chr12 53385912 N DEL 5
SRR1766473.6123300 chr12 53385634 N chr12 53385953 N DEL 5
SRR1766453.5330784 chr12 53385642 N chr12 53385961 N DEL 9
SRR1766442.42093179 chr4 162764161 N chr4 162764228 N DUP 22
SRR1766445.10545933 chr4 162764161 N chr4 162764228 N DUP 28
SRR1766446.4231808 chr4 162764120 N chr4 162764228 N DUP 30
SRR1766484.9703071 chr4 162764120 N chr4 162764228 N DUP 30
SRR1766445.6231410 chr4 162764160 N chr4 162764209 N DUP 37
SRR1766466.3922666 chr4 162764120 N chr4 162764228 N DUP 24
SRR1766476.10399494 chr4 162764120 N chr4 162764228 N DUP 24
SRR1766465.7415466 chr4 162764120 N chr4 162764228 N DUP 29
SRR1766476.10864049 chr4 162764120 N chr4 162764228 N DUP 29
SRR1766468.575116 chr4 162764160 N chr4 162764209 N DUP 34
SRR1766456.5541965 chr4 162764160 N chr4 162764209 N DUP 36
SRR1766464.10343395 chr4 162764160 N chr4 162764209 N DUP 36
SRR1766483.5105017 chr4 162764143 N chr4 162764201 N DEL 23
SRR1766446.4776360 chr4 162764143 N chr4 162764201 N DEL 21
SRR1766477.9642725 chr4 162764143 N chr4 162764201 N DEL 21
SRR1766462.59031 chr4 162764143 N chr4 162764201 N DEL 21
SRR1766484.9098791 chr4 162764116 N chr4 162764199 N DEL 12
SRR1766443.1572423 chr4 162764143 N chr4 162764201 N DEL 23
SRR1766456.815454 chr4 162764125 N chr4 162764199 N DEL 14
SRR1766455.7585734 chr4 162764143 N chr4 162764201 N DEL 23
SRR1766447.7595681 chr4 162764125 N chr4 162764199 N DEL 14
SRR1766479.3682614 chr4 162764115 N chr4 162764207 N DEL 9
SRR1766479.4210118 chr4 162764118 N chr4 162764210 N DEL 6
SRR1766482.2426197 chr4 162764122 N chr4 162764214 N DEL 2
SRR1766462.297208 chr4 162764116 N chr4 162764208 N DEL 8
SRR1766481.12441686 chr4 162764116 N chr4 162764208 N DEL 8
SRR1766471.4590922 chr7 73509087 N chr7 73509397 N DEL 3
SRR1766452.740028 chr7 73509058 N chr7 73509368 N DEL 5
SRR1766465.246786 chr14 67700822 N chr14 67701132 N DEL 4
SRR1766476.10614659 chr14 67700855 N chr14 67701166 N DEL 5
SRR1766470.9437047 chr14 67700868 N chr14 67701174 N DEL 11
SRR1766478.1303720 chr14 67700618 N chr14 67700928 N DEL 5
SRR1766480.6959696 chr2 70107363 N chr2 70107431 N DUP 2
SRR1766480.878275 chr10 68503004 N chr10 68503089 N DEL 12
SRR1766480.2338559 chr10 68502982 N chr10 68503105 N DEL 3
SRR1766483.6900094 chr5 474337 N chr5 474440 N DEL 7
SRR1766463.4421973 chr5 474440 N chr5 474640 N DUP 2
SRR1766458.2057405 chr6 994146 N chr6 994210 N DUP 1
SRR1766461.10562237 chr6 994146 N chr6 994210 N DUP 10
SRR1766443.559355 chr7 157324342 N chr7 157324674 N DUP 5
SRR1766477.3807290 chr7 157324688 N chr7 157325000 N DEL 5
SRR1766484.10722071 chr7 157324644 N chr7 157324954 N DUP 1
SRR1766449.7080122 chr7 157324630 N chr7 157324940 N DUP 5
SRR1766478.6980619 chr7 157324657 N chr7 157324967 N DUP 2
SRR1766454.9100429 chr7 157324657 N chr7 157324967 N DUP 5
SRR1766451.4652891 chr7 157324682 N chr7 157324994 N DEL 5
SRR1766460.10152860 chr7 157324682 N chr7 157324994 N DEL 5
SRR1766473.7978047 chr7 157324697 N chr7 157325009 N DEL 15
SRR1766464.2574685 chr7 157324696 N chr7 157325008 N DEL 5
SRR1766452.806529 chr7 157324675 N chr7 157324987 N DEL 5
SRR1766442.13136366 chr7 157324697 N chr7 157325009 N DEL 10
SRR1766483.5680166 chr7 157324702 N chr7 157325014 N DEL 5
SRR1766464.561889 chr7 157324385 N chr7 157325030 N DEL 12
SRR1766462.5228266 chr7 157324692 N chr7 157325004 N DEL 4
SRR1766442.33744957 chr20 64105723 N chr20 64105875 N DEL 20
SRR1766483.9561670 chr20 64105722 N chr20 64105874 N DEL 20
SRR1766461.8523351 chr20 64105722 N chr20 64105874 N DEL 20
SRR1766468.5538195 chr20 64105681 N chr20 64105875 N DEL 20
SRR1766477.6259834 chr3 188179144 N chr3 188179197 N DUP 6
SRR1766468.5475635 chr3 188179159 N chr3 188179258 N DEL 1
SRR1766483.8244552 chr14 34735123 N chr14 34735250 N DEL 11
SRR1766467.1220833 chr14 34735115 N chr14 34735256 N DEL 5
SRR1766471.5447847 chr14 34735116 N chr14 34735259 N DEL 9
SRR1766453.10892011 chr14 34735123 N chr14 34735288 N DEL 11
SRR1766457.3754226 chr14 34735116 N chr14 34735273 N DEL 7
SRR1766466.4769805 chr14 34735113 N chr14 34735274 N DEL 5
SRR1766442.8429989 chr14 34735237 N chr14 34735298 N DEL 5
SRR1766482.12340820 chr14 34735114 N chr14 34735299 N DEL 4
SRR1766452.2675250 chr14 34735106 N chr14 34735315 N DEL 6
SRR1766450.9148354 chr9 134523988 N chr9 134524247 N DUP 6
SRR1766471.7665878 chr9 134523986 N chr9 134524185 N DUP 5
SRR1766450.9702322 chr9 134523967 N chr9 134524038 N DEL 5
SRR1766448.1616070 chr9 134523935 N chr9 134524194 N DUP 5
SRR1766457.9320523 chr9 134523932 N chr9 134524191 N DUP 5
SRR1766480.1702292 chr9 134524046 N chr9 134524175 N DUP 10
SRR1766479.7397739 chr9 134524128 N chr9 134524187 N DUP 10
SRR1766445.6411802 chr9 134523932 N chr9 134524191 N DUP 10
SRR1766463.94800 chr9 134524146 N chr9 134524205 N DUP 5
SRR1766461.279125 chr9 134524128 N chr9 134524187 N DUP 5
SRR1766454.636191 chr9 134524146 N chr9 134524205 N DUP 5
SRR1766453.4178465 chr6 522335 N chr6 522533 N DEL 5
SRR1766466.6111114 chr6 522354 N chr6 522748 N DEL 15
SRR1766470.11179145 chr6 522464 N chr6 522564 N DEL 1
SRR1766455.8439651 chr6 522586 N chr6 522685 N DEL 1
SRR1766447.2393390 chr6 522549 N chr6 522842 N DUP 2
SRR1766464.1432952 chr6 522376 N chr6 522770 N DEL 6
SRR1766445.656603 chr6 522428 N chr6 522822 N DEL 4
SRR1766480.3745003 chr12 58320336 N chr12 58320437 N DUP 7
SRR1766451.398276 chr12 58320336 N chr12 58320437 N DUP 7
SRR1766467.6109314 chr13 113375287 N chr13 113375528 N DEL 5
SRR1766486.9232122 chr13 113375300 N chr13 113375981 N DEL 10
SRR1766442.16716254 chr13 113375340 N chr13 113376001 N DEL 10
SRR1766459.3527291 chr13 113375263 N chr13 113375352 N DUP 5
SRR1766484.6218978 chr13 113375303 N chr13 113375624 N DEL 5
SRR1766466.8833002 chr13 113375420 N chr13 113376001 N DEL 10
SRR1766453.1685489 chr13 113375367 N chr13 113375608 N DEL 10
SRR1766442.18034647 chr13 113375420 N chr13 113376001 N DEL 10
SRR1766452.8786077 chr13 113375360 N chr13 113375681 N DEL 5
SRR1766485.3821950 chr13 113375382 N chr13 113375623 N DEL 5
SRR1766483.1007781 chr13 113375420 N chr13 113376001 N DEL 10
SRR1766465.3232313 chr13 113375519 N chr13 113375918 N DUP 5
SRR1766467.9101855 chr13 113375367 N chr13 113375926 N DUP 5
SRR1766469.7187815 chr13 113375533 N chr13 113375932 N DUP 1
SRR1766477.2345401 chr13 113375519 N chr13 113375918 N DUP 5
SRR1766458.824786 chr13 113375289 N chr13 113375598 N DUP 16
SRR1766474.9347228 chr13 113375599 N chr13 113375918 N DUP 5
SRR1766463.8563728 chr13 113375602 N chr13 113375921 N DUP 10
SRR1766482.12157498 chr13 113375580 N chr13 113376001 N DEL 5
SRR1766467.6109314 chr13 113375282 N chr13 113375613 N DEL 1
SRR1766444.2461363 chr13 113375679 N chr13 113375918 N DUP 5
SRR1766443.1149995 chr13 113375679 N chr13 113375918 N DUP 5
SRR1766471.340189 chr13 113375528 N chr13 113375927 N DUP 5
SRR1766444.2461363 chr13 113375529 N chr13 113375928 N DUP 5
SRR1766442.7748246 chr13 113376001 N chr13 113376080 N DUP 15
SRR1766473.5647016 chr13 113376001 N chr13 113376080 N DUP 15
SRR1766446.8369414 chr13 113375580 N chr13 113376001 N DEL 10
SRR1766442.593321 chr13 113375740 N chr13 113376001 N DEL 4
SRR1766475.8314229 chr13 113375529 N chr13 113375850 N DEL 5
SRR1766474.9347228 chr13 113375839 N chr13 113375918 N DUP 5
SRR1766459.3527291 chr13 113375849 N chr13 113375928 N DUP 5
SRR1766463.8786286 chr13 113375839 N chr13 113375998 N DUP 15
SRR1766473.9224426 chr13 113375525 N chr13 113375846 N DEL 5
SRR1766482.9950323 chr13 113375839 N chr13 113375918 N DUP 5
SRR1766474.4980775 chr13 113375839 N chr13 113375918 N DUP 5
SRR1766448.6773321 chr13 113375327 N chr13 113375966 N DUP 5
SRR1766466.8833002 chr13 113375357 N chr13 113375918 N DEL 5
SRR1766477.276055 chr13 113375706 N chr13 113375947 N DEL 5
SRR1766458.824786 chr13 113375337 N chr13 113375958 N DEL 13
SRR1766461.5918936 chr13 113375679 N chr13 113376018 N DUP 5
SRR1766486.9232122 chr13 113375839 N chr13 113376018 N DUP 5
SRR1766476.1778747 chr13 113375839 N chr13 113376018 N DUP 5
SRR1766483.1007781 chr13 113375341 N chr13 113376082 N DEL 5
SRR1766467.2006353 chr13 113375997 N chr13 113376138 N DEL 6
SRR1766477.730531 chr13 113375969 N chr13 113376257 N DUP 5
SRR1766448.3891786 chr13 113376174 N chr13 113376400 N DUP 5
SRR1766475.10405569 chr13 113375370 N chr13 113376250 N DEL 5
SRR1766452.381912 chr13 113376041 N chr13 113376349 N DEL 10
SRR1766485.10171440 chr2 68012916 N chr2 68013033 N DEL 5
SRR1766452.5403440 chr12 2177645 N chr12 2177714 N DUP 2
SRR1766460.5768967 chr6 71316412 N chr6 71316473 N DUP 10
SRR1766476.5189228 chr6 71316412 N chr6 71316473 N DUP 10
SRR1766444.5008869 chr18 3113361 N chr18 3113452 N DUP 5
SRR1766455.7317657 chr18 3113361 N chr18 3113452 N DUP 5
SRR1766483.1945455 chr18 3113373 N chr18 3113486 N DEL 15
SRR1766468.2567035 chr18 3113359 N chr18 3113492 N DEL 6
SRR1766482.12819358 chr3 77323092 N chr3 77323144 N DUP 14
SRR1766470.5413413 chr3 77323092 N chr3 77323144 N DUP 10
SRR1766482.5469074 chr3 77323092 N chr3 77323173 N DUP 20
SRR1766481.4646853 chr3 77323092 N chr3 77323231 N DUP 5
SRR1766475.3383508 chr3 77323092 N chr3 77323231 N DUP 14
SRR1766460.8179183 chr3 77323072 N chr3 77323153 N DUP 10
SRR1766452.10560426 chr3 77323092 N chr3 77323202 N DUP 8
SRR1766453.6593551 chr3 77323092 N chr3 77323144 N DUP 14
SRR1766478.4434323 chr3 77323092 N chr3 77323202 N DUP 10
SRR1766475.10073472 chr3 77323094 N chr3 77323146 N DUP 10
SRR1766480.1027218 chr3 77323092 N chr3 77323144 N DUP 12
SRR1766465.6317734 chr3 77323072 N chr3 77323211 N DUP 10
SRR1766464.7925165 chr3 77323092 N chr3 77323231 N DUP 12
SRR1766475.1021030 chr3 77323092 N chr3 77323144 N DUP 18
SRR1766459.1207565 chr3 77323068 N chr3 77323236 N DUP 12
SRR1766450.6971141 chr3 77323094 N chr3 77323204 N DUP 12
SRR1766445.2207246 chr3 77322920 N chr3 77323076 N DEL 2
SRR1766475.7501766 chr3 77323068 N chr3 77323236 N DUP 13
SRR1766478.2237840 chr3 77323078 N chr3 77323227 N DUP 7
SRR1766474.6846091 chr3 77323097 N chr3 77323219 N DEL 5
SRR1766479.8293449 chr3 77323097 N chr3 77323219 N DEL 5
SRR1766468.3098755 chr3 77322918 N chr3 77323219 N DEL 5
SRR1766480.4069988 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766471.6636310 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766468.7840055 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766480.6578666 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766471.8305279 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766451.7845618 chrY 10790402 N chrY 10790643 N DEL 12
SRR1766447.9381161 chrY 10790347 N chrY 10790667 N DEL 2
SRR1766462.7983021 chrY 10790386 N chrY 10790480 N DUP 30
SRR1766452.2963636 chr2 38479868 N chr2 38480021 N DEL 11
SRR1766479.1095609 chr2 38479874 N chr2 38480031 N DEL 3
SRR1766470.7845645 chr19 14636153 N chr19 14636289 N DUP 4
SRR1766455.3814826 chr19 14636153 N chr19 14636289 N DUP 4
SRR1766446.7143820 chr19 14636153 N chr19 14636289 N DUP 8
SRR1766450.3678986 chr19 14636173 N chr19 14636299 N DEL 15
SRR1766453.9491509 chr19 14636175 N chr19 14636301 N DEL 13
SRR1766466.6225683 chr19 14636176 N chr19 14636302 N DEL 12
SRR1766442.21322860 chr19 14636177 N chr19 14636303 N DEL 11
SRR1766458.5319495 chr19 14636216 N chr19 14636310 N DEL 4
SRR1766479.8754798 chr19 14636216 N chr19 14636310 N DEL 4
SRR1766444.4722992 chr19 14636179 N chr19 14636305 N DEL 9
SRR1766474.2218712 chr18 22740454 N chr18 22740521 N DUP 46
SRR1766472.2340108 chr18 22740454 N chr18 22740521 N DUP 46
SRR1766467.9015539 chr18 22740454 N chr18 22740521 N DUP 46
SRR1766476.2570549 chr18 22740477 N chr18 22740571 N DUP 11
SRR1766461.3979564 chr18 22740477 N chr18 22740571 N DUP 12
SRR1766470.11076688 chr18 22740478 N chr18 22740572 N DUP 11
SRR1766479.7642685 chr18 22740480 N chr18 22740574 N DUP 13
SRR1766447.3482777 chr12 7197438 N chr12 7197611 N DUP 3
SRR1766469.4024029 chr12 7197464 N chr12 7197615 N DUP 9
SRR1766479.13293243 chr12 7197426 N chr12 7197528 N DUP 12
SRR1766444.4710132 chr12 7197426 N chr12 7197528 N DUP 12
SRR1766453.3652266 chr12 7197426 N chr12 7197528 N DUP 17
SRR1766446.10526335 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766486.8071106 chr12 7197426 N chr12 7197528 N DUP 20
SRR1766478.5771996 chr12 7197490 N chr12 7197541 N DUP 10
SRR1766442.17743676 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766467.8277990 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766483.7669952 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766483.7090183 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766464.2949238 chr12 7197464 N chr12 7197517 N DUP 22
SRR1766462.11102186 chr12 7197464 N chr12 7197544 N DUP 27
SRR1766486.11792641 chr12 7197427 N chr12 7197580 N DUP 23
SRR1766478.3221258 chr12 7197427 N chr12 7197580 N DUP 28
SRR1766459.6053149 chr12 7197464 N chr12 7197544 N DUP 27
SRR1766460.4289330 chr12 7197484 N chr12 7197563 N DUP 28
SRR1766457.550630 chr12 7197464 N chr12 7197570 N DUP 31
SRR1766479.5202926 chr12 7197464 N chr12 7197570 N DUP 31
SRR1766484.5798433 chr12 7197515 N chr12 7197588 N DUP 11
SRR1766474.10345640 chr12 7197523 N chr12 7197575 N DEL 8
SRR1766457.550630 chr12 7197523 N chr12 7197575 N DEL 8
SRR1766454.10278459 chr12 7197471 N chr12 7197649 N DUP 5
SRR1766467.8998667 chr12 7197482 N chr12 7197564 N DUP 25
SRR1766465.7470978 chr12 7197523 N chr12 7197575 N DEL 5
SRR1766475.7449761 chr12 7197454 N chr12 7197582 N DEL 11
SRR1766454.6180553 chr12 7197454 N chr12 7197582 N DEL 10
SRR1766449.8470532 chr12 7197454 N chr12 7197582 N DEL 10
SRR1766442.34667529 chr12 7197592 N chr12 7197690 N DUP 5
SRR1766485.7670183 chr4 3362782 N chr4 3362951 N DUP 5
SRR1766466.6367117 chr4 3362782 N chr4 3362951 N DUP 5
SRR1766485.2364746 chr18 21577177 N chr18 21577804 N DEL 1
SRR1766448.769230 chr18 21577158 N chr18 21577784 N DUP 5
SRR1766470.4351337 chr10 82098397 N chr10 82098473 N DEL 13
SRR1766449.1348248 chr10 82098400 N chr10 82098476 N DEL 12
SRR1766454.2598736 chr1 167806412 N chr1 167806567 N DEL 5
SRR1766464.6310723 chr1 167806409 N chr1 167806641 N DEL 5
SRR1766470.6383648 chr1 167806422 N chr1 167806500 N DEL 1
SRR1766442.23965795 chr1 167806422 N chr1 167806500 N DEL 1
SRR1766461.4992520 chr1 167806422 N chr1 167806500 N DEL 5
SRR1766455.151795 chr1 167806422 N chr1 167806500 N DEL 5
SRR1766463.10800530 chr1 167806412 N chr1 167806490 N DEL 5
SRR1766453.2639819 chr1 167806412 N chr1 167806490 N DEL 10
SRR1766445.5225586 chr1 167806422 N chr1 167806500 N DEL 5
SRR1766453.3175698 chr1 167806422 N chr1 167806500 N DEL 5
SRR1766460.2660085 chr1 167806422 N chr1 167806500 N DEL 5
SRR1766452.449035 chr1 167806422 N chr1 167806500 N DEL 5
SRR1766449.10448864 chr1 167806422 N chr1 167806500 N DEL 5
SRR1766473.4912186 chr1 167806409 N chr1 167806487 N DEL 10
SRR1766477.605377 chr1 167806422 N chr1 167806500 N DEL 5
SRR1766477.9812848 chr1 167806454 N chr1 167806530 N DUP 5
SRR1766452.5863141 chr1 167806460 N chr1 167806536 N DUP 4
SRR1766461.4710836 chr1 167806423 N chr1 167806576 N DUP 2
SRR1766442.17793730 chr1 167806497 N chr1 167806575 N DEL 5
SRR1766448.57472 chr1 167806497 N chr1 167806575 N DEL 5
SRR1766454.2598736 chr1 167806497 N chr1 167806575 N DEL 5
SRR1766453.2639819 chr1 167806497 N chr1 167806575 N DEL 5
SRR1766471.5388906 chr1 167806497 N chr1 167806575 N DEL 5
SRR1766475.6425172 chr1 167806448 N chr1 167806603 N DEL 5
SRR1766473.4912186 chr1 167806448 N chr1 167806603 N DEL 5
SRR1766481.8633892 chr1 167806448 N chr1 167806603 N DEL 5
SRR1766454.1615089 chr1 167806458 N chr1 167806613 N DEL 5
SRR1766442.3191675 chr1 167806435 N chr1 167806743 N DEL 1
SRR1766479.2708904 chrX 1581657 N chrX 1582003 N DEL 1
SRR1766448.5642393 chrX 1581740 N chrX 1581880 N DEL 5
SRR1766457.7969891 chrX 1581712 N chrX 1582062 N DEL 5
SRR1766445.2601244 chrX 1581645 N chrX 1581718 N DEL 5
SRR1766450.2462552 chrX 1581852 N chrX 1582057 N DUP 14
SRR1766464.7355476 chrX 1581853 N chrX 1581991 N DUP 5
SRR1766460.7878058 chrX 1581758 N chrX 1581967 N DUP 1
SRR1766460.3221417 chrX 1581806 N chrX 1581946 N DEL 5
SRR1766445.7645559 chrX 1581852 N chrX 1582057 N DUP 5
SRR1766442.39951709 chrX 1581852 N chrX 1582057 N DUP 7
SRR1766442.28468290 chrX 1581852 N chrX 1582057 N DUP 7
SRR1766451.4256155 chrX 1581852 N chrX 1582057 N DUP 9
SRR1766478.10249118 chrX 1581852 N chrX 1582057 N DUP 9
SRR1766483.10365137 chrX 1581852 N chrX 1582057 N DUP 9
SRR1766482.12541918 chrX 1581852 N chrX 1582057 N DUP 9
SRR1766465.9514419 chrX 1582021 N chrX 1582161 N DEL 9
SRR1766442.28469307 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766462.8568193 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766466.10020583 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766486.8495807 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766462.9075244 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766442.42650235 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766445.4425448 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766479.11555393 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766452.2680434 chrX 1581712 N chrX 1582062 N DEL 9
SRR1766456.2615026 chrX 1581737 N chrX 1582087 N DEL 2
SRR1766466.2064314 chrX 1581640 N chrX 1582062 N DEL 9
SRR1766451.6790877 chrX 1581640 N chrX 1582062 N DEL 9
SRR1766448.5642393 chrX 1581640 N chrX 1582062 N DEL 9
SRR1766486.429408 chrX 1581640 N chrX 1582062 N DEL 9
SRR1766454.5133122 chrX 1581642 N chrX 1582064 N DEL 9
SRR1766460.6086991 chrX 1581644 N chrX 1582066 N DEL 9
SRR1766479.2708904 chrX 1581644 N chrX 1582066 N DEL 9
SRR1766442.13690542 chrX 1581717 N chrX 1582067 N DEL 9
SRR1766483.339772 chrX 1581718 N chrX 1582068 N DEL 9
SRR1766484.4236420 chrX 1581718 N chrX 1582068 N DEL 9
SRR1766443.8897487 chrX 1581719 N chrX 1582069 N DEL 8
SRR1766478.8970075 chrX 1581798 N chrX 1582080 N DEL 5
SRR1766455.6152714 chrX 1581645 N chrX 1582126 N DEL 3
SRR1766477.56560 chrX 1581811 N chrX 1582161 N DEL 5
SRR1766463.5827519 chrX 1581676 N chrX 1582161 N DEL 5
SRR1766483.1927469 chrX 1581687 N chrX 1582172 N DEL 4
SRR1766472.5364005 chrX 1581786 N chrX 1581991 N DUP 2
SRR1766465.4657839 chrX 1581786 N chrX 1581991 N DUP 3
SRR1766452.4859997 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766480.6115145 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766459.10889104 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766472.10460707 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766463.4764536 chrX 1582251 N chrX 1582454 N DUP 1
SRR1766478.7168662 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766462.6916880 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766455.1601781 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766450.6416148 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766469.9336191 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766442.15762121 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766442.4019487 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766455.5042480 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766442.21472712 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766442.28286574 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766485.6479064 chrX 1581811 N chrX 1582361 N DUP 5
SRR1766445.7838684 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766468.1846912 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766460.7878058 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766448.5020950 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766451.738595 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766471.3588677 chrX 1581789 N chrX 1581994 N DUP 5
SRR1766483.10446028 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766475.1991190 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766442.21999361 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766442.28469307 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766446.8722417 chrX 1581786 N chrX 1581991 N DUP 5
SRR1766486.7058298 chrX 1582161 N chrX 1582362 N DUP 5
SRR1766454.1017545 chrX 1582161 N chrX 1582362 N DUP 5
SRR1766475.4943487 chrX 1582161 N chrX 1582362 N DUP 5
SRR1766471.3529461 chrX 1581677 N chrX 1582162 N DEL 10
SRR1766445.6281273 chrX 1582161 N chrX 1582362 N DUP 5
SRR1766474.51499 chrX 1582161 N chrX 1582362 N DUP 5
SRR1766471.11551969 chrX 1581686 N chrX 1582373 N DEL 10
SRR1766442.38534548 chrX 1582034 N chrX 1582376 N DEL 1
SRR1766457.8959440 chrX 1581821 N chrX 1582373 N DEL 5
SRR1766472.10559970 chrX 1581821 N chrX 1582373 N DEL 5
SRR1766464.9383842 chrX 1581821 N chrX 1582373 N DEL 5
SRR1766483.10365137 chrX 1581821 N chrX 1582373 N DEL 5
SRR1766475.772120 chrX 1581821 N chrX 1582373 N DEL 5
SRR1766479.11432521 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766479.10596792 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766456.3219212 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766456.4973337 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766465.9691157 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766462.4018810 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766470.4802638 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766442.39951709 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766482.12541918 chrX 1581686 N chrX 1582373 N DEL 5
SRR1766447.1734778 chrX 1581689 N chrX 1582376 N DEL 5
SRR1766457.7423084 chrX 1581693 N chrX 1582380 N DEL 5
SRR1766458.5033157 chrX 1581697 N chrX 1582384 N DEL 4
SRR1766456.4277990 chrX 1581699 N chrX 1582386 N DEL 2
SRR1766484.9893013 chrX 1581639 N chrX 1582398 N DEL 5
SRR1766460.3327054 chr8 82824891 N chr8 82824962 N DEL 7
SRR1766442.14520520 chr10 2669910 N chr10 2669993 N DEL 3
SRR1766467.8154289 chrX 943209 N chrX 943275 N DUP 5
SRR1766469.11124434 chrX 943283 N chrX 943499 N DUP 5
SRR1766442.35398340 chrX 943215 N chrX 943343 N DEL 6
SRR1766465.6043000 chr16 11499269 N chr16 11499453 N DEL 2
SRR1766456.6043241 chr6 166824827 N chr6 166824926 N DEL 14
SRR1766461.1932987 chr6 166824810 N chr6 166824903 N DEL 15
SRR1766468.2685443 chr6 166824860 N chr6 166824957 N DEL 11
SRR1766475.10985322 chr6 166824795 N chr6 166824860 N DUP 13
SRR1766486.6579404 chr6 166824831 N chr6 166824926 N DEL 22
SRR1766469.44660 chr6 166824926 N chr6 166824989 N DUP 18
SRR1766475.10985322 chr6 166824718 N chr6 166824928 N DEL 7
SRR1766455.901312 chr6 166824834 N chr6 166824967 N DEL 9
SRR1766473.4503709 chr6 166824722 N chr6 166824932 N DEL 5
SRR1766456.6043241 chr6 166824823 N chr6 166824934 N DEL 5
SRR1766461.4567677 chr6 166824769 N chr6 166824938 N DEL 3
SRR1766480.3254381 chr6 166824770 N chr6 166824939 N DEL 2
SRR1766465.4488605 chr6 166824771 N chr6 166824940 N DEL 1
SRR1766479.5464903 chr6 166824776 N chr6 166824967 N DEL 12
SRR1766459.3169022 chr6 166824776 N chr6 166824967 N DEL 12
SRR1766448.2568363 chr6 166824721 N chr6 166824973 N DEL 5
SRR1766456.5674649 chr6 166824721 N chr6 166824973 N DEL 5
SRR1766463.1047278 chr6 166824829 N chr6 166824982 N DEL 5
SRR1766464.6625571 chr6 166824727 N chr6 166824979 N DEL 3
SRR1766444.1809950 chrY 6081086 N chrY 6081407 N DEL 5
SRR1766467.7704282 chrY 6081085 N chrY 6081406 N DEL 21
SRR1766471.4730322 chrY 6081147 N chrY 6081468 N DEL 2
SRR1766486.10503348 chr17 43634060 N chr17 43634113 N DUP 6
SRR1766442.32955485 chr16 904181 N chr16 904320 N DUP 5
SRR1766478.5181105 chr16 904000 N chr16 904323 N DUP 6
SRR1766483.7451286 chr16 904008 N chr16 904331 N DUP 6
SRR1766448.2171547 chr12 132446237 N chr12 132446390 N DEL 5
SRR1766484.157717 chr12 132446223 N chr12 132446374 N DUP 5
SRR1766448.1832658 chr12 132446223 N chr12 132446374 N DUP 5
SRR1766460.8552835 chr12 132446223 N chr12 132446374 N DUP 5
SRR1766467.953269 chr12 132446250 N chr12 132446403 N DEL 2
SRR1766452.6151028 chr3 147778950 N chr3 147779045 N DEL 6
SRR1766479.12059830 chr7 61610310 N chr7 61610822 N DUP 5
SRR1766449.8097491 chr7 61610245 N chr7 61610321 N DEL 5
SRR1766485.7585292 chr7 61610125 N chr7 61610543 N DEL 13
SRR1766479.1141777 chr5 21344703 N chr5 21344773 N DUP 5
SRR1766445.1778680 chr5 21344823 N chr5 21344926 N DEL 5
SRR1766478.9332922 chr5 21344737 N chr5 21344816 N DEL 7
SRR1766454.6379474 chr5 21344829 N chr5 21344912 N DEL 17
SRR1766453.551323 chr5 21344829 N chr5 21344912 N DEL 17
SRR1766449.3101329 chr5 21344829 N chr5 21344912 N DEL 17
SRR1766472.11132225 chrX 375661 N chrX 375758 N DEL 4
SRR1766469.10585343 chrX 375453 N chrX 375692 N DUP 5
SRR1766448.4851324 chr10 16646011 N chr10 16646070 N DUP 8
SRR1766485.4826104 chr10 16646011 N chr10 16646070 N DUP 11
SRR1766477.3528578 chr10 16646011 N chr10 16646070 N DUP 12
SRR1766442.21891090 chr10 16646011 N chr10 16646070 N DUP 15
SRR1766447.10488370 chr10 16646011 N chr10 16646112 N DUP 11
SRR1766448.1342968 chr10 16646011 N chr10 16646112 N DUP 16
SRR1766445.5527388 chr10 16646015 N chr10 16646130 N DUP 8
SRR1766462.772773 chr10 16646072 N chr10 16646129 N DEL 2
SRR1766475.586435 chr10 16646073 N chr10 16646156 N DEL 23
SRR1766464.1106556 chr10 16646073 N chr10 16646156 N DEL 13
SRR1766481.1837505 chr10 14015339 N chr10 14015410 N DEL 9
SRR1766455.6479385 chr10 14015197 N chr10 14015415 N DEL 5
SRR1766470.7827514 chr21 30484466 N chr21 30484537 N DEL 5
SRR1766442.43428699 chr21 30484466 N chr21 30484537 N DEL 5
SRR1766464.8053156 chr21 30484466 N chr21 30484537 N DEL 5
SRR1766450.4709109 chr21 30484469 N chr21 30484540 N DEL 5
SRR1766484.1003446 chr21 30484470 N chr21 30484541 N DEL 5
SRR1766455.5237890 chr21 30484473 N chr21 30484544 N DEL 5
SRR1766455.6479315 chr21 30484473 N chr21 30484544 N DEL 5
SRR1766464.7789299 chr17 77885469 N chr17 77885665 N DEL 10
SRR1766442.4631638 chr17 77885548 N chr17 77885641 N DEL 6
SRR1766461.4281064 chr17 77885458 N chr17 77885692 N DUP 5
SRR1766472.9158598 chr7 158349790 N chr7 158349839 N DUP 5
SRR1766473.3233689 chr7 158349790 N chr7 158349839 N DUP 5
SRR1766442.39731535 chr7 158349790 N chr7 158349839 N DUP 5
SRR1766473.10497524 chr7 158349790 N chr7 158349839 N DUP 5
SRR1766456.429460 chr7 158349790 N chr7 158349839 N DUP 5
SRR1766483.9026879 chr7 158349861 N chr7 158349961 N DUP 5
SRR1766469.994884 chr7 158349819 N chr7 158349971 N DEL 5
SRR1766466.8164647 chr7 158349769 N chr7 158349971 N DEL 5
SRR1766472.8245438 chr7 158349777 N chr7 158349979 N DEL 5
SRR1766478.8359513 chr8 6680909 N chr8 6680979 N DUP 5
SRR1766480.6760403 chr8 6680830 N chr8 6680902 N DEL 5
SRR1766466.7115941 chr8 6680806 N chr8 6680908 N DEL 5
SRR1766467.7910307 chr8 6680939 N chr8 6681013 N DUP 5
SRR1766448.2868102 chr18 79969480 N chr18 79969533 N DEL 5
SRR1766464.9228770 chr7 27987447 N chr7 27987732 N DUP 7
SRR1766445.8408246 chr8 117973949 N chr8 117974037 N DUP 9
SRR1766446.1990774 chr13 87990186 N chr13 87990243 N DEL 32
SRR1766443.10189656 chr13 87990186 N chr13 87990243 N DEL 56
SRR1766469.7932559 chr13 87990186 N chr13 87990243 N DEL 57
SRR1766457.5232709 chr13 87990186 N chr13 87990243 N DEL 60
SRR1766463.7962679 chr13 87990186 N chr13 87990243 N DEL 53
SRR1766455.7092090 chr13 87990186 N chr13 87990243 N DEL 42
SRR1766445.812646 chr13 87990186 N chr13 87990243 N DEL 41
SRR1766462.1762920 chr13 87990186 N chr13 87990243 N DEL 36
SRR1766464.3248739 chr13 87990186 N chr13 87990243 N DEL 35
SRR1766468.495698 chr13 87990186 N chr13 87990243 N DEL 18
SRR1766479.9892609 chr13 87990186 N chr13 87990243 N DEL 15
SRR1766475.4352322 chr13 87990186 N chr13 87990243 N DEL 13
SRR1766449.3646662 chr13 87990186 N chr13 87990243 N DEL 13
SRR1766458.1705585 chr13 87990186 N chr13 87990243 N DEL 12
SRR1766474.4565614 chr13 87990189 N chr13 87990246 N DEL 9
SRR1766447.5873933 chr13 87990189 N chr13 87990246 N DEL 9
SRR1766453.2974310 chr13 87990190 N chr13 87990247 N DEL 9
SRR1766444.1227352 chr3 197876949 N chr3 197877022 N DEL 5
SRR1766478.1361215 chr3 197876949 N chr3 197877022 N DEL 5
SRR1766443.5551694 chr3 197876949 N chr3 197877022 N DEL 5
SRR1766476.6584642 chr3 197876949 N chr3 197877022 N DEL 5
SRR1766466.7710239 chr3 197876949 N chr3 197877022 N DEL 5
SRR1766448.9017750 chr3 197876963 N chr3 197877036 N DEL 1
SRR1766447.731041 chr3 197876976 N chr3 197877335 N DUP 5
SRR1766442.30816434 chr3 197877155 N chr3 197877336 N DEL 5
SRR1766479.8078858 chr3 197877155 N chr3 197877336 N DEL 5
SRR1766443.7016715 chr3 197877048 N chr3 197877335 N DUP 5
SRR1766484.10676322 chr3 197876956 N chr3 197877099 N DUP 5
SRR1766449.10094500 chr3 197877048 N chr3 197877335 N DUP 5
SRR1766474.10425239 chr3 197876975 N chr3 197877336 N DEL 5
SRR1766442.30816434 chr3 197877264 N chr3 197877335 N DUP 5
SRR1766443.5551694 chr3 197877048 N chr3 197877335 N DUP 5
SRR1766442.25179336 chr3 197877048 N chr3 197877335 N DUP 5
SRR1766463.875109 chr3 197877048 N chr3 197877335 N DUP 5
SRR1766467.1482159 chr3 197877048 N chr3 197877335 N DUP 5
SRR1766457.2280535 chr3 197877336 N chr3 197877659 N DUP 5
SRR1766462.1164322 chr3 197877060 N chr3 197877743 N DUP 5
SRR1766473.2847703 chr3 197876976 N chr3 197877335 N DUP 5
SRR1766463.4770637 chr3 197877171 N chr3 197877712 N DEL 4
SRR1766445.5802720 chr3 197877135 N chr3 197877712 N DEL 5
SRR1766442.29893613 chr3 197877135 N chr3 197877712 N DEL 5
SRR1766442.4193457 chr3 197877135 N chr3 197877712 N DEL 5
SRR1766471.1564158 chr3 197877135 N chr3 197877712 N DEL 5
SRR1766442.10766529 chr3 197877336 N chr3 197877661 N DEL 10
SRR1766480.2547678 chr3 197877099 N chr3 197877712 N DEL 5
SRR1766459.4277807 chr3 197877063 N chr3 197877712 N DEL 10
SRR1766442.35079802 chr3 197877099 N chr3 197877712 N DEL 5
SRR1766460.9958473 chr3 197877099 N chr3 197877712 N DEL 5
SRR1766462.5157039 chr3 197877099 N chr3 197877712 N DEL 5
SRR1766472.2421086 chr3 197877099 N chr3 197877712 N DEL 5
SRR1766485.9857312 chr3 197877099 N chr3 197877712 N DEL 5
SRR1766450.607177 chr3 197876991 N chr3 197877712 N DEL 5
SRR1766465.8320984 chr3 197876991 N chr3 197877712 N DEL 5
SRR1766473.3639750 chr3 197876991 N chr3 197877712 N DEL 5
SRR1766451.8991757 chr3 197876999 N chr3 197877720 N DEL 5
SRR1766475.1160353 chr22 46290645 N chr22 46290791 N DEL 5
SRR1766446.2219432 chr22 48992309 N chr22 48992407 N DEL 9
SRR1766474.7674137 chr22 48992310 N chr22 48992408 N DEL 9
SRR1766447.3577550 chr22 48992362 N chr22 48992448 N DEL 1
SRR1766450.4222228 chr2 240961895 N chr2 240962123 N DUP 5
SRR1766467.4482619 chr21 44404129 N chr21 44404466 N DUP 3
SRR1766442.26499947 chr21 44404130 N chr21 44404467 N DUP 2
SRR1766470.6113389 chr8 142116253 N chr8 142116746 N DEL 15
SRR1766449.9909730 chr8 142116241 N chr8 142116434 N DEL 8
SRR1766460.9100588 chr8 142116260 N chr8 142116737 N DEL 5
SRR1766484.1887313 chr8 142116246 N chr8 142116431 N DEL 5
SRR1766460.879122 chr8 142116186 N chr8 142116269 N DUP 10
SRR1766461.9765918 chr8 142116267 N chr8 142116736 N DEL 19
SRR1766451.76931 chr8 142116303 N chr8 142116736 N DEL 7
SRR1766474.5479588 chr8 142116194 N chr8 142116309 N DUP 13
SRR1766477.6161398 chr8 142115942 N chr8 142116333 N DUP 9
SRR1766442.45343044 chr8 142116268 N chr8 142116345 N DEL 10
SRR1766461.10807979 chr8 142116230 N chr8 142116437 N DUP 5
SRR1766459.5024419 chr8 142116422 N chr8 142116675 N DEL 6
SRR1766486.10295875 chr8 142116246 N chr8 142116435 N DEL 21
SRR1766442.23242165 chr8 142116109 N chr8 142116433 N DEL 13
SRR1766481.7044046 chr8 142116043 N chr8 142116443 N DEL 3
SRR1766477.671722 chr8 142116179 N chr8 142116484 N DEL 4
SRR1766457.2735558 chr8 142116473 N chr8 142116550 N DEL 9
SRR1766479.8061485 chr8 142116231 N chr8 142116556 N DEL 9
SRR1766459.136911 chr8 142115961 N chr8 142116570 N DEL 10
SRR1766460.879122 chr8 142116628 N chr8 142116783 N DUP 18
SRR1766447.10103305 chr8 142116245 N chr8 142116650 N DEL 5
SRR1766463.2268455 chr8 142116225 N chr8 142116764 N DUP 3
SRR1766449.5310206 chr8 142116225 N chr8 142116764 N DUP 5
SRR1766481.7044046 chr8 142116225 N chr8 142116764 N DUP 5
SRR1766460.5955407 chr8 142116250 N chr8 142116791 N DEL 5
SRR1766467.9812726 chr8 142116250 N chr8 142116791 N DEL 5
SRR1766474.7036554 chr8 142116250 N chr8 142116791 N DEL 5
SRR1766469.848220 chr8 142116250 N chr8 142116791 N DEL 5
SRR1766446.7967599 chr8 142116250 N chr8 142116791 N DEL 5
SRR1766449.1491774 chr8 142115958 N chr8 142116791 N DEL 5
SRR1766469.4816792 chr8 142115958 N chr8 142116791 N DEL 5
SRR1766443.7504265 chr8 142115958 N chr8 142116791 N DEL 5
SRR1766478.7448931 chr8 142115958 N chr8 142116791 N DEL 5
SRR1766442.33595812 chr8 142116045 N chr8 142116797 N DEL 5
SRR1766468.125922 chr2 141324176 N chr2 141324263 N DEL 5
SRR1766448.1102754 chr19 7640004 N chr19 7640135 N DUP 8
SRR1766484.10191319 chr19 7640169 N chr19 7640376 N DEL 3
SRR1766457.1348101 chr19 7640147 N chr19 7640632 N DEL 14
SRR1766467.10960619 chr19 7640132 N chr19 7640619 N DEL 7
SRR1766446.9366976 chr19 7640185 N chr19 7640260 N DEL 5
SRR1766461.9420238 chr19 7640206 N chr19 7640505 N DEL 11
SRR1766459.10825638 chr19 7640266 N chr19 7640671 N DEL 2
SRR1766450.8703190 chr19 7640270 N chr19 7640593 N DEL 1
SRR1766459.2345881 chr19 7640270 N chr19 7640593 N DEL 4
SRR1766466.4464312 chr19 7640273 N chr19 7640628 N DEL 5
SRR1766453.10121645 chr19 7640259 N chr19 7640486 N DEL 2
SRR1766468.6484053 chr19 7640218 N chr19 7640645 N DUP 5
SRR1766474.7384139 chr19 7640383 N chr19 7640454 N DEL 2
SRR1766472.10252237 chr19 7640284 N chr19 7640687 N DUP 5
SRR1766479.8359434 chr19 7640293 N chr19 7640462 N DUP 6
SRR1766484.10426568 chr19 7640336 N chr19 7640661 N DUP 4
SRR1766442.31602047 chr19 7640109 N chr19 7640334 N DEL 5
SRR1766482.7113450 chr19 7640356 N chr19 7640645 N DUP 12
SRR1766480.2630266 chr19 7640460 N chr19 7640575 N DEL 6
SRR1766471.11517789 chr19 7640290 N chr19 7640369 N DEL 10
SRR1766450.10496323 chr19 7640327 N chr19 7640496 N DUP 9
SRR1766442.32229991 chr19 7640327 N chr19 7640496 N DUP 9
SRR1766451.287711 chr19 7640395 N chr19 7640660 N DUP 8
SRR1766442.14653607 chr19 7640438 N chr19 7640687 N DUP 13
SRR1766465.1676595 chr19 7640414 N chr19 7640645 N DUP 9
SRR1766466.1290398 chr19 7640115 N chr19 7640468 N DEL 1
SRR1766471.6561278 chr19 7640018 N chr19 7640515 N DEL 5
SRR1766463.1473794 chr19 7640335 N chr19 7640538 N DEL 18
SRR1766456.3708421 chr19 7640581 N chr19 7640652 N DUP 3
SRR1766447.4780252 chr19 7640293 N chr19 7640542 N DEL 11
SRR1766474.1694267 chr19 7640462 N chr19 7640571 N DEL 8
SRR1766448.3873239 chr19 7640594 N chr19 7640645 N DUP 8
SRR1766483.7795068 chr19 7640600 N chr19 7640661 N DUP 10
SRR1766457.1348101 chr19 7640327 N chr19 7640618 N DEL 15
SRR1766483.6278071 chr19 7640195 N chr19 7640624 N DEL 7
SRR1766446.2767360 chr19 7640291 N chr19 7640628 N DEL 11
SRR1766444.2741862 chr19 7640097 N chr19 7640636 N DEL 5
SRR1766462.6250909 chr6 167575839 N chr6 167575987 N DEL 10
SRR1766465.3444603 chr6 167575839 N chr6 167575987 N DEL 8
SRR1766447.5567148 chr6 167575831 N chr6 167576000 N DEL 2
SRR1766453.10629345 chr14 87964237 N chr14 87964298 N DEL 2
SRR1766480.1510414 chr14 87964237 N chr14 87964298 N DEL 5
SRR1766473.4261016 chr14 87964237 N chr14 87964298 N DEL 5
SRR1766442.11565169 chr14 87964228 N chr14 87964287 N DUP 5
SRR1766461.10283133 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766442.18698955 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766470.1241109 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766468.6828619 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766450.7043120 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766472.881253 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766477.10423829 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766453.4048779 chr14 87964227 N chr14 87964286 N DUP 5
SRR1766461.5007509 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766473.8392587 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766485.11848538 chr14 87964218 N chr14 87964277 N DUP 5
SRR1766460.4729469 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766459.11235383 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766443.6547947 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766478.3943116 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766452.8489192 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766483.8791873 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766457.8147653 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766450.1629133 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766456.3280815 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766449.8845176 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766486.527201 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766462.7145271 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766467.11352228 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766471.1568680 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766442.593284 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766449.3223263 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766459.5854221 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766447.2234847 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766468.6562681 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766482.9492861 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766482.12922659 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766486.8781190 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766452.6372598 chr14 87964298 N chr14 87964357 N DUP 5
SRR1766444.5113360 chr14 87964237 N chr14 87964298 N DEL 5
SRR1766483.10519496 chr14 87964237 N chr14 87964298 N DEL 5
SRR1766467.1655427 chr14 87964237 N chr14 87964298 N DEL 5
SRR1766442.14802336 chr14 87964237 N chr14 87964298 N DEL 5
SRR1766468.2999378 chr14 87964238 N chr14 87964299 N DEL 5
SRR1766442.21672152 chr14 87964239 N chr14 87964300 N DEL 5
SRR1766453.4644222 chr8 1698394 N chr8 1698450 N DUP 7
SRR1766455.5286534 chr8 1698454 N chr8 1698512 N DEL 5
SRR1766447.3412355 chr8 1698544 N chr8 1698690 N DEL 5
SRR1766461.6206713 chr8 1698452 N chr8 1698508 N DUP 5
SRR1766451.2668165 chr8 1698562 N chr8 1699055 N DEL 8
SRR1766446.588066 chr8 1698487 N chr8 1698631 N DUP 10
SRR1766450.3425732 chr8 1698660 N chr8 1699096 N DEL 5
SRR1766442.12704653 chr8 1698660 N chr8 1699096 N DEL 5
SRR1766477.10707876 chr8 1698652 N chr8 1699088 N DEL 15
SRR1766472.10156255 chr8 1698388 N chr8 1698617 N DEL 7
SRR1766451.2157039 chr8 1698740 N chr8 1699088 N DEL 5
SRR1766467.5260057 chr8 1698670 N chr8 1698757 N DUP 5
SRR1766477.2277245 chr8 1698518 N chr8 1698664 N DEL 10
SRR1766465.6279546 chr8 1698407 N chr8 1698698 N DEL 20
SRR1766481.10438027 chr8 1698461 N chr8 1698807 N DUP 5
SRR1766442.36913523 chr8 1698664 N chr8 1698808 N DUP 5
SRR1766461.6908107 chr8 1698752 N chr8 1698808 N DUP 22
SRR1766484.93610 chr8 1698664 N chr8 1698808 N DUP 10
SRR1766478.6232040 chr8 1698752 N chr8 1698808 N DUP 10
SRR1766455.2025403 chr8 1698664 N chr8 1698808 N DUP 20
SRR1766448.4390109 chr8 1698394 N chr8 1698854 N DUP 5
SRR1766447.5521092 chr8 1698709 N chr8 1698765 N DUP 22
SRR1766453.1875414 chr8 1698450 N chr8 1698798 N DEL 30
SRR1766484.93610 chr8 1698410 N chr8 1698758 N DEL 5
SRR1766447.3412355 chr8 1698440 N chr8 1698788 N DEL 15
SRR1766481.4696832 chr8 1698418 N chr8 1698766 N DEL 6
SRR1766454.6774206 chr8 1698483 N chr8 1698774 N DEL 5
SRR1766483.4656267 chr8 1698483 N chr8 1698774 N DEL 5
SRR1766452.175877 chr8 1698439 N chr8 1698787 N DEL 2
SRR1766442.18425688 chr8 1698476 N chr8 1698910 N DUP 5
SRR1766474.3682491 chr8 1698411 N chr8 1698816 N DEL 4
SRR1766457.7471931 chr8 1698536 N chr8 1698827 N DEL 5
SRR1766462.6099946 chr8 1698587 N chr8 1698847 N DEL 5
SRR1766466.10462504 chr8 1698786 N chr8 1698982 N DUP 7
SRR1766477.10707876 chr8 1698407 N chr8 1698895 N DEL 6
SRR1766459.8806486 chr8 1698808 N chr8 1698923 N DEL 15
SRR1766442.42143536 chr8 1698830 N chr8 1698945 N DEL 5
SRR1766448.3198592 chr8 1698473 N chr8 1698935 N DEL 10
SRR1766447.6950828 chr8 1698870 N chr8 1698985 N DEL 5
SRR1766453.2407385 chr8 1698435 N chr8 1698985 N DEL 5
SRR1766467.10088998 chr8 1698508 N chr8 1699087 N DUP 5
SRR1766442.21944096 chr8 1698498 N chr8 1699103 N DUP 5
SRR1766457.1967128 chr8 1698561 N chr8 1699023 N DEL 15
SRR1766465.2082162 chr8 1698707 N chr8 1699055 N DEL 5
SRR1766451.2668165 chr8 1698536 N chr8 1699060 N DEL 1
SRR1766480.7862629 chr8 1698691 N chr8 1699070 N DEL 1
SRR1766458.5687517 chr8 1698447 N chr8 1699085 N DEL 5
SRR1766477.8006940 chr8 1699025 N chr8 1699088 N DEL 5
SRR1766482.10900186 chr8 1698879 N chr8 1699113 N DEL 5
SRR1766465.416450 chr8 1698879 N chr8 1699113 N DEL 5
SRR1766457.8364109 chr8 1698532 N chr8 1699113 N DEL 6
SRR1766443.2781559 chr8 1698532 N chr8 1699113 N DEL 5
SRR1766484.5068096 chr8 1698532 N chr8 1699113 N DEL 5
SRR1766479.1983418 chr8 1698532 N chr8 1699113 N DEL 5
SRR1766484.11241231 chr8 1698532 N chr8 1699113 N DEL 5
SRR1766442.29334801 chr18 78755796 N chr18 78755972 N DUP 12
SRR1766471.2193416 chr18 78755792 N chr18 78755968 N DUP 10
SRR1766449.2394043 chr18 78755818 N chr18 78755973 N DUP 5
SRR1766465.6559008 chr18 78755813 N chr18 78755968 N DUP 3
SRR1766480.4328314 chr18 78755872 N chr18 78756029 N DEL 25
SRR1766475.615956 chr9 137861489 N chr9 137861569 N DEL 5
SRR1766442.40012687 chr9 137861493 N chr9 137861710 N DEL 13
SRR1766478.3188328 chr9 137861503 N chr9 137861714 N DEL 7
SRR1766479.11899665 chr9 137861506 N chr9 137861571 N DEL 1
SRR1766474.6683467 chr9 137861492 N chr9 137861542 N DUP 2
SRR1766462.8470861 chr5 1543492 N chr5 1543670 N DUP 6
SRR1766460.3535056 chr5 1543593 N chr5 1543690 N DUP 2
SRR1766442.19638477 chr5 1543478 N chr5 1543685 N DEL 3
SRR1766442.742115 chrY 10773275 N chrY 10773371 N DEL 13
SRR1766468.5919514 chr8 79730462 N chr8 79730545 N DUP 6
SRR1766454.7344130 chr8 79730445 N chr8 79730574 N DUP 1
SRR1766464.2190590 chr8 79730478 N chr8 79730609 N DUP 10
SRR1766443.3156513 chr5 180312202 N chr5 180312347 N DEL 2
SRR1766457.7522940 chr5 180312182 N chr5 180312359 N DEL 7
SRR1766477.361206 chr5 49687 N chr5 49778 N DEL 1
SRR1766472.9134466 chr5 49687 N chr5 49778 N DEL 4
SRR1766477.3911342 chr5 49687 N chr5 49778 N DEL 11
SRR1766481.4145111 chr5 49687 N chr5 49778 N DEL 11
SRR1766466.1475842 chr14 102942963 N chr14 102943126 N DUP 4
SRR1766463.5437201 chr14 102942797 N chr14 102943122 N DEL 6
SRR1766482.6251085 chr14 102942906 N chr14 102943071 N DEL 3
SRR1766442.44095027 chr14 102942908 N chr14 102943073 N DEL 1
SRR1766443.7223220 chr4 117740001 N chr4 117740063 N DUP 20
SRR1766486.714908 chr4 117740001 N chr4 117740063 N DUP 20
SRR1766481.1396643 chr4 117740001 N chr4 117740063 N DUP 26
SRR1766453.5765675 chr4 117740001 N chr4 117740063 N DUP 27
SRR1766485.2393910 chr4 117740001 N chr4 117740063 N DUP 34
SRR1766471.2332312 chr4 117740001 N chr4 117740063 N DUP 36
SRR1766448.1984575 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766442.113303 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766462.4751505 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766470.7062168 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766467.6169663 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766455.7778042 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766442.23983098 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766464.5262491 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766442.11958196 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766445.9433921 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766469.2490008 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766465.11141919 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766477.4403156 chr4 117740001 N chr4 117740063 N DUP 37
SRR1766459.1191571 chr4 117740001 N chr4 117740063 N DUP 39
SRR1766442.46781775 chr4 117740001 N chr4 117740063 N DUP 41
SRR1766442.22613791 chr4 117740053 N chr4 117740136 N DEL 14
SRR1766455.4700077 chr4 117740055 N chr4 117740138 N DEL 12
SRR1766465.5813673 chr4 117740055 N chr4 117740138 N DEL 12
SRR1766477.1375051 chr4 117740054 N chr4 117740137 N DEL 13
SRR1766442.8627486 chr4 117740059 N chr4 117740142 N DEL 8
SRR1766475.11288262 chr4 117740060 N chr4 117740143 N DEL 7
SRR1766447.8751724 chr4 117740226 N chr4 117740320 N DEL 8
SRR1766474.8583943 chr4 117740226 N chr4 117740320 N DEL 9
SRR1766476.1504280 chr4 117740226 N chr4 117740320 N DEL 9
SRR1766471.2358954 chr4 117740226 N chr4 117740320 N DEL 10
SRR1766442.10497564 chr4 117740226 N chr4 117740320 N DEL 11
SRR1766458.3851732 chr4 117740226 N chr4 117740320 N DEL 24
SRR1766462.8081067 chr4 117740226 N chr4 117740320 N DEL 24
SRR1766484.9652404 chr4 117740226 N chr4 117740320 N DEL 26
SRR1766458.1000470 chr4 117740226 N chr4 117740320 N DEL 26
SRR1766467.607608 chr4 117740226 N chr4 117740320 N DEL 26
SRR1766468.7713097 chr4 117740226 N chr4 117740320 N DEL 29
SRR1766474.1401520 chr4 117740226 N chr4 117740320 N DEL 30
SRR1766462.5862362 chr4 117740226 N chr4 117740320 N DEL 30
SRR1766464.4587641 chr4 117740226 N chr4 117740320 N DEL 31
SRR1766464.6645833 chr4 117740226 N chr4 117740320 N DEL 32
SRR1766465.8520346 chr4 117740240 N chr4 117740334 N DEL 1
SRR1766453.2545477 chr4 117740228 N chr4 117740322 N DEL 13
SRR1766455.8877986 chr4 117740232 N chr4 117740326 N DEL 9
SRR1766465.762195 chr4 117740227 N chr4 117740321 N DEL 14
SRR1766450.5377606 chr4 117740233 N chr4 117740327 N DEL 8
SRR1766450.4606567 chr16 89342033 N chr16 89342206 N DUP 20
SRR1766447.10828257 chr16 89342064 N chr16 89342195 N DUP 2
SRR1766456.3302408 chr16 89342052 N chr16 89342183 N DUP 6
SRR1766465.6312542 chr16 89341991 N chr16 89342163 N DEL 4
SRR1766448.9274559 chr16 89342136 N chr16 89342227 N DEL 48
SRR1766467.11546382 chr16 89342136 N chr16 89342227 N DEL 38
SRR1766477.4580543 chr16 89342136 N chr16 89342227 N DEL 44
SRR1766448.733517 chr16 89342136 N chr16 89342227 N DEL 25
SRR1766448.8949338 chr16 89342136 N chr16 89342227 N DEL 23
SRR1766465.211241 chr16 89342136 N chr16 89342227 N DEL 19
SRR1766462.8886384 chr16 89342136 N chr16 89342227 N DEL 18
SRR1766466.5641529 chr16 89342011 N chr16 89342231 N DEL 8
SRR1766446.7650567 chrX 1297301 N chrX 1297473 N DEL 7
SRR1766472.5213963 chrX 1297285 N chrX 1297398 N DUP 3
SRR1766485.8654523 chrX 1297286 N chrX 1297399 N DUP 2
SRR1766485.8500084 chrX 1297359 N chrX 1297415 N DUP 5
SRR1766469.8009412 chrX 1297296 N chrX 1297580 N DUP 5
SRR1766444.3895079 chrX 1297381 N chrX 1297496 N DEL 5
SRR1766444.3318161 chrX 1297273 N chrX 1297386 N DUP 9
SRR1766442.13007365 chrX 1297296 N chrX 1297580 N DUP 5
SRR1766472.10773969 chrX 1297339 N chrX 1297452 N DUP 10
SRR1766467.7000389 chrX 1297273 N chrX 1297329 N DUP 5
SRR1766445.9602061 chrX 1297339 N chrX 1297395 N DUP 5
SRR1766444.5561551 chrX 1297273 N chrX 1297329 N DUP 5
SRR1766442.16069429 chrX 1297273 N chrX 1297329 N DUP 5
SRR1766474.10119131 chrX 1297309 N chrX 1297593 N DUP 2
SRR1766483.8250036 chrX 1297363 N chrX 1297533 N DUP 5
SRR1766442.10509576 chrX 1297339 N chrX 1297395 N DUP 5
SRR1766455.4138885 chrX 1297342 N chrX 1297398 N DUP 5
SRR1766478.4910135 chrX 1297339 N chrX 1297395 N DUP 5
SRR1766444.4129254 chrX 1297339 N chrX 1297395 N DUP 5
SRR1766484.6416978 chrX 1297285 N chrX 1297398 N DUP 1
SRR1766476.10407791 chrX 1297415 N chrX 1297473 N DEL 10
SRR1766455.901455 chrX 1297360 N chrX 1297416 N DUP 5
SRR1766445.5498862 chrX 1297273 N chrX 1297443 N DUP 10
SRR1766445.59329 chrX 1297410 N chrX 1297466 N DUP 5
SRR1766452.4171265 chrX 1297412 N chrX 1297468 N DUP 5
SRR1766443.1933880 chrX 1297340 N chrX 1297453 N DUP 10
SRR1766442.20723698 chrX 1297339 N chrX 1297452 N DUP 10
SRR1766486.7493480 chrX 1297409 N chrX 1297465 N DUP 5
SRR1766450.2340510 chrX 1297409 N chrX 1297465 N DUP 5
SRR1766470.10770788 chrX 1297409 N chrX 1297465 N DUP 10
SRR1766475.9927873 chrX 1297423 N chrX 1297479 N DUP 5
SRR1766470.2021591 chrX 1297294 N chrX 1297409 N DEL 9
SRR1766442.6447563 chrX 1297409 N chrX 1297465 N DUP 5
SRR1766445.4130578 chrX 1297273 N chrX 1297443 N DUP 5
SRR1766458.5227782 chrX 1297303 N chrX 1297418 N DEL 5
SRR1766463.6357 chrX 1297294 N chrX 1297409 N DEL 5
SRR1766486.3736299 chrX 1297294 N chrX 1297409 N DEL 5
SRR1766460.9536043 chrX 1297472 N chrX 1297528 N DUP 5
SRR1766477.7472782 chrX 1297472 N chrX 1297585 N DUP 5
SRR1766473.9731125 chrX 1297339 N chrX 1297509 N DUP 5
SRR1766445.8876915 chrX 1297263 N chrX 1297547 N DUP 12
SRR1766474.4541691 chrX 1297473 N chrX 1297529 N DUP 10
SRR1766464.3259875 chrX 1297472 N chrX 1297528 N DUP 5
SRR1766442.29116909 chrX 1297472 N chrX 1297528 N DUP 5
SRR1766454.8963487 chrX 1297486 N chrX 1297542 N DUP 10
SRR1766442.36238930 chrX 1297300 N chrX 1297472 N DEL 5
SRR1766463.3610676 chr3 60860390 N chr3 60860455 N DUP 11
SRR1766479.13600969 chr3 60860390 N chr3 60860455 N DUP 11
SRR1766472.3986952 chr3 60860390 N chr3 60860455 N DUP 11
SRR1766473.817752 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766454.2085433 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766444.1734587 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766448.7267246 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766460.10344168 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766477.10564264 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766465.5888777 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766483.7088928 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766448.9888280 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766444.1734587 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766473.9139992 chr3 60860423 N chr3 60860532 N DUP 10
SRR1766479.13726865 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766452.6164498 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766471.697922 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766462.5195647 chr13 35124677 N chr13 35124778 N DUP 6
SRR1766442.15532860 chr13 35124677 N chr13 35124778 N DUP 7
SRR1766464.9739716 chr13 35124677 N chr13 35124778 N DUP 9
SRR1766466.6274090 chr13 35124677 N chr13 35124778 N DUP 9
SRR1766462.4032350 chr13 35124778 N chr13 35124915 N DEL 12
SRR1766467.11041177 chr13 35124778 N chr13 35124915 N DEL 12
SRR1766483.2108351 chr13 35124698 N chr13 35124803 N DEL 7
SRR1766455.5139011 chr13 35124698 N chr13 35124803 N DEL 5
SRR1766460.3201285 chr13 35124805 N chr13 35124938 N DUP 5
SRR1766460.172793 chr13 35124811 N chr13 35124900 N DUP 5
SRR1766452.1913603 chr13 35124689 N chr13 35124814 N DEL 4
SRR1766459.1688739 chr13 35124691 N chr13 35124816 N DEL 2
SRR1766442.39915366 chr13 35124691 N chr13 35124816 N DEL 2
SRR1766476.1607148 chr6 62854108 N chr6 62854482 N DUP 5
SRR1766449.10079999 chr6 62854700 N chr6 62854852 N DUP 2
SRR1766448.9754101 chr6 62854724 N chr6 62854878 N DEL 5
SRR1766463.1989128 chr6 62854724 N chr6 62854878 N DEL 5
SRR1766452.8324457 chr6 62854420 N chr6 62854878 N DEL 5
SRR1766486.2200783 chr16 56566849 N chr16 56566926 N DUP 7
SRR1766456.1892722 chr12 39713610 N chr12 39713759 N DUP 10
SRR1766463.5244109 chr1 151601053 N chr1 151601300 N DUP 5
SRR1766455.2668786 chr1 151601046 N chr1 151601218 N DEL 3
SRR1766468.1198636 chr1 151601112 N chr1 151601283 N DEL 5
SRR1766442.14454341 chr6 155029272 N chr6 155029446 N DUP 5
SRR1766459.4340733 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766447.9969623 chr6 155029279 N chr6 155029428 N DUP 5
SRR1766481.3204764 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766442.19153552 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766460.1123536 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766457.3130520 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766463.9624436 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766484.2793484 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766451.3092731 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766458.3718914 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766450.3499149 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766449.4462807 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766469.7001720 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766456.5712257 chr6 155029354 N chr6 155029428 N DUP 5
SRR1766448.2470067 chr6 155029301 N chr6 155029352 N DEL 5
SRR1766456.827698 chr6 155029309 N chr6 155029360 N DEL 5
SRR1766447.11309676 chr6 155029341 N chr6 155029442 N DEL 5
SRR1766482.8600926 chr6 155029341 N chr6 155029442 N DEL 5
SRR1766481.10148901 chr6 155029316 N chr6 155029442 N DEL 5
SRR1766451.1991579 chr6 155029316 N chr6 155029442 N DEL 5
SRR1766448.10741316 chr6 155029291 N chr6 155029442 N DEL 5
SRR1766459.4322947 chr6 155029291 N chr6 155029442 N DEL 5
SRR1766479.2189361 chr6 155029291 N chr6 155029442 N DEL 5
SRR1766452.2424982 chr6 155029291 N chr6 155029442 N DEL 5
SRR1766447.934860 chr6 155029300 N chr6 155029451 N DEL 5
SRR1766442.34077466 chr12 130091658 N chr12 130091944 N DUP 5
SRR1766474.10691167 chr12 130091882 N chr12 130092092 N DUP 1
SRR1766484.8291433 chr12 130091796 N chr12 130091998 N DUP 5
SRR1766461.5533596 chr4 31749526 N chr4 31749576 N DUP 9
SRR1766461.9738282 chr11 64271206 N chr11 64271282 N DEL 6
SRR1766486.6511335 chr6 21797739 N chr6 21798089 N DEL 6
SRR1766462.4979903 chr6 21797856 N chr6 21797931 N DUP 5
SRR1766470.231487 chr6 21797969 N chr6 21798124 N DUP 5
SRR1766465.2601458 chr8 123315143 N chr8 123315495 N DEL 19
SRR1766442.21173843 chr8 123315143 N chr8 123315495 N DEL 20
SRR1766463.10957138 chr8 123315143 N chr8 123315495 N DEL 15
SRR1766456.4660246 chr8 123315143 N chr8 123315495 N DEL 20
SRR1766446.4033195 chr8 123315143 N chr8 123315495 N DEL 20
SRR1766473.3739623 chr8 123315265 N chr8 123315393 N DEL 1
SRR1766461.9696750 chr8 123315298 N chr8 123315957 N DEL 10
SRR1766461.9696750 chr8 123315305 N chr8 123315757 N DUP 10
SRR1766442.27991436 chr8 123315128 N chr8 123315276 N DEL 5
SRR1766466.5565595 chr8 123315314 N chr8 123315973 N DEL 7
SRR1766453.9408663 chr8 123315184 N chr8 123315585 N DEL 24
SRR1766485.4406859 chr8 123315190 N chr8 123315591 N DEL 13
SRR1766478.9536311 chr8 123315696 N chr8 123315750 N DEL 7
SRR1766466.4885941 chr8 123315673 N chr8 123316106 N DUP 10
SRR1766467.418309 chr8 123315396 N chr8 123315670 N DEL 5
SRR1766455.647993 chr8 123315223 N chr8 123315673 N DEL 8
SRR1766447.9461078 chr8 123315128 N chr8 123315676 N DEL 2
SRR1766472.3312019 chr8 123315128 N chr8 123315676 N DEL 2
SRR1766459.5475016 chr8 123315739 N chr8 123315867 N DEL 5
SRR1766447.11439771 chr8 123315696 N chr8 123315750 N DEL 7
SRR1766453.234582 chr8 123315696 N chr8 123315750 N DEL 9
SRR1766453.600780 chr8 123315248 N chr8 123315956 N DEL 5
SRR1766480.1413409 chr8 123315203 N chr8 123315960 N DEL 10
SRR1766485.1522065 chr8 123315209 N chr8 123315761 N DEL 4
SRR1766483.6352542 chr8 123315396 N chr8 123315850 N DEL 5
SRR1766479.13595924 chr8 123315872 N chr8 123316076 N DUP 5
SRR1766470.5008901 chr8 123315779 N chr8 123315983 N DUP 1
SRR1766459.3367184 chr8 123315357 N chr8 123315938 N DEL 5
SRR1766461.9996824 chr8 123315315 N chr8 123315392 N DUP 9
SRR1766465.4373280 chr8 123315276 N chr8 123316061 N DUP 7
SRR1766482.2037079 chr8 123315315 N chr8 123315392 N DUP 7
SRR1766451.94572 chr8 123315280 N chr8 123316065 N DUP 7
SRR1766443.2470571 chr8 123315730 N chr8 123316060 N DUP 11
SRR1766458.4382914 chr8 123315403 N chr8 123316061 N DEL 7
SRR1766442.26256524 chr8 123315403 N chr8 123316061 N DEL 7
SRR1766470.5608889 chr8 123315403 N chr8 123316061 N DEL 7
SRR1766458.3264261 chr8 123315403 N chr8 123316061 N DEL 7
SRR1766474.10031121 chr8 123315403 N chr8 123316061 N DEL 7
SRR1766460.1902377 chr8 123316063 N chr8 123316112 N DUP 8
SRR1766469.968090 chr8 123315227 N chr8 123316061 N DEL 7
SRR1766485.9532452 chr7 157439615 N chr7 157439770 N DEL 1
SRR1766485.10803759 chr7 157439460 N chr7 157439648 N DUP 4
SRR1766453.6678034 chr7 157439560 N chr7 157439664 N DUP 5
SRR1766449.10069429 chr7 157439560 N chr7 157439664 N DUP 5
SRR1766456.4058385 chr7 157439563 N chr7 157439931 N DUP 5
SRR1766450.606632 chr7 157439567 N chr7 157439935 N DUP 5
SRR1766459.8987944 chr7 157439570 N chr7 157439938 N DUP 5
SRR1766468.2429682 chr7 157439736 N chr7 157440000 N DEL 4
SRR1766484.9264159 chr7 157439776 N chr7 157439832 N DEL 6
SRR1766442.23239024 chr7 157439769 N chr7 157439825 N DEL 12
SRR1766448.2188717 chr7 157439773 N chr7 157439829 N DEL 5
SRR1766477.7695057 chr7 157439664 N chr7 157439825 N DEL 5
SRR1766442.43384812 chr7 157439776 N chr7 157439832 N DEL 5
SRR1766461.2169182 chr7 157439439 N chr7 157440017 N DUP 6
SRR1766471.9493631 chr7 157439725 N chr7 157439987 N DUP 5
SRR1766466.7060871 chr7 157439665 N chr7 157439930 N DEL 5
SRR1766455.5141976 chr7 157439483 N chr7 157439937 N DEL 5
SRR1766451.8174199 chr7 157439578 N chr7 157440104 N DUP 9
SRR1766463.10058916 chr7 157439691 N chr7 157440119 N DUP 5
SRR1766471.2054337 chr7 157439596 N chr7 157440124 N DEL 10
SRR1766472.5289661 chr7 157439598 N chr7 157440126 N DEL 9
SRR1766482.9649051 chr7 157439466 N chr7 157440134 N DEL 5
SRR1766455.4477233 chrX 40616946 N chrX 40616995 N DUP 6
SRR1766458.1257881 chrX 40616950 N chrX 40617023 N DUP 32
SRR1766454.618763 chrY 10976009 N chrY 10976111 N DEL 10
SRR1766455.6011185 chrY 10976009 N chrY 10976111 N DEL 10
SRR1766471.3670895 chrY 10976007 N chrY 10976119 N DEL 7
SRR1766473.7568319 chrY 10976103 N chrY 10976299 N DUP 5
SRR1766469.10857532 chrX 818511 N chrX 818836 N DUP 5
SRR1766475.768835 chrX 818492 N chrX 818546 N DEL 22
SRR1766476.5977634 chrX 818457 N chrX 818546 N DEL 20
SRR1766484.3957404 chrX 818457 N chrX 818546 N DEL 23
SRR1766449.10556070 chrX 818457 N chrX 818546 N DEL 15
SRR1766472.7772488 chrX 818428 N chrX 818546 N DEL 15
SRR1766485.2356778 chrX 818444 N chrX 818579 N DEL 2
SRR1766444.2927061 chrX 818434 N chrX 818552 N DEL 9
SRR1766478.1192260 chrX 818436 N chrX 818554 N DEL 7
SRR1766446.2502928 chrX 818573 N chrX 819011 N DUP 8
SRR1766446.1074889 chrX 818457 N chrX 818546 N DEL 17
SRR1766455.2207311 chrX 818457 N chrX 818546 N DEL 20
SRR1766449.4400899 chrX 818457 N chrX 818546 N DEL 22
SRR1766484.12259432 chrX 818457 N chrX 818546 N DEL 24
SRR1766475.4774066 chrX 818577 N chrX 818737 N DUP 5
SRR1766468.5874703 chrX 818377 N chrX 818632 N DEL 3
SRR1766459.2909969 chrX 818819 N chrX 818895 N DUP 8
SRR1766469.304078 chr14 21657486 N chr14 21657593 N DEL 1
SRR1766446.5661685 chr14 21657486 N chr14 21657593 N DEL 4
SRR1766479.12420950 chr11 1873732 N chr11 1873803 N DUP 5
SRR1766442.39483175 chr22 46609037 N chr22 46609156 N DEL 5
SRR1766475.976711 chr22 46609045 N chr22 46609164 N DEL 10
SRR1766471.5010619 chr22 46609067 N chr22 46609123 N DUP 7
SRR1766478.143743 chr22 46609061 N chr22 46609178 N DUP 3
SRR1766477.5624255 chr8 139997444 N chr8 139997696 N DEL 5
SRR1766482.6805526 chr8 139997532 N chr8 139998121 N DEL 6
SRR1766442.15231913 chr8 139997335 N chr8 139997451 N DEL 5
SRR1766478.10582109 chr8 139997585 N chr8 139998015 N DEL 5
SRR1766450.1492479 chr8 139997718 N chr8 139997787 N DEL 1
SRR1766459.2499329 chr8 139997718 N chr8 139997787 N DEL 4
SRR1766455.4851743 chr8 139997414 N chr8 139997732 N DUP 10
SRR1766469.5150890 chr8 139997342 N chr8 139997640 N DEL 10
SRR1766480.7119414 chr8 139997662 N chr8 139998044 N DUP 8
SRR1766473.3550911 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766450.6602475 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766469.11170539 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766472.4366138 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766478.6555588 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766472.4366138 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766485.2210979 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766462.9239351 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766466.3733020 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766470.10369951 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766442.670641 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766447.5321447 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766484.3639334 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766444.4991464 chr8 139997723 N chr8 139997814 N DEL 5
SRR1766465.3236566 chr8 139997799 N chr8 139998093 N DEL 5
SRR1766478.10436843 chr8 139997735 N chr8 139997802 N DUP 6
SRR1766455.4815858 chr8 139997837 N chr8 139997928 N DEL 3
SRR1766450.3435331 chr8 139997827 N chr8 139997940 N DEL 5
SRR1766454.7224073 chr8 139997836 N chr8 139997927 N DEL 5
SRR1766475.7447168 chr8 139997836 N chr8 139997927 N DEL 5
SRR1766459.10936949 chr8 139997433 N chr8 139997865 N DEL 5
SRR1766447.10926585 chr8 139997836 N chr8 139997927 N DEL 5
SRR1766466.7196880 chr8 139997846 N chr8 139997937 N DEL 5
SRR1766479.13483865 chr8 139997836 N chr8 139997927 N DEL 5
SRR1766452.6211400 chr8 139997846 N chr8 139997937 N DEL 5
SRR1766467.3039504 chr8 139997836 N chr8 139997927 N DEL 5
SRR1766467.1265267 chr8 139997846 N chr8 139997937 N DEL 5
SRR1766470.3425506 chr8 139997690 N chr8 139997939 N DEL 3
SRR1766449.2248925 chr8 139997343 N chr8 139998047 N DEL 5
SRR1766475.8817472 chr8 139997690 N chr8 139998051 N DEL 5
SRR1766442.10485619 chr8 139997432 N chr8 139998067 N DEL 5
SRR1766473.952350 chr8 139997443 N chr8 139998210 N DUP 5
SRR1766477.11004873 chr8 139997440 N chr8 139998166 N DEL 5
SRR1766486.2197339 chr1 8952119 N chr1 8952435 N DUP 5
SRR1766466.4301354 chr1 173913876 N chr1 173914097 N DUP 5
SRR1766470.1980768 chr19 57137967 N chr19 57138264 N DEL 5
SRR1766453.8521863 chr19 57138063 N chr19 57138228 N DEL 6
SRR1766449.4570193 chr19 57137989 N chr19 57138060 N DUP 8
SRR1766469.10089654 chr19 57137989 N chr19 57138068 N DUP 5
SRR1766442.15979870 chr19 57138034 N chr19 57138141 N DUP 2
SRR1766445.3513444 chr19 57138016 N chr19 57138178 N DUP 14
SRR1766465.6743129 chr19 57138060 N chr19 57138116 N DUP 13
SRR1766475.7586315 chr19 57137986 N chr19 57138146 N DUP 12
SRR1766469.5791321 chr19 57137992 N chr19 57138139 N DUP 5
SRR1766469.10762129 chr19 57138052 N chr19 57138155 N DUP 10
SRR1766474.60635 chr19 57138024 N chr19 57138099 N DUP 13
SRR1766463.3412795 chr19 57138057 N chr19 57138133 N DUP 12
SRR1766481.5417566 chr19 57138007 N chr19 57138134 N DUP 4
SRR1766448.10590751 chr19 57137994 N chr19 57138067 N DEL 2
SRR1766457.8388299 chr19 57137986 N chr19 57138130 N DUP 7
SRR1766442.35089032 chr19 57138028 N chr19 57138152 N DUP 12
SRR1766463.4717118 chr19 57138033 N chr19 57138098 N DEL 4
SRR1766453.8693804 chr19 57138038 N chr19 57138139 N DEL 6
SRR1766442.38839232 chr19 57138011 N chr19 57138242 N DUP 14
SRR1766470.9249561 chr19 57138052 N chr19 57138231 N DUP 15
SRR1766451.1614682 chr7 68509466 N chr7 68509569 N DUP 1
SRR1766452.8471900 chrY 11032148 N chrY 11032419 N DUP 5
SRR1766473.8086953 chr13 20392562 N chr13 20392613 N DEL 6
SRR1766464.9957028 chr13 20392643 N chr13 20392886 N DEL 5
SRR1766459.3720 chr13 20392522 N chr13 20392660 N DUP 4
SRR1766480.4911187 chr13 20392525 N chr13 20392751 N DUP 5
SRR1766453.2115359 chr13 20392636 N chr13 20392750 N DUP 1
SRR1766482.11233668 chr13 20392716 N chr13 20392897 N DUP 1
SRR1766470.2270859 chr13 20392644 N chr13 20392863 N DUP 5
SRR1766484.9364275 chr22 42087669 N chr22 42088275 N DEL 1
SRR1766468.5777039 chr22 42087670 N chr22 42087976 N DEL 26
SRR1766473.8208453 chr22 42087669 N chr22 42088275 N DEL 20
SRR1766486.2777480 chr22 42087768 N chr22 42088374 N DEL 5
SRR1766472.2081827 chr22 42087844 N chr22 42088450 N DEL 10
SRR1766471.6319322 chr22 42087820 N chr22 42088424 N DUP 15
SRR1766447.5439204 chr22 42087916 N chr22 42088836 N DEL 3
SRR1766475.4032484 chr22 42087671 N chr22 42087975 N DUP 2
SRR1766458.5155559 chr22 42088023 N chr22 42088324 N DEL 36
SRR1766443.2575371 chr22 42087670 N chr22 42087976 N DEL 13
SRR1766472.8615351 chr22 42088257 N chr22 42088871 N DEL 5
SRR1766447.1295310 chr22 42088261 N chr22 42088871 N DEL 4
SRR1766453.5082174 chr22 42087726 N chr22 42088332 N DEL 10
SRR1766475.405940 chr5 95360576 N chr5 95360665 N DUP 14
SRR1766452.2519904 chr1 80700055 N chr1 80700156 N DEL 6
SRR1766442.21271732 chr1 80700055 N chr1 80700156 N DEL 6
SRR1766453.9961730 chr1 80700055 N chr1 80700156 N DEL 6
SRR1766468.5358476 chr1 80700056 N chr1 80700157 N DEL 6
SRR1766479.10728980 chr1 80700056 N chr1 80700157 N DEL 6
SRR1766471.5277653 chr15 97058369 N chr15 97058474 N DEL 1
SRR1766479.12623699 chr9 20417278 N chr9 20417443 N DEL 10
SRR1766466.11283389 chr9 20417146 N chr9 20417459 N DEL 20
SRR1766479.4174472 chrX 2166513 N chrX 2166576 N DEL 19
SRR1766459.10891684 chr14 32199763 N chr14 32199950 N DUP 3
SRR1766479.3797457 chr14 32199856 N chr14 32199953 N DUP 4
SRR1766466.834244 chr14 32199842 N chr14 32199958 N DEL 2
SRR1766451.8161233 chr9 119249974 N chr9 119250235 N DUP 5
SRR1766473.6198366 chr9 119250198 N chr9 119250259 N DEL 12
SRR1766442.39941293 chr9 119250088 N chr9 119250175 N DUP 1
SRR1766467.10720879 chr9 119250117 N chr9 119250188 N DUP 7
SRR1766474.11425769 chr5 15935450 N chr5 15935735 N DEL 4
SRR1766477.10629360 chr5 15935450 N chr5 15935735 N DEL 8
SRR1766456.708743 chr5 15935502 N chr5 15935787 N DEL 11
SRR1766466.7598979 chr14 34350232 N chr14 34350323 N DEL 10
SRR1766478.3735069 chr14 34349684 N chr14 34349840 N DEL 5
SRR1766469.9186669 chr14 34349958 N chr14 34350472 N DEL 10
SRR1766464.905893 chr14 34349446 N chr14 34350323 N DEL 5
SRR1766467.6724816 chr14 34349508 N chr14 34350071 N DUP 9
SRR1766475.7682053 chr14 34349666 N chr14 34349820 N DUP 5
SRR1766461.6769123 chr14 34349666 N chr14 34349820 N DUP 5
SRR1766482.13066334 chr14 34349682 N chr14 34349838 N DEL 5
SRR1766471.4002404 chr14 34349685 N chr14 34349841 N DEL 5
SRR1766442.27310654 chr14 34349680 N chr14 34349836 N DEL 5
SRR1766482.807045 chr14 34349687 N chr14 34349843 N DEL 4
SRR1766461.6617292 chr14 34349666 N chr14 34349820 N DUP 5
SRR1766442.10551951 chr14 34349666 N chr14 34349820 N DUP 5
SRR1766474.1345334 chr14 34350188 N chr14 34350247 N DUP 10
SRR1766484.11739419 chr14 34350188 N chr14 34350247 N DUP 10
SRR1766443.7042458 chr14 34350202 N chr14 34350323 N DEL 1
SRR1766461.6617292 chr14 34350232 N chr14 34350293 N DEL 10
SRR1766471.11192317 chr4 2430211 N chr4 2430401 N DEL 5
SRR1766459.8217098 chr4 2430211 N chr4 2430401 N DEL 5
SRR1766471.3624699 chr4 2430258 N chr4 2430322 N DEL 3
SRR1766463.1835312 chr4 2430239 N chr4 2430303 N DEL 5
SRR1766467.8803067 chr4 2430239 N chr4 2430303 N DEL 5
SRR1766466.6752984 chr4 2430240 N chr4 2430302 N DUP 10
SRR1766457.1214383 chr4 2430240 N chr4 2430302 N DUP 10
SRR1766459.4076190 chr4 2430242 N chr4 2430304 N DUP 9
SRR1766461.3257283 chr4 2430251 N chr4 2430313 N DUP 4
SRR1766442.41072175 chr4 2430274 N chr4 2430464 N DEL 5
SRR1766442.9222722 chr4 2430274 N chr4 2430464 N DEL 5
SRR1766442.43504385 chr4 2430274 N chr4 2430590 N DEL 5
SRR1766484.3306783 chr4 2430240 N chr4 2430302 N DUP 1
SRR1766470.182592 chr4 2430211 N chr4 2430590 N DEL 5
SRR1766476.6408816 chr4 2430211 N chr4 2430590 N DEL 5
SRR1766447.9505125 chr4 2430211 N chr4 2430590 N DEL 5
SRR1766472.2765096 chr4 2430211 N chr4 2430590 N DEL 5
SRR1766445.1595153 chr4 2430240 N chr4 2430302 N DUP 5
SRR1766486.5403168 chr4 2430220 N chr4 2430599 N DEL 6
SRR1766486.9435272 chr4 2430230 N chr4 2430294 N DEL 5
SRR1766442.20545169 chr4 2430302 N chr4 2430429 N DEL 5
SRR1766468.4224943 chr4 2430232 N chr4 2430296 N DEL 5
SRR1766467.884437 chr4 2430302 N chr4 2430429 N DEL 5
SRR1766480.5259121 chr4 2430240 N chr4 2430302 N DUP 5
SRR1766464.4500254 chr4 2430302 N chr4 2430429 N DEL 5
SRR1766475.11468194 chr4 2430337 N chr4 2430464 N DEL 3
SRR1766442.38568939 chr4 2430337 N chr4 2430464 N DEL 5
SRR1766462.3980863 chr4 2430240 N chr4 2430302 N DUP 10
SRR1766464.2511304 chr4 2430212 N chr4 2430400 N DUP 5
SRR1766480.2293355 chr4 2430230 N chr4 2430357 N DEL 5
SRR1766448.10564696 chr4 2430211 N chr4 2430401 N DEL 5
SRR1766449.21631 chr4 2430230 N chr4 2430609 N DEL 10
SRR1766459.1021521 chr4 2430274 N chr4 2430464 N DEL 5
SRR1766486.6383824 chr4 2430239 N chr4 2430303 N DEL 5
SRR1766444.679140 chr4 2430274 N chr4 2430464 N DEL 5
SRR1766442.44733692 chr4 2430275 N chr4 2430463 N DUP 5
SRR1766470.10527019 chr4 2430275 N chr4 2430463 N DUP 5
SRR1766442.12189952 chr4 2430274 N chr4 2430464 N DEL 5
SRR1766442.14571662 chr4 2430274 N chr4 2430464 N DEL 5
SRR1766472.2315687 chr4 2430316 N chr4 2430443 N DEL 1
SRR1766475.4602288 chr4 2430316 N chr4 2430443 N DEL 1
SRR1766442.20750782 chr4 2430274 N chr4 2430464 N DEL 5
SRR1766454.4358932 chr4 2430268 N chr4 2430584 N DEL 1
SRR1766448.5165837 chr4 2430268 N chr4 2430584 N DEL 2
SRR1766442.46558909 chr4 2430294 N chr4 2430419 N DUP 5
SRR1766482.4172599 chr4 2430429 N chr4 2430491 N DUP 5
SRR1766484.3807853 chr4 2430233 N chr4 2430486 N DEL 5
SRR1766462.10163703 chr4 2430337 N chr4 2430527 N DEL 5
SRR1766480.7590847 chr4 2430337 N chr4 2430527 N DEL 5
SRR1766442.31183505 chr4 2430337 N chr4 2430527 N DEL 5
SRR1766476.6230796 chr4 2430337 N chr4 2430527 N DEL 5
SRR1766449.6035769 chr4 2430337 N chr4 2430527 N DEL 5
SRR1766447.8204148 chr4 2430274 N chr4 2430527 N DEL 5
SRR1766481.2332007 chr4 2430274 N chr4 2430527 N DEL 5
SRR1766481.2332007 chr4 2430216 N chr4 2430532 N DEL 5
SRR1766483.5504906 chr4 2430302 N chr4 2430429 N DEL 5
SRR1766473.782496 chr4 2430337 N chr4 2430464 N DEL 10
SRR1766446.1767298 chr4 2430310 N chr4 2430437 N DEL 5
SRR1766483.10806468 chr4 2430230 N chr4 2430609 N DEL 5
SRR1766455.9398218 chr4 2430404 N chr4 2430594 N DEL 3
SRR1766471.11192317 chr4 2430337 N chr4 2430653 N DEL 5
SRR1766457.8278912 chr4 2430230 N chr4 2430672 N DEL 10
SRR1766444.679140 chr4 2430410 N chr4 2430726 N DEL 10
SRR1766464.2511304 chr4 2430410 N chr4 2430726 N DEL 5
SRR1766480.6588329 chr4 2430410 N chr4 2430726 N DEL 5
SRR1766442.35745760 chr4 2430227 N chr4 2430732 N DEL 5
SRR1766480.1687803 chr5 160504972 N chr5 160505148 N DEL 11
SRR1766447.4715364 chr5 160504952 N chr5 160505163 N DUP 6
SRR1766463.6215726 chr5 160504982 N chr5 160505154 N DUP 6
SRR1766464.1605111 chr5 160504862 N chr5 160505105 N DUP 5
SRR1766479.3893736 chr5 160505108 N chr5 160505221 N DEL 5
SRR1766446.10602129 chr5 160505108 N chr5 160505221 N DEL 6
SRR1766465.2906374 chr5 160505039 N chr5 160505161 N DUP 7
SRR1766460.6535811 chr5 160505112 N chr5 160505183 N DUP 5
SRR1766475.7188699 chr5 160505121 N chr5 160505232 N DUP 4
SRR1766456.6443496 chr5 160504879 N chr5 160505124 N DEL 1
SRR1766481.4632384 chr5 160505156 N chr5 160505232 N DUP 5
SRR1766459.3814504 chr5 160504928 N chr5 160505251 N DEL 5
SRR1766475.6382382 chr5 2219178 N chr5 2219793 N DEL 7
SRR1766467.5910894 chr5 2219205 N chr5 2219890 N DEL 2
SRR1766479.10029685 chr5 2219396 N chr5 2219780 N DEL 4
SRR1766485.1301976 chr5 2219387 N chr5 2219816 N DUP 3
SRR1766464.2434616 chr5 2219541 N chr5 2219795 N DEL 6
SRR1766472.11821186 chr5 2219487 N chr5 2219537 N DUP 10
SRR1766452.8939342 chr5 2219412 N chr5 2219600 N DUP 7
SRR1766480.8641988 chr22 46194965 N chr22 46195295 N DEL 20
SRR1766479.3452364 chr22 46194703 N chr22 46195026 N DUP 7
SRR1766442.46038382 chr22 46194970 N chr22 46195300 N DEL 20
SRR1766476.732756 chr22 46194970 N chr22 46195300 N DEL 15
SRR1766457.4210451 chr12 39712193 N chr12 39712530 N DUP 1
SRR1766482.13134835 chr12 39712193 N chr12 39712530 N DUP 1
SRR1766443.10275616 chr12 39712193 N chr12 39712530 N DUP 1
SRR1766485.2451622 chr12 39712174 N chr12 39712311 N DEL 7
SRR1766475.4798919 chr12 39712355 N chr12 39712458 N DUP 2
SRR1766478.10327167 chr12 39712315 N chr12 39712512 N DUP 13
SRR1766442.41243329 chr12 39712252 N chr12 39712513 N DUP 14
SRR1766460.3625296 chr12 39712561 N chr12 39712620 N DEL 8
SRR1766475.10588741 chr12 39712188 N chr12 39712485 N DEL 2
SRR1766473.1740543 chr12 39712188 N chr12 39712485 N DEL 1
SRR1766467.5678987 chr12 39712477 N chr12 39712544 N DEL 7
SRR1766463.8808939 chr12 39712265 N chr12 39712544 N DEL 3
SRR1766471.8788883 chr12 39712527 N chr12 39712642 N DEL 46
SRR1766477.11092086 chr10 7526686 N chr10 7526923 N DEL 1
SRR1766444.3363549 chr10 7526771 N chr10 7526828 N DUP 11
SRR1766455.6347094 chr10 7526771 N chr10 7526828 N DUP 12
SRR1766467.10990244 chr10 7526850 N chr10 7526983 N DUP 16
SRR1766462.1802173 chr10 7526781 N chr10 7526923 N DUP 12
SRR1766486.2647662 chr10 7526782 N chr10 7526924 N DUP 11
SRR1766481.4088628 chr10 7526840 N chr10 7526973 N DUP 21
SRR1766478.7249718 chr10 7526840 N chr10 7526973 N DUP 20
SRR1766453.7469241 chr10 7526840 N chr10 7526973 N DUP 20
SRR1766479.10906004 chr10 7526850 N chr10 7526983 N DUP 14
SRR1766460.4603530 chr10 7526740 N chr10 7526962 N DEL 6
SRR1766442.42882839 chr10 7526647 N chr10 7526979 N DEL 5
SRR1766462.1261323 chr10 7526668 N chr10 7527004 N DEL 1
SRR1766458.1714965 chr4 187024897 N chr4 187025040 N DEL 5
SRR1766450.7304544 chr4 187024973 N chr4 187025117 N DUP 3
SRR1766478.8089751 chr4 187024965 N chr4 187025109 N DEL 6
SRR1766471.7152244 chr9 137034440 N chr9 137034500 N DEL 1
SRR1766444.6567973 chr1 169737562 N chr1 169737618 N DEL 6
SRR1766472.1992594 chr13 113588899 N chr13 113588951 N DUP 5
SRR1766482.494686 chr13 113588899 N chr13 113588951 N DUP 5
SRR1766475.10398764 chr13 113588899 N chr13 113588951 N DUP 5
SRR1766476.6559939 chr18 47541662 N chr18 47541796 N DEL 4
SRR1766450.8441946 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766447.6330704 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766463.7736540 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766442.42485774 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766458.4848613 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766465.4970216 chr18 47541666 N chr18 47541800 N DEL 5
SRR1766479.11644161 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766442.39962950 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766485.959769 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766479.5585035 chr18 47541662 N chr18 47541796 N DEL 5
SRR1766460.5581142 chr18 47541662 N chr18 47541796 N DEL 7
SRR1766456.1079309 chr18 47541667 N chr18 47541801 N DEL 5
SRR1766459.3421580 chr12 117409564 N chr12 117409733 N DUP 1
SRR1766469.3895796 chr16 34583301 N chr16 34583420 N DEL 5
SRR1766476.2346164 chr16 34583311 N chr16 34583430 N DEL 3
SRR1766468.5144228 chr16 34583291 N chr16 34583362 N DUP 11
SRR1766457.8491967 chr16 34583311 N chr16 34583430 N DEL 5
SRR1766481.258881 chr16 34583311 N chr16 34583430 N DEL 5
SRR1766469.5829954 chr16 34583299 N chr16 34583393 N DUP 10
SRR1766447.399638 chr16 34583247 N chr16 34583318 N DUP 4
SRR1766464.835346 chr16 34583360 N chr16 34583456 N DEL 7
SRR1766481.11362387 chr16 34583334 N chr16 34583430 N DEL 4
SRR1766466.2453444 chr11 129580634 N chr11 129580754 N DEL 5
SRR1766445.1579622 chr11 129580634 N chr11 129580754 N DEL 5
SRR1766482.1732122 chr11 129580604 N chr11 129580675 N DUP 7
SRR1766486.9300017 chr11 129580620 N chr11 129580693 N DEL 5
SRR1766460.9970825 chr16 34754099 N chr16 34754219 N DUP 1
SRR1766449.6263814 chr9 80122947 N chr9 80123104 N DEL 6
SRR1766451.4286354 chr9 80122819 N chr9 80123403 N DUP 13
SRR1766481.9801896 chr9 80122819 N chr9 80123403 N DUP 13
SRR1766463.4934093 chr12 132528849 N chr12 132528922 N DEL 5
SRR1766462.5146556 chr22 15583248 N chr22 15583406 N DEL 1
SRR1766453.7158381 chr12 56075892 N chr12 56075991 N DEL 4
SRR1766482.6329777 chr12 56076049 N chr12 56076323 N DEL 5
SRR1766443.963052 chr12 56076306 N chr12 56076463 N DEL 3
SRR1766448.9800347 chr20 4089793 N chr20 4089850 N DEL 4
SRR1766446.2671068 chr14 79471020 N chr14 79471073 N DEL 5
SRR1766465.2562958 chr14 79471048 N chr14 79471103 N DEL 7
SRR1766477.8275190 chr14 79471048 N chr14 79471111 N DEL 15
SRR1766473.9396436 chr14 79471048 N chr14 79471111 N DEL 15
SRR1766442.27450871 chr14 79471059 N chr14 79471112 N DEL 4
SRR1766442.43452959 chr5 27427103 N chr5 27427167 N DUP 5
SRR1766442.22524350 chr5 27427103 N chr5 27427167 N DUP 5
SRR1766473.8165683 chr5 27427118 N chr5 27427206 N DUP 2
SRR1766472.11497897 chr5 27427118 N chr5 27427254 N DUP 3
SRR1766447.8171471 chr5 27427118 N chr5 27427254 N DUP 5
SRR1766476.7796081 chr5 27427137 N chr5 27427203 N DEL 5
SRR1766466.4019976 chr5 27427137 N chr5 27427203 N DEL 5
SRR1766459.5021042 chr5 27427137 N chr5 27427203 N DEL 5
SRR1766470.5375732 chr5 27427137 N chr5 27427203 N DEL 5
SRR1766453.3549622 chr5 27427137 N chr5 27427203 N DEL 5
SRR1766449.719669 chr5 27427138 N chr5 27427204 N DEL 4
SRR1766448.8505674 chr5 27427141 N chr5 27427207 N DEL 1
SRR1766485.3875644 chr5 27427137 N chr5 27427227 N DEL 5
SRR1766473.4736452 chr5 27427131 N chr5 27427221 N DEL 5
SRR1766484.3401157 chr5 27427131 N chr5 27427221 N DEL 5
SRR1766469.10408934 chr5 27427137 N chr5 27427227 N DEL 5
SRR1766470.2705063 chr5 27427137 N chr5 27427227 N DEL 5
SRR1766450.10523635 chr5 27427134 N chr5 27427224 N DEL 5
SRR1766485.8228915 chr5 27427137 N chr5 27427227 N DEL 5
SRR1766446.9324842 chr5 27427136 N chr5 27427226 N DEL 5
SRR1766451.2386677 chr5 27427137 N chr5 27427227 N DEL 5
SRR1766460.1967473 chr5 27427161 N chr5 27427234 N DEL 2
SRR1766465.11270907 chr5 27427137 N chr5 27427251 N DEL 5
SRR1766476.3753264 chr5 27427137 N chr5 27427251 N DEL 5
SRR1766457.981034 chr5 27427137 N chr5 27427251 N DEL 5
SRR1766455.5925878 chr5 27427162 N chr5 27427259 N DEL 1
SRR1766468.1654842 chr5 27427137 N chr5 27427275 N DEL 5
SRR1766485.4834032 chr5 27427137 N chr5 27427275 N DEL 5
SRR1766473.10254767 chr5 27427137 N chr5 27427275 N DEL 5
SRR1766477.6818586 chr5 27427137 N chr5 27427275 N DEL 5
SRR1766442.34427762 chr5 27427137 N chr5 27427275 N DEL 5
SRR1766467.11534793 chr5 27427138 N chr5 27427276 N DEL 4
SRR1766442.22299305 chr5 27427137 N chr5 27427299 N DEL 5
SRR1766460.3737794 chr5 27427137 N chr5 27427299 N DEL 5
SRR1766483.1789792 chr5 27427137 N chr5 27427299 N DEL 5
SRR1766452.956752 chr5 27427139 N chr5 27427301 N DEL 3
SRR1766472.10102489 chr18 79582411 N chr18 79582983 N DEL 4
SRR1766445.9257875 chr18 79582259 N chr18 79582434 N DEL 5
SRR1766454.2130715 chr18 79582727 N chr18 79582842 N DEL 7
SRR1766442.28059024 chr18 79582745 N chr18 79582856 N DUP 1
SRR1766472.4482790 chr18 79582668 N chr18 79582886 N DUP 3
SRR1766447.9487277 chr18 79582668 N chr18 79582886 N DUP 4
SRR1766452.2626559 chr18 79582668 N chr18 79582886 N DUP 4
SRR1766479.7682002 chr18 79582682 N chr18 79582902 N DEL 5
SRR1766449.6088393 chr16 34891886 N chr16 34891993 N DUP 5
SRR1766442.263812 chr1 189005976 N chr1 189006065 N DEL 5
SRR1766475.7203554 chr1 189005976 N chr1 189006065 N DEL 5
SRR1766475.4760898 chr1 103182937 N chr1 103183074 N DEL 8
SRR1766477.2851986 chr1 103183005 N chr1 103183074 N DEL 2
SRR1766458.524905 chr1 103183005 N chr1 103183074 N DEL 4
SRR1766453.522661 chr1 103183005 N chr1 103183074 N DEL 7
SRR1766481.8050794 chr1 103183005 N chr1 103183074 N DEL 7
SRR1766462.2887283 chr1 103183005 N chr1 103183074 N DEL 8
SRR1766481.8309394 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766478.9892453 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766469.8403513 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766484.11461911 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766471.7683050 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766466.10648705 chr1 103182937 N chr1 103183074 N DEL 5
SRR1766446.7103859 chr1 103182903 N chr1 103183074 N DEL 5
SRR1766442.34738564 chr1 103182903 N chr1 103183074 N DEL 5
SRR1766471.10708940 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766447.10788821 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766458.4102203 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766461.9033213 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766468.2323489 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766465.10276724 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766463.9579616 chr1 103182903 N chr1 103183074 N DEL 5
SRR1766446.7768499 chr1 103182903 N chr1 103183074 N DEL 5
SRR1766442.30073744 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766482.229753 chr1 103182903 N chr1 103183074 N DEL 5
SRR1766445.1783199 chr1 103182903 N chr1 103183074 N DEL 5
SRR1766443.7093167 chr1 103182903 N chr1 103183074 N DEL 5
SRR1766476.7013938 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766451.10333380 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766450.2528682 chr1 103182903 N chr1 103183074 N DEL 5
SRR1766442.42097907 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766443.2810271 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766445.3539154 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766456.6131194 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766467.4136555 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766471.6545430 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766475.3192630 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766449.7045159 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766468.868237 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766457.7278639 chr1 103183005 N chr1 103183074 N DEL 10
SRR1766463.5211377 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766455.6850370 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766472.2065535 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766460.10663906 chr1 103183005 N chr1 103183074 N DEL 7
SRR1766447.2095690 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766465.5582290 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766453.6555998 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766459.1904025 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766458.5732347 chr1 103182869 N chr1 103183074 N DEL 5
SRR1766446.3222093 chr1 103182835 N chr1 103183074 N DEL 5
SRR1766454.6967935 chr1 103182838 N chr1 103183077 N DEL 5
SRR1766460.1194443 chr1 103182838 N chr1 103183077 N DEL 5
SRR1766469.5283563 chr1 103182839 N chr1 103183078 N DEL 5
SRR1766477.6784770 chr1 103182847 N chr1 103183086 N DEL 3
SRR1766467.9357630 chr1 103182849 N chr1 103183088 N DEL 1
SRR1766486.1891716 chr20 45646267 N chr20 45646464 N DEL 5
SRR1766467.4330076 chr20 45646280 N chr20 45646360 N DEL 5
SRR1766446.2988704 chr22 38807555 N chr22 38807730 N DUP 5
SRR1766442.9410197 chr22 38807544 N chr22 38807769 N DUP 1
SRR1766476.10408718 chr22 38807534 N chr22 38807760 N DUP 8
SRR1766454.2991766 chr22 38807762 N chr22 38807890 N DEL 8
SRR1766467.1108090 chr22 38807715 N chr22 38807941 N DUP 10
SRR1766482.8769076 chr22 38807719 N chr22 38807947 N DUP 2
SRR1766483.7620423 chr22 38807642 N chr22 38807819 N DUP 2
SRR1766445.6245464 chr22 38807642 N chr22 38807819 N DUP 4
SRR1766453.10819496 chr22 38807642 N chr22 38807819 N DUP 5
SRR1766471.865666 chr22 38807515 N chr22 38807868 N DUP 5
SRR1766445.10478702 chr22 38807701 N chr22 38807802 N DEL 5
SRR1766445.8533467 chr14 56564609 N chr14 56564790 N DUP 1
SRR1766459.602651 chr1 175101910 N chr1 175102190 N DEL 5
SRR1766478.3190021 chr21 43975394 N chr21 43975447 N DUP 1
SRR1766442.42784834 chr10 92393378 N chr10 92393566 N DEL 5
SRR1766446.2492785 chr10 92393323 N chr10 92393556 N DEL 42
SRR1766474.1830864 chr10 92393338 N chr10 92393409 N DUP 5
SRR1766482.8824310 chr10 92393410 N chr10 92393509 N DUP 1
SRR1766481.11892151 chr10 92393343 N chr10 92393499 N DEL 6
SRR1766483.3971877 chr10 92393448 N chr10 92393539 N DEL 25
SRR1766446.10531661 chr10 92393448 N chr10 92393539 N DEL 19
SRR1766459.1943428 chr10 92393448 N chr10 92393539 N DEL 19
SRR1766460.416714 chr10 92393448 N chr10 92393539 N DEL 17
SRR1766442.15865456 chr10 92393404 N chr10 92393547 N DEL 7
SRR1766479.8012268 chr10 92393345 N chr10 92393555 N DEL 5
SRR1766468.3170598 chr10 92393398 N chr10 92393588 N DEL 4
SRR1766446.1919366 chr5 38821159 N chr5 38821251 N DUP 1
SRR1766471.11886399 chr5 38821159 N chr5 38821251 N DUP 2
SRR1766442.3553532 chr1 121836673 N chr1 121836942 N DEL 5
SRR1766458.4663378 chr1 121836673 N chr1 121836942 N DEL 5
SRR1766467.7524003 chr1 121836673 N chr1 121836942 N DEL 5
SRR1766443.4849970 chr1 121836673 N chr1 121836942 N DEL 5
SRR1766442.31762470 chr1 121836742 N chr1 121837011 N DEL 5
SRR1766460.5833895 chr1 121836742 N chr1 121837011 N DEL 5
SRR1766461.4623692 chr1 121836709 N chr1 121836976 N DUP 1
SRR1766483.10697640 chr1 121836807 N chr1 121837076 N DEL 5
SRR1766460.2117324 chr1 121836808 N chr1 121837075 N DUP 5
SRR1766480.5448552 chr1 121836808 N chr1 121837075 N DUP 5
SRR1766479.3045702 chr1 121836808 N chr1 121837075 N DUP 5
SRR1766457.5720111 chr1 121836808 N chr1 121837075 N DUP 5
SRR1766463.531716 chr1 121836891 N chr1 121837160 N DEL 1
SRR1766481.10808095 chr1 121836808 N chr1 121837075 N DUP 5
SRR1766461.10146253 chr1 121836808 N chr1 121837075 N DUP 5
SRR1766471.2645221 chr1 121836808 N chr1 121837075 N DUP 5
SRR1766465.6748128 chr1 121836808 N chr1 121837075 N DUP 5
SRR1766447.4733284 chr1 121836740 N chr1 121837007 N DUP 5
SRR1766452.5947986 chr1 121836740 N chr1 121837007 N DUP 5
SRR1766442.3553532 chr1 121836740 N chr1 121837007 N DUP 5
SRR1766458.4663378 chr1 121836740 N chr1 121837007 N DUP 5
SRR1766480.294430 chr1 121836740 N chr1 121837007 N DUP 5
SRR1766481.180414 chr1 121836740 N chr1 121837007 N DUP 5
SRR1766457.1502512 chr1 121836675 N chr1 121836944 N DEL 5
SRR1766471.7003000 chr2 217512943 N chr2 217513150 N DEL 5
SRR1766443.6371759 chr6 158155033 N chr6 158155130 N DEL 5
SRR1766479.6574 chr10 108880281 N chr10 108880339 N DUP 15
SRR1766442.39887904 chr10 108880281 N chr10 108880339 N DUP 16
SRR1766469.1876082 chr10 108880143 N chr10 108880352 N DEL 4
SRR1766461.10030268 chr10 108880297 N chr10 108880354 N DEL 3
SRR1766442.33690140 chr14 101245270 N chr14 101245325 N DEL 3
SRR1766468.7765869 chr14 101245272 N chr14 101245831 N DEL 5
SRR1766463.2446612 chr14 101245298 N chr14 101245911 N DEL 5
SRR1766469.5260493 chr14 101245308 N chr14 101245831 N DEL 5
SRR1766461.9158422 chr14 101245290 N chr14 101245651 N DEL 35
SRR1766470.10752330 chr14 101245334 N chr14 101245533 N DEL 5
SRR1766449.9274970 chr14 101245298 N chr14 101245911 N DEL 5
SRR1766481.6677747 chr14 101245334 N chr14 101245533 N DEL 5
SRR1766464.8372563 chr14 101245334 N chr14 101245533 N DEL 5
SRR1766484.5095045 chr14 101245334 N chr14 101245533 N DEL 5
SRR1766463.6114574 chr14 101245352 N chr14 101245911 N DEL 10
SRR1766463.10018286 chr14 101245362 N chr14 101245435 N DEL 5
SRR1766478.1825873 chr14 101245352 N chr14 101245911 N DEL 10
SRR1766465.9327965 chr14 101245352 N chr14 101245533 N DEL 15
SRR1766484.7439924 chr14 101245362 N chr14 101245435 N DEL 11
SRR1766452.2424098 chr14 101245344 N chr14 101245831 N DEL 14
SRR1766446.311057 chr14 101245939 N chr14 101246622 N DUP 28
SRR1766481.8432542 chr14 101245352 N chr14 101245911 N DEL 15
SRR1766460.4815622 chr14 101245373 N chr14 101246724 N DEL 27
SRR1766458.7111845 chr14 101245334 N chr14 101245425 N DEL 23
SRR1766468.7765869 chr14 101245356 N chr14 101245735 N DEL 24
SRR1766478.9702500 chr14 101245344 N chr14 101245831 N DEL 15
SRR1766446.420543 chr14 101245345 N chr14 101245544 N DEL 10
SRR1766471.3162563 chr14 101245217 N chr14 101245290 N DEL 5
SRR1766479.13375974 chr14 101245271 N chr14 101245324 N DUP 12
SRR1766443.5828807 chr14 101245271 N chr14 101245342 N DUP 16
SRR1766454.2135611 chr14 101245399 N chr14 101245904 N DEL 5
SRR1766462.1978821 chr14 101245345 N chr14 101245904 N DEL 15
SRR1766466.4792661 chr14 101245370 N chr14 101245821 N DEL 15
SRR1766470.1638359 chr14 101245345 N chr14 101245578 N DUP 10
SRR1766470.5716333 chr14 101245298 N chr14 101245533 N DEL 19
SRR1766453.879915 chr14 101245352 N chr14 101245911 N DEL 5
SRR1766462.5726561 chr14 101245219 N chr14 101245328 N DEL 9
SRR1766486.5168337 chr14 101245301 N chr14 101245444 N DUP 5
SRR1766485.4283071 chr14 101245423 N chr14 101245944 N DUP 15
SRR1766474.3378948 chr14 101245273 N chr14 101245902 N DUP 15
SRR1766486.5330697 chr14 101246382 N chr14 101246707 N DEL 20
SRR1766442.1229275 chr14 101245291 N chr14 101245902 N DUP 10
SRR1766443.8250472 chr14 101245452 N chr14 101245921 N DEL 5
SRR1766477.2479649 chr14 101245380 N chr14 101245883 N DUP 5
SRR1766485.359779 chr14 101245307 N chr14 101245380 N DEL 7
SRR1766467.8505432 chr14 101245307 N chr14 101245380 N DEL 5
SRR1766452.9003871 chr14 101245442 N chr14 101245821 N DEL 6
SRR1766470.1825605 chr14 101245273 N chr14 101245470 N DUP 14
SRR1766481.1297127 chr14 101245451 N chr14 101246100 N DEL 20
SRR1766450.7194758 chr14 101245332 N chr14 101245423 N DEL 13
SRR1766467.9106655 chr14 101245393 N chr14 101245446 N DUP 2
SRR1766483.9148776 chr14 101245964 N chr14 101246379 N DEL 20
SRR1766449.8007059 chr14 101245892 N chr14 101246379 N DEL 15
SRR1766482.5168333 chr14 101245478 N chr14 101245533 N DEL 25
SRR1766442.42666224 chr14 101245460 N chr14 101246379 N DEL 29
SRR1766444.5923801 chr14 101245496 N chr14 101245821 N DEL 24
SRR1766486.114319 chr14 101245460 N chr14 101246379 N DEL 31
SRR1766448.8377048 chr14 101245332 N chr14 101245423 N DEL 5
SRR1766465.1116988 chr14 101245308 N chr14 101245435 N DEL 15
SRR1766442.30835632 chr14 101245321 N chr14 101245518 N DUP 5
SRR1766445.1439541 chr14 101245327 N chr14 101245470 N DUP 25
SRR1766479.10761570 chr14 101245291 N chr14 101245506 N DUP 5
SRR1766484.2331466 chr14 101245281 N chr14 101245426 N DEL 14
SRR1766486.8858851 chr14 101245318 N chr14 101245515 N DUP 10
SRR1766446.2136184 chr14 101245290 N chr14 101245435 N DEL 13
SRR1766476.1774820 chr14 101245221 N chr14 101245438 N DEL 12
SRR1766476.339565 chr14 101245460 N chr14 101245533 N DEL 5
SRR1766442.30835632 chr14 101245536 N chr14 101246203 N DEL 15
SRR1766442.38613342 chr14 101245281 N chr14 101245532 N DUP 10
SRR1766462.2549889 chr14 101245282 N chr14 101245497 N DUP 7
SRR1766463.7734475 chr14 101245282 N chr14 101245497 N DUP 21
SRR1766466.8893021 chr14 101245303 N chr14 101246454 N DUP 13
SRR1766473.5689713 chr14 101245435 N chr14 101245542 N DUP 10
SRR1766460.8212328 chr14 101245496 N chr14 101245821 N DEL 14
SRR1766459.3519443 chr14 101245299 N chr14 101245480 N DEL 5
SRR1766462.8603687 chr14 101245548 N chr14 101246215 N DEL 10
SRR1766442.8271609 chr14 101245380 N chr14 101245577 N DUP 5
SRR1766452.3284318 chr14 101245597 N chr14 101245904 N DEL 3
SRR1766459.6957271 chr14 101245572 N chr14 101245717 N DEL 7
SRR1766479.13375974 chr14 101245453 N chr14 101245508 N DEL 10
SRR1766446.6671085 chr14 101245380 N chr14 101245577 N DUP 5
SRR1766454.599539 chr14 101245560 N chr14 101245939 N DEL 20
SRR1766447.5452777 chr14 101245435 N chr14 101245614 N DUP 10
SRR1766458.6651298 chr14 101245271 N chr14 101245558 N DUP 15
SRR1766484.333605 chr14 101245380 N chr14 101245577 N DUP 5
SRR1766465.11064262 chr14 101245273 N chr14 101245578 N DUP 16
SRR1766454.2135611 chr14 101246005 N chr14 101246708 N DEL 15
SRR1766442.15262427 chr14 101245221 N chr14 101245528 N DEL 10
SRR1766442.42286057 chr14 101245452 N chr14 101245543 N DEL 10
SRR1766445.4212652 chr14 101245591 N chr14 101245896 N DUP 15
SRR1766470.2488826 chr14 101245597 N chr14 101245904 N DEL 13
SRR1766471.10148455 chr14 101245292 N chr14 101245545 N DEL 3
SRR1766481.1297127 chr14 101245482 N chr14 101245591 N DEL 10
SRR1766462.3256831 chr14 101245496 N chr14 101245605 N DEL 5
SRR1766478.2367219 chr14 101245623 N chr14 101246864 N DUP 15
SRR1766478.9781159 chr14 101245597 N chr14 101245904 N DEL 20
SRR1766471.8152510 chr14 101245258 N chr14 101245311 N DUP 3
SRR1766478.6037459 chr14 101245362 N chr14 101245633 N DEL 25
SRR1766477.3098970 chr14 101245380 N chr14 101245451 N DUP 18
SRR1766442.5700407 chr14 101245533 N chr14 101245658 N DUP 15
SRR1766452.5029579 chr14 101245426 N chr14 101245695 N DUP 5
SRR1766484.5742455 chr14 101245282 N chr14 101245695 N DUP 1
SRR1766447.7848055 chr14 101245640 N chr14 101245821 N DEL 18
SRR1766442.21797007 chr14 101245640 N chr14 101246379 N DEL 5
SRR1766482.415829 chr14 101245636 N chr14 101245887 N DUP 20
SRR1766481.6398813 chr14 101245695 N chr14 101245768 N DEL 5
SRR1766470.1895312 chr14 101245318 N chr14 101245695 N DUP 20
SRR1766472.6341740 chr14 101245314 N chr14 101245621 N DEL 15
SRR1766485.8047111 chr14 101245314 N chr14 101245621 N DEL 15
SRR1766451.3254329 chr14 101245633 N chr14 101245686 N DUP 10
SRR1766450.4364560 chr14 101245358 N chr14 101245431 N DEL 10
SRR1766477.2542897 chr14 101245633 N chr14 101245884 N DUP 20
SRR1766463.5282942 chr14 101245623 N chr14 101245694 N DUP 15
SRR1766469.6404545 chr14 101245280 N chr14 101245623 N DEL 15
SRR1766477.1493530 chr14 101245308 N chr14 101245633 N DEL 20
SRR1766442.36906202 chr14 101245633 N chr14 101245686 N DUP 15
SRR1766478.7884671 chr14 101245672 N chr14 101246769 N DUP 6
SRR1766442.2944098 chr14 101245723 N chr14 101245904 N DEL 10
SRR1766452.2250233 chr14 101245274 N chr14 101245507 N DUP 15
SRR1766464.1808613 chr14 101245282 N chr14 101245713 N DUP 10
SRR1766471.9908205 chr14 101245464 N chr14 101245519 N DEL 5
SRR1766471.10588742 chr14 101245307 N chr14 101246100 N DEL 15
SRR1766486.7838220 chr14 101245297 N chr14 101245622 N DEL 5
SRR1766479.6759241 chr14 101245293 N chr14 101245654 N DEL 20
SRR1766449.1638059 chr14 101245722 N chr14 101246353 N DEL 5
SRR1766447.8209277 chr14 101245624 N chr14 101246829 N DUP 14
SRR1766455.449102 chr14 101245297 N chr14 101245640 N DEL 5
SRR1766470.8788501 chr14 101245464 N chr14 101245663 N DEL 5
SRR1766442.21797007 chr14 101245282 N chr14 101245713 N DUP 10
SRR1766453.6240820 chr14 101245273 N chr14 101245704 N DUP 20
SRR1766479.10761570 chr14 101245394 N chr14 101245665 N DEL 5
SRR1766450.7728881 chr14 101245516 N chr14 101245731 N DUP 5
SRR1766442.33690140 chr14 101245374 N chr14 101245717 N DEL 26
SRR1766458.3178253 chr14 101245282 N chr14 101245785 N DUP 5
SRR1766463.6114574 chr14 101245401 N chr14 101245726 N DEL 15
SRR1766486.6495742 chr14 101245706 N chr14 101245903 N DUP 10
SRR1766465.3000192 chr14 101245351 N chr14 101246738 N DEL 30
SRR1766458.7111845 chr14 101245598 N chr14 101245725 N DEL 5
SRR1766484.10457121 chr14 101245374 N chr14 101245735 N DEL 30
SRR1766446.1672006 chr14 101245309 N chr14 101245812 N DUP 10
SRR1766442.33696470 chr14 101245802 N chr14 101245911 N DEL 5
SRR1766454.7690490 chr14 101245281 N chr14 101245748 N DUP 15
SRR1766484.5382012 chr14 101245776 N chr14 101245831 N DEL 20
SRR1766447.9871520 chr14 101245370 N chr14 101245749 N DEL 26
SRR1766482.5168333 chr14 101245370 N chr14 101246487 N DEL 25
SRR1766459.8727129 chr14 101245289 N chr14 101245792 N DUP 15
SRR1766446.6468754 chr14 101245281 N chr14 101245732 N DEL 4
SRR1766464.8372563 chr14 101245352 N chr14 101245749 N DEL 10
SRR1766483.1597335 chr14 101245298 N chr14 101245749 N DEL 12
SRR1766454.2060420 chr14 101245767 N chr14 101245892 N DUP 14
SRR1766481.8432542 chr14 101245298 N chr14 101245749 N DEL 10
SRR1766446.6150418 chr14 101245298 N chr14 101246487 N DEL 15
SRR1766465.5700396 chr14 101245282 N chr14 101245785 N DUP 10
SRR1766457.8017718 chr14 101245310 N chr14 101245813 N DUP 5
SRR1766484.11203081 chr14 101245812 N chr14 101245921 N DEL 5
SRR1766442.10043082 chr14 101245812 N chr14 101245921 N DEL 5
SRR1766442.44680682 chr14 101245812 N chr14 101245921 N DEL 5
SRR1766482.6533115 chr14 101245785 N chr14 101245912 N DEL 5
SRR1766474.3378948 chr14 101245864 N chr14 101246639 N DEL 2
SRR1766478.9702500 chr14 101245864 N chr14 101246639 N DEL 5
SRR1766444.5923801 chr14 101245353 N chr14 101245786 N DEL 5
SRR1766452.3284318 chr14 101245504 N chr14 101245793 N DEL 5
SRR1766442.1229275 chr14 101245504 N chr14 101245793 N DEL 5
SRR1766446.6150418 chr14 101245829 N chr14 101246316 N DEL 10
SRR1766468.5097685 chr14 101245309 N chr14 101245902 N DUP 5
SRR1766478.1825873 chr14 101245488 N chr14 101245831 N DEL 20
SRR1766448.7476190 chr14 101245831 N chr14 101245884 N DUP 22
SRR1766481.5165580 chr14 101245317 N chr14 101245892 N DUP 22
SRR1766485.7749809 chr14 101245821 N chr14 101245892 N DUP 20
SRR1766478.11319565 chr14 101245293 N chr14 101245834 N DEL 20
SRR1766465.439369 chr14 101245317 N chr14 101245460 N DUP 10
SRR1766457.6100005 chr14 101245831 N chr14 101245884 N DUP 25
SRR1766454.8144665 chr14 101245298 N chr14 101245821 N DEL 15
SRR1766447.5452777 chr14 101245294 N chr14 101245817 N DEL 10
SRR1766467.2066155 chr14 101245823 N chr14 101246830 N DUP 11
SRR1766477.2321932 chr14 101245346 N chr14 101245527 N DEL 17
SRR1766481.10341623 chr14 101245290 N chr14 101245831 N DEL 13
SRR1766460.8212328 chr14 101245295 N chr14 101245836 N DEL 5
SRR1766466.4792661 chr14 101245352 N chr14 101246487 N DEL 19
SRR1766485.4283071 chr14 101245297 N chr14 101245838 N DEL 5
SRR1766466.10752342 chr14 101245333 N chr14 101246324 N DEL 10
SRR1766459.5305497 chr14 101245821 N chr14 101246036 N DUP 10
SRR1766479.9225617 chr14 101245291 N chr14 101245902 N DUP 5
SRR1766478.9074782 chr14 101245275 N chr14 101245886 N DUP 10
SRR1766463.10018286 chr14 101245271 N chr14 101245378 N DUP 18
SRR1766450.4428949 chr14 101245271 N chr14 101245378 N DUP 17
SRR1766453.6407873 chr14 101245274 N chr14 101245903 N DUP 10
SRR1766442.5693907 chr14 101245362 N chr14 101245453 N DEL 14
SRR1766473.5689713 chr14 101245271 N chr14 101245360 N DUP 10
SRR1766469.5260493 chr14 101245271 N chr14 101245378 N DUP 17
SRR1766462.2601057 chr14 101245279 N chr14 101245908 N DUP 10
SRR1766449.6654833 chr14 101245353 N chr14 101245786 N DEL 5
SRR1766453.6407873 chr14 101245496 N chr14 101245911 N DEL 15
SRR1766442.221807 chr14 101245579 N chr14 101245904 N DEL 5
SRR1766479.6506790 chr14 101245278 N chr14 101245349 N DUP 15
SRR1766449.9274970 chr14 101245586 N chr14 101245911 N DEL 10
SRR1766442.20819856 chr14 101245384 N chr14 101245889 N DEL 5
SRR1766486.1210980 chr14 101245370 N chr14 101245911 N DEL 15
SRR1766477.3098970 chr14 101245332 N chr14 101246089 N DEL 10
SRR1766463.3487261 chr14 101245887 N chr14 101246660 N DUP 5
SRR1766461.4940491 chr14 101245455 N chr14 101245888 N DEL 5
SRR1766454.7375551 chr14 101245271 N chr14 101245954 N DUP 10
SRR1766476.5417618 chr14 101245435 N chr14 101245992 N DUP 5
SRR1766478.6525055 chr14 101245281 N chr14 101245928 N DUP 9
SRR1766484.7439924 chr14 101245344 N chr14 101245939 N DEL 10
SRR1766450.7194758 chr14 101245425 N chr14 101245964 N DUP 15
SRR1766463.7734475 chr14 101245460 N chr14 101245911 N DEL 10
SRR1766449.9894398 chr14 101246000 N chr14 101246091 N DEL 5
SRR1766466.3621639 chr14 101245974 N chr14 101246101 N DEL 10
SRR1766449.1277676 chr14 101245831 N chr14 101245992 N DUP 19
SRR1766486.11512295 chr14 101245821 N chr14 101246000 N DUP 16
SRR1766454.599539 chr14 101245288 N chr14 101245919 N DEL 5
SRR1766450.8037774 chr14 101245317 N chr14 101245442 N DUP 12
SRR1766484.2565051 chr14 101245831 N chr14 101245992 N DUP 24
SRR1766450.2080379 chr14 101245487 N chr14 101246100 N DEL 20
SRR1766470.10752330 chr14 101245308 N chr14 101245939 N DEL 10
SRR1766442.5700407 chr14 101245362 N chr14 101245831 N DEL 22
SRR1766473.1702017 chr14 101245298 N chr14 101245929 N DEL 5
SRR1766484.7193371 chr14 101246136 N chr14 101246605 N DEL 25
SRR1766442.10000842 chr14 101245281 N chr14 101245948 N DEL 10
SRR1766483.4238392 chr14 101245974 N chr14 101246101 N DEL 10
SRR1766452.5029579 chr14 101245326 N chr14 101245939 N DEL 5
SRR1766469.1549462 chr14 101245289 N chr14 101245938 N DEL 5
SRR1766476.2111411 chr14 101245453 N chr14 101245884 N DUP 5
SRR1766442.19273876 chr14 101245285 N chr14 101245952 N DEL 2
SRR1766468.31014 chr14 101245271 N chr14 101245378 N DUP 15
SRR1766470.2488826 chr14 101245453 N chr14 101245884 N DUP 5
SRR1766464.1808613 chr14 101245217 N chr14 101245956 N DEL 5
SRR1766484.4202834 chr14 101245901 N chr14 101246010 N DEL 5
SRR1766445.7595154 chr14 101245901 N chr14 101246010 N DEL 5
SRR1766466.7587906 chr14 101245478 N chr14 101245533 N DEL 20
SRR1766462.8603687 chr14 101245901 N chr14 101246010 N DEL 5
SRR1766460.2051043 chr14 101245327 N chr14 101246046 N DUP 20
SRR1766443.11096063 chr14 101245308 N chr14 101245453 N DEL 14
SRR1766450.3353896 chr14 101245913 N chr14 101246074 N DUP 10
SRR1766442.38613342 chr14 101245865 N chr14 101246010 N DEL 7
SRR1766482.1173970 chr14 101246076 N chr14 101246707 N DEL 5
SRR1766484.333605 chr14 101246076 N chr14 101246707 N DEL 5
SRR1766442.42286057 chr14 101246076 N chr14 101246707 N DEL 5
SRR1766467.11787800 chr14 101245307 N chr14 101246010 N DEL 5
SRR1766459.6926832 chr14 101245307 N chr14 101246010 N DEL 5
SRR1766485.4558320 chr14 101246076 N chr14 101246707 N DEL 5
SRR1766465.11064262 chr14 101245536 N chr14 101246707 N DEL 10
SRR1766473.6728132 chr14 101245819 N chr14 101246088 N DUP 5
SRR1766443.6819343 chr14 101246087 N chr14 101246214 N DEL 15
SRR1766458.6651298 chr14 101245440 N chr14 101246017 N DEL 5
SRR1766470.396866 chr14 101246076 N chr14 101246473 N DEL 10
SRR1766464.937969 chr14 101245819 N chr14 101246088 N DUP 5
SRR1766442.10043082 chr14 101245857 N chr14 101246038 N DEL 5
SRR1766451.7085099 chr14 101245819 N chr14 101246088 N DUP 5
SRR1766479.11943828 chr14 101245819 N chr14 101246088 N DUP 10
SRR1766459.8727129 chr14 101245548 N chr14 101246089 N DEL 5
SRR1766479.9740464 chr14 101245631 N chr14 101246100 N DEL 5
SRR1766451.4681008 chr14 101245448 N chr14 101246061 N DEL 5
SRR1766455.5129217 chr14 101246163 N chr14 101246560 N DEL 10
SRR1766447.10219899 chr14 101245831 N chr14 101246136 N DUP 15
SRR1766446.2915964 chr14 101245831 N chr14 101246154 N DUP 30
SRR1766484.761616 chr14 101245307 N chr14 101246100 N DEL 10
SRR1766483.7188093 chr14 101245663 N chr14 101246130 N DUP 3
SRR1766483.10452952 chr14 101245433 N chr14 101246100 N DEL 5
SRR1766468.5097685 chr14 101245325 N chr14 101246100 N DEL 10
SRR1766445.1207403 chr14 101245460 N chr14 101246379 N DEL 15
SRR1766486.11512295 chr14 101246100 N chr14 101246603 N DUP 15
SRR1766470.1895312 chr14 101245325 N chr14 101246100 N DEL 10
SRR1766445.7569450 chr14 101245442 N chr14 101246379 N DEL 10
SRR1766463.4513275 chr14 101245946 N chr14 101246379 N DEL 15
SRR1766451.3372057 chr14 101245274 N chr14 101246173 N DUP 20
SRR1766459.3667085 chr14 101245433 N chr14 101246100 N DEL 5
SRR1766442.33696470 chr14 101245289 N chr14 101246100 N DEL 13
SRR1766470.396866 chr14 101245442 N chr14 101246379 N DEL 10
SRR1766464.6546876 chr14 101245442 N chr14 101246379 N DEL 10
SRR1766486.8692356 chr14 101245447 N chr14 101246114 N DEL 1
SRR1766484.5742455 chr14 101246110 N chr14 101246829 N DUP 5
SRR1766479.11989098 chr14 101245273 N chr14 101246172 N DUP 5
SRR1766484.2989722 chr14 101245271 N chr14 101245378 N DUP 15
SRR1766454.54597 chr14 101245497 N chr14 101246128 N DEL 5
SRR1766479.13146486 chr14 101245273 N chr14 101246172 N DUP 5
SRR1766459.5795576 chr14 101245371 N chr14 101246164 N DEL 5
SRR1766445.6693034 chr14 101245273 N chr14 101246172 N DUP 5
SRR1766445.9123263 chr14 101246109 N chr14 101246216 N DUP 2
SRR1766471.9908205 chr14 101245579 N chr14 101246174 N DEL 10
SRR1766477.7198085 chr14 101245717 N chr14 101246238 N DUP 5
SRR1766442.42250094 chr14 101245368 N chr14 101246215 N DEL 10
SRR1766459.424307 chr14 101245831 N chr14 101246226 N DUP 5
SRR1766458.3178253 chr14 101245318 N chr14 101245515 N DUP 10
SRR1766477.6589584 chr14 101245822 N chr14 101246217 N DUP 6
SRR1766466.3621639 chr14 101245316 N chr14 101246163 N DEL 5
SRR1766471.10486227 chr14 101245746 N chr14 101246215 N DEL 5
SRR1766471.3573507 chr14 101245896 N chr14 101246203 N DEL 20
SRR1766469.4685021 chr14 101245746 N chr14 101246215 N DEL 5
SRR1766453.6240820 chr14 101245587 N chr14 101246182 N DEL 15
SRR1766471.10486227 chr14 101245271 N chr14 101245756 N DUP 20
SRR1766470.7784038 chr14 101245590 N chr14 101246185 N DEL 7
SRR1766453.879915 chr14 101245694 N chr14 101246217 N DEL 15
SRR1766442.2944098 chr14 101245746 N chr14 101246215 N DEL 5
SRR1766442.44680682 chr14 101245767 N chr14 101246236 N DEL 5
SRR1766442.36720550 chr14 101246271 N chr14 101246540 N DUP 5
SRR1766457.8017718 chr14 101245370 N chr14 101246217 N DEL 16
SRR1766485.8742473 chr14 101245598 N chr14 101246193 N DEL 4
SRR1766485.980861 chr14 101245381 N chr14 101246244 N DUP 5
SRR1766479.5642890 chr14 101245299 N chr14 101246270 N DUP 20
SRR1766472.5230379 chr14 101245782 N chr14 101246251 N DEL 5
SRR1766463.4718845 chr14 101245904 N chr14 101246263 N DUP 5
SRR1766459.4420228 chr14 101246274 N chr14 101246707 N DEL 5
SRR1766449.6654833 chr14 101245296 N chr14 101246215 N DEL 10
SRR1766455.5129217 chr14 101245932 N chr14 101246473 N DEL 16
SRR1766477.1367445 chr14 101245321 N chr14 101246222 N DEL 5
SRR1766468.2840145 chr14 101245904 N chr14 101246281 N DUP 15
SRR1766456.3516764 chr14 101245819 N chr14 101246286 N DUP 8
SRR1766475.10583976 chr14 101245717 N chr14 101246346 N DUP 5
SRR1766477.6709766 chr14 101245327 N chr14 101246298 N DUP 10
SRR1766461.3588899 chr14 101245334 N chr14 101246289 N DEL 10
SRR1766482.4872556 chr14 101245821 N chr14 101246306 N DUP 19
SRR1766486.5168337 chr14 101245525 N chr14 101245902 N DUP 20
SRR1766453.10345893 chr14 101245821 N chr14 101246306 N DUP 5
SRR1766452.9309309 chr14 101245273 N chr14 101246298 N DUP 20
SRR1766476.2111411 chr14 101245332 N chr14 101246287 N DEL 5
SRR1766449.5020930 chr14 101245334 N chr14 101245533 N DEL 10
SRR1766464.10117287 chr14 101245291 N chr14 101246352 N DUP 5
SRR1766466.8118570 chr14 101245911 N chr14 101246360 N DUP 5
SRR1766454.11030453 chr14 101245271 N chr14 101245468 N DUP 10
SRR1766457.7217813 chr14 101246101 N chr14 101246334 N DUP 25
SRR1766449.9894398 chr14 101245450 N chr14 101246279 N DEL 6
SRR1766454.7690490 chr14 101245314 N chr14 101246287 N DEL 10
SRR1766450.8366300 chr14 101245478 N chr14 101246217 N DEL 25
SRR1766484.6202096 chr14 101245451 N chr14 101246316 N DEL 5
SRR1766443.7847574 chr14 101245345 N chr14 101245452 N DUP 15
SRR1766454.7375551 chr14 101245451 N chr14 101246316 N DEL 5
SRR1766484.5382012 chr14 101245300 N chr14 101246291 N DEL 10
SRR1766478.9972357 chr14 101245911 N chr14 101246360 N DUP 5
SRR1766460.1657224 chr14 101245273 N chr14 101246352 N DUP 20
SRR1766451.3254329 chr14 101245326 N chr14 101246317 N DEL 17
SRR1766475.8846686 chr14 101245344 N chr14 101246317 N DEL 19
SRR1766442.5693907 chr14 101245451 N chr14 101246316 N DEL 5
SRR1766453.4744671 chr14 101245451 N chr14 101246316 N DEL 5
SRR1766478.10684306 chr14 101246100 N chr14 101246387 N DUP 5
SRR1766475.1637672 chr14 101245831 N chr14 101246280 N DUP 20
SRR1766486.10137409 chr14 101245443 N chr14 101246326 N DEL 5
SRR1766478.5042180 chr14 101245642 N chr14 101246433 N DUP 3
SRR1766475.10583976 chr14 101245866 N chr14 101246101 N DEL 20
SRR1766456.3516764 chr14 101245478 N chr14 101246379 N DEL 15
SRR1766457.6100005 chr14 101245496 N chr14 101246379 N DEL 10
SRR1766461.4449336 chr14 101245295 N chr14 101246376 N DEL 4
SRR1766454.6052678 chr14 101245298 N chr14 101246379 N DEL 8
SRR1766468.6715708 chr14 101245283 N chr14 101246452 N DUP 15
SRR1766448.10853759 chr14 101245831 N chr14 101246460 N DUP 5
SRR1766476.8860572 chr14 101245282 N chr14 101246451 N DUP 5
SRR1766471.7528543 chr14 101245290 N chr14 101246011 N DEL 10
SRR1766482.4872556 chr14 101245273 N chr14 101245902 N DUP 10
SRR1766464.2378079 chr14 101245889 N chr14 101246178 N DEL 10
SRR1766467.3866580 chr14 101246109 N chr14 101246720 N DUP 5
SRR1766443.7847574 chr14 101246119 N chr14 101246226 N DUP 5
SRR1766463.4433866 chr14 101245353 N chr14 101246434 N DEL 5
SRR1766473.6728132 chr14 101245452 N chr14 101246425 N DEL 10
SRR1766449.1277676 chr14 101245998 N chr14 101246485 N DEL 25
SRR1766443.11096063 chr14 101245704 N chr14 101246335 N DEL 5
SRR1766475.8846686 chr14 101245533 N chr14 101245766 N DUP 6
SRR1766448.7476190 chr14 101245299 N chr14 101246434 N DEL 5
SRR1766485.7749809 chr14 101245548 N chr14 101246485 N DEL 5
SRR1766464.8365604 chr14 101245452 N chr14 101246425 N DEL 5
SRR1766479.5642890 chr14 101245579 N chr14 101246444 N DEL 10
SRR1766476.3644173 chr14 101245332 N chr14 101246449 N DEL 5
SRR1766477.11449956 chr14 101245793 N chr14 101246260 N DUP 2
SRR1766486.699950 chr14 101245299 N chr14 101246452 N DEL 20
SRR1766450.8037774 chr14 101245793 N chr14 101246260 N DUP 5
SRR1766479.9225617 chr14 101245453 N chr14 101246444 N DEL 10
SRR1766458.7379630 chr14 101245793 N chr14 101246260 N DUP 5
SRR1766442.704320 chr14 101245350 N chr14 101246485 N DEL 30
SRR1766482.4051031 chr14 101245793 N chr14 101246260 N DUP 5
SRR1766442.42250094 chr14 101245692 N chr14 101246485 N DEL 15
SRR1766445.9123263 chr14 101245793 N chr14 101246260 N DUP 5
SRR1766481.11495774 chr14 101245314 N chr14 101246485 N DEL 12
SRR1766486.4776314 chr14 101245921 N chr14 101246550 N DUP 10
SRR1766465.4071350 chr14 101245309 N chr14 101246550 N DUP 15
SRR1766457.5778614 chr14 101245680 N chr14 101246473 N DEL 6
SRR1766479.11943828 chr14 101245676 N chr14 101246487 N DEL 10
SRR1766444.5740043 chr14 101245328 N chr14 101246551 N DUP 15
SRR1766459.2447632 chr14 101245320 N chr14 101246473 N DEL 10
SRR1766461.10770513 chr14 101245271 N chr14 101246242 N DUP 23
SRR1766442.33647476 chr14 101245296 N chr14 101246485 N DEL 10
SRR1766460.1657224 chr14 101245289 N chr14 101246478 N DEL 5
SRR1766451.3372057 chr14 101245293 N chr14 101246482 N DEL 5
SRR1766442.36720550 chr14 101246281 N chr14 101246552 N DEL 15
SRR1766459.5305497 chr14 101245424 N chr14 101246487 N DEL 1
SRR1766469.9614842 chr14 101246295 N chr14 101246546 N DUP 10
SRR1766445.449651 chr14 101245423 N chr14 101246556 N DUP 5
SRR1766469.10123512 chr14 101246163 N chr14 101246542 N DEL 5
SRR1766447.7848055 chr14 101246163 N chr14 101246542 N DEL 5
SRR1766480.6181736 chr14 101246299 N chr14 101246552 N DEL 10
SRR1766459.8386373 chr14 101245370 N chr14 101246271 N DEL 5
SRR1766442.38014091 chr14 101246163 N chr14 101246542 N DEL 5
SRR1766461.7594490 chr14 101245865 N chr14 101246604 N DEL 10
SRR1766480.5941280 chr14 101245786 N chr14 101245965 N DUP 5
SRR1766473.784334 chr14 101245785 N chr14 101246542 N DEL 5
SRR1766451.7085099 chr14 101245759 N chr14 101246604 N DUP 2
SRR1766443.6819343 chr14 101245271 N chr14 101246638 N DUP 5
SRR1766477.6589584 chr14 101246570 N chr14 101246623 N DUP 16
SRR1766442.466758 chr14 101245471 N chr14 101246552 N DEL 10
SRR1766462.340158 chr14 101245322 N chr14 101246547 N DEL 5
SRR1766448.6487499 chr14 101245497 N chr14 101246542 N DEL 5
SRR1766465.7672721 chr14 101245281 N chr14 101246648 N DUP 5
SRR1766445.6693034 chr14 101245497 N chr14 101246542 N DEL 5
SRR1766445.449651 chr14 101245579 N chr14 101246552 N DEL 5
SRR1766461.3588899 chr14 101245667 N chr14 101246638 N DUP 5
SRR1766469.9614842 chr14 101245499 N chr14 101246544 N DEL 5
SRR1766452.9309309 chr14 101245579 N chr14 101246552 N DEL 5
SRR1766483.10452952 chr14 101245579 N chr14 101246552 N DEL 5
SRR1766485.980861 chr14 101245361 N chr14 101246604 N DEL 25
SRR1766450.3267099 chr14 101245502 N chr14 101246547 N DEL 5
SRR1766442.31600668 chr14 101245481 N chr14 101246580 N DEL 15
SRR1766465.4071350 chr14 101246559 N chr14 101246666 N DUP 20
SRR1766481.9721316 chr14 101245865 N chr14 101246604 N DEL 10
SRR1766462.2601057 chr14 101245496 N chr14 101246091 N DEL 20
SRR1766467.11302991 chr14 101245831 N chr14 101246570 N DEL 5
SRR1766459.424307 chr14 101245691 N chr14 101246610 N DEL 11
SRR1766481.7379630 chr14 101245831 N chr14 101246570 N DEL 5
SRR1766444.5740043 chr14 101245973 N chr14 101246604 N DEL 14
SRR1766485.11852955 chr14 101245291 N chr14 101246570 N DEL 13
SRR1766478.1274699 chr14 101245831 N chr14 101246570 N DEL 5
SRR1766461.7059478 chr14 101245832 N chr14 101246571 N DEL 5
SRR1766479.6506790 chr14 101245865 N chr14 101246604 N DEL 10
SRR1766460.2051043 chr14 101245296 N chr14 101246575 N DEL 5
SRR1766463.3487261 chr14 101245865 N chr14 101246604 N DEL 10
SRR1766457.7217813 chr14 101245361 N chr14 101246604 N DEL 13
SRR1766473.7540291 chr14 101245287 N chr14 101246584 N DEL 1
SRR1766477.6709766 chr14 101245287 N chr14 101246584 N DEL 1
SRR1766445.8922334 chr14 101245307 N chr14 101246604 N DEL 7
SRR1766442.8835869 chr14 101245307 N chr14 101246604 N DEL 5
SRR1766456.1886143 chr14 101245273 N chr14 101246676 N DUP 15
SRR1766483.7188093 chr14 101246100 N chr14 101246603 N DUP 15
SRR1766455.8583754 chr14 101246135 N chr14 101246782 N DUP 20
SRR1766452.6714314 chr14 101245533 N chr14 101246342 N DUP 10
SRR1766484.2565051 chr14 101245299 N chr14 101246632 N DEL 5
SRR1766442.38014091 chr14 101245796 N chr14 101246140 N DEL 6
SRR1766447.10219899 chr14 101245219 N chr14 101246642 N DEL 10
SRR1766484.7193371 chr14 101245920 N chr14 101246695 N DEL 10
SRR1766469.5943272 chr14 101245758 N chr14 101246731 N DEL 10
SRR1766466.8118570 chr14 101245464 N chr14 101246689 N DEL 20
SRR1766477.11449956 chr14 101245749 N chr14 101246738 N DUP 2
SRR1766457.6551052 chr14 101245749 N chr14 101246738 N DUP 5
SRR1766478.9972357 chr14 101245296 N chr14 101246701 N DEL 3
SRR1766464.937969 chr14 101245632 N chr14 101246497 N DEL 15
SRR1766467.5270396 chr14 101245302 N chr14 101246707 N DEL 5
SRR1766480.5941280 chr14 101245291 N chr14 101246714 N DEL 5
SRR1766475.10771606 chr14 101245921 N chr14 101246046 N DUP 20
SRR1766479.11989098 chr14 101245460 N chr14 101245749 N DEL 12
SRR1766484.962215 chr14 101245921 N chr14 101246802 N DUP 10
SRR1766450.8366300 chr14 101246440 N chr14 101246783 N DEL 5
SRR1766453.10345893 chr14 101246026 N chr14 101246819 N DEL 20
SRR1766456.1886143 chr14 101245828 N chr14 101246819 N DEL 5
SRR1766461.1928104 chr14 101245828 N chr14 101246819 N DEL 5
SRR1766486.4776314 chr14 101245828 N chr14 101246819 N DEL 5
SRR1766472.10525016 chr14 101245828 N chr14 101246819 N DEL 5
SRR1766444.6541026 chr14 101245828 N chr14 101246819 N DEL 5
SRR1766448.6738318 chr14 101245828 N chr14 101246819 N DEL 5
SRR1766483.5403524 chr14 101245828 N chr14 101246819 N DEL 5
SRR1766451.10639888 chr14 101245829 N chr14 101246820 N DEL 5
SRR1766454.4898158 chr14 101245831 N chr14 101246822 N DEL 5
SRR1766469.3868910 chr14 101245444 N chr14 101246831 N DEL 3
SRR1766486.1145252 chr14 101245285 N chr14 101246872 N DEL 8
SRR1766477.10855281 chr9 136894055 N chr9 136894353 N DEL 5
SRR1766467.763469 chr14 105570118 N chr14 105570233 N DUP 3
SRR1766470.10502638 chr14 105570234 N chr14 105570953 N DEL 5
SRR1766472.1116421 chr14 105570216 N chr14 105570792 N DEL 10
SRR1766447.6654874 chr14 105570186 N chr14 105570434 N DUP 5
SRR1766475.11117611 chr14 105570346 N chr14 105570562 N DEL 5
SRR1766475.5687126 chr14 105570250 N chr14 105570824 N DUP 1
SRR1766456.4720148 chr14 105570267 N chr14 105570755 N DUP 8
SRR1766484.11682379 chr14 105570373 N chr14 105570587 N DUP 5
SRR1766467.8234464 chr14 105570129 N chr14 105570397 N DEL 4
SRR1766474.235107 chr14 105570578 N chr14 105570810 N DEL 3
SRR1766442.1054140 chr14 105570516 N chr14 105570907 N DUP 2
SRR1766453.10683707 chr14 105570458 N chr14 105570671 N DUP 4
SRR1766471.9229233 chr14 105570250 N chr14 105570630 N DEL 3
SRR1766480.2697945 chr14 105570482 N chr14 105570693 N DEL 4
SRR1766457.9137224 chr14 105570133 N chr14 105570729 N DEL 10
SRR1766466.1836384 chr14 105570370 N chr14 105570752 N DEL 2
SRR1766472.10362227 chr14 105570232 N chr14 105570738 N DEL 5
SRR1766481.3077636 chr14 105570147 N chr14 105570875 N DUP 4
SRR1766454.2626927 chr14 105570233 N chr14 105570809 N DEL 3
SRR1766482.6252426 chrX 1561288 N chrX 1561403 N DUP 5
SRR1766483.5054508 chr7 154627144 N chr7 154627332 N DUP 5
SRR1766456.3758465 chr4 186043204 N chr4 186043271 N DEL 2
SRR1766442.5327475 chr4 186043172 N chr4 186043569 N DEL 1
SRR1766447.3878045 chr4 186043204 N chr4 186043337 N DEL 7
SRR1766475.8711322 chr4 186043172 N chr4 186043569 N DEL 5
SRR1766468.3116910 chr4 186043172 N chr4 186043569 N DEL 5
SRR1766477.6505316 chr4 186043172 N chr4 186043569 N DEL 5
SRR1766476.5271563 chr4 186043172 N chr4 186043569 N DEL 5
SRR1766476.10887086 chr4 186043259 N chr4 186043326 N DEL 5
SRR1766458.1776442 chr4 186043259 N chr4 186043326 N DEL 5
SRR1766464.7136723 chr4 186043601 N chr4 186043666 N DUP 15
SRR1766475.7816568 chr4 186043304 N chr4 186043437 N DEL 10
SRR1766463.7479151 chr4 186043282 N chr4 186043415 N DEL 5
SRR1766486.5801268 chr4 186043150 N chr4 186043415 N DEL 5
SRR1766486.4531391 chr4 186043305 N chr4 186043370 N DUP 5
SRR1766470.4585423 chr4 186043305 N chr4 186043370 N DUP 5
SRR1766465.9179805 chr4 186043305 N chr4 186043370 N DUP 5
SRR1766450.4459579 chr4 186043305 N chr4 186043370 N DUP 5
SRR1766460.5727324 chr4 186043348 N chr4 186043415 N DEL 3
SRR1766471.3322185 chr4 186043238 N chr4 186043305 N DEL 5
SRR1766456.868846 chr4 186043238 N chr4 186043305 N DEL 5
SRR1766460.4646960 chr4 186043238 N chr4 186043305 N DEL 5
SRR1766448.1811238 chr4 186043238 N chr4 186043305 N DEL 5
SRR1766483.11943886 chr4 186043238 N chr4 186043305 N DEL 5
SRR1766457.7558562 chr4 186043246 N chr4 186043313 N DEL 5
SRR1766467.3901981 chr4 186043348 N chr4 186043415 N DEL 5
SRR1766469.9994843 chr4 186043348 N chr4 186043415 N DEL 5
SRR1766483.1614004 chr4 186043348 N chr4 186043415 N DEL 5
SRR1766461.8856532 chr4 186043348 N chr4 186043415 N DEL 5
SRR1766467.5874479 chr4 186043437 N chr4 186043700 N DUP 10
SRR1766442.10113989 chr4 186043247 N chr4 186043314 N DEL 5
SRR1766452.4801303 chr4 186043181 N chr4 186043380 N DEL 5
SRR1766460.5895270 chr4 186043441 N chr4 186043704 N DUP 5
SRR1766472.1843896 chr4 186043415 N chr4 186043480 N DUP 5
SRR1766462.7205122 chr4 186043415 N chr4 186043480 N DUP 5
SRR1766463.3158830 chr4 186043518 N chr4 186043651 N DEL 10
SRR1766469.5299728 chr4 186043415 N chr4 186043480 N DUP 5
SRR1766479.5879682 chr4 186043415 N chr4 186043480 N DUP 5
SRR1766485.11424197 chr4 186043415 N chr4 186043480 N DUP 5
SRR1766476.9138369 chr4 186043415 N chr4 186043678 N DUP 6
SRR1766444.191234 chr4 186043321 N chr4 186043452 N DUP 3
SRR1766453.1447611 chr4 186043150 N chr4 186043415 N DEL 5
SRR1766442.1032264 chr4 186043150 N chr4 186043415 N DEL 5
SRR1766452.2571034 chr4 186043415 N chr4 186043480 N DUP 3
SRR1766467.8721292 chr4 186043284 N chr4 186043417 N DEL 5
SRR1766473.11820393 chr4 186043220 N chr4 186043419 N DEL 5
SRR1766474.10451272 chr4 186043220 N chr4 186043419 N DEL 5
SRR1766442.34808183 chr4 186043224 N chr4 186043423 N DEL 5
SRR1766443.8574927 chr4 186043415 N chr4 186043480 N DUP 5
SRR1766442.17837543 chr4 186043415 N chr4 186043480 N DUP 5
SRR1766442.30594265 chr4 186043188 N chr4 186043453 N DEL 5
SRR1766455.9305778 chr4 186043260 N chr4 186043523 N DUP 10
SRR1766462.6306000 chr4 186043259 N chr4 186043524 N DEL 10
SRR1766448.6935736 chr4 186043386 N chr4 186043651 N DEL 5
SRR1766481.5667782 chr4 186043408 N chr4 186043541 N DEL 5
SRR1766459.2494339 chr4 186043172 N chr4 186043633 N DUP 5
SRR1766454.3969859 chr4 186043123 N chr4 186043520 N DEL 5
SRR1766485.10524278 chr4 186043408 N chr4 186043541 N DEL 5
SRR1766462.2959477 chr4 186043541 N chr4 186043672 N DUP 6
SRR1766480.8697591 chr4 186043386 N chr4 186043585 N DEL 10
SRR1766480.8697591 chr4 186043144 N chr4 186043541 N DEL 7
SRR1766465.10926803 chr4 186043144 N chr4 186043541 N DEL 7
SRR1766471.8010748 chr4 186043145 N chr4 186043542 N DEL 5
SRR1766469.5666379 chr4 186043150 N chr4 186043547 N DEL 5
SRR1766442.20102227 chr4 186043151 N chr4 186043548 N DEL 5
SRR1766466.8060160 chr4 186043284 N chr4 186043549 N DEL 2
SRR1766477.3506960 chr4 186043415 N chr4 186043612 N DUP 5
SRR1766472.1101242 chr4 186043222 N chr4 186043553 N DEL 3
SRR1766445.2089099 chr4 186043601 N chr4 186043666 N DUP 5
SRR1766442.5327475 chr4 186043601 N chr4 186043666 N DUP 5
SRR1766448.1301692 chr4 186043601 N chr4 186043666 N DUP 5
SRR1766481.6339221 chr4 186043601 N chr4 186043666 N DUP 5
SRR1766465.2122427 chr4 186043601 N chr4 186043666 N DUP 5
SRR1766480.8671340 chr4 186043601 N chr4 186043666 N DUP 5
SRR1766477.660611 chr4 186043338 N chr4 186043603 N DEL 5
SRR1766461.906185 chr4 186043148 N chr4 186043611 N DEL 5
SRR1766481.704717 chr4 186043284 N chr4 186043615 N DEL 1
SRR1766479.6263200 chr4 186043259 N chr4 186043656 N DEL 5
SRR1766478.5566508 chr4 186043502 N chr4 186043701 N DEL 5
SRR1766473.10007304 chr4 186043127 N chr4 186043656 N DEL 5
SRR1766464.10779901 chr4 186043383 N chr4 186043714 N DEL 10
SRR1766478.8058522 chr4 186043370 N chr4 186043701 N DEL 5
SRR1766442.17802145 chr4 186043238 N chr4 186043701 N DEL 5
SRR1766477.6505316 chr4 186043651 N chr4 186043716 N DUP 5
SRR1766450.2393247 chr4 186043679 N chr4 186043746 N DEL 15
SRR1766461.7047770 chr4 186043704 N chr4 186043771 N DEL 8
SRR1766460.7700387 chr4 186043502 N chr4 186043767 N DEL 5
SRR1766479.6263200 chr4 186043481 N chr4 186043746 N DEL 5
SRR1766458.4194726 chr4 186043151 N chr4 186043746 N DEL 5
SRR1766453.10031499 chr4 186043151 N chr4 186043746 N DEL 5
SRR1766460.5727324 chr4 186043226 N chr4 186043755 N DEL 5
SRR1766477.5455519 chr2 60467224 N chr2 60467297 N DEL 5
SRR1766482.10171891 chr2 60467236 N chr2 60467870 N DEL 5
SRR1766470.690237 chr2 60467245 N chr2 60468161 N DEL 5
SRR1766471.1006136 chr2 60467226 N chr2 60467299 N DEL 5
SRR1766486.8748168 chr2 60467221 N chr2 60467274 N DUP 11
SRR1766443.7941489 chr2 60467221 N chr2 60467337 N DUP 15
SRR1766459.3145847 chr2 60467371 N chr2 60468065 N DEL 1
SRR1766462.608256 chr2 60467288 N chr2 60467476 N DUP 7
SRR1766471.5731134 chr2 60468151 N chr2 60468228 N DUP 13
SRR1766453.765743 chr2 60467238 N chr2 60467434 N DEL 5
SRR1766486.91312 chr2 60467296 N chr2 60467598 N DUP 12
SRR1766480.8030291 chr2 60467281 N chr2 60467583 N DUP 15
SRR1766471.1687300 chr2 60467307 N chr2 60467588 N DUP 16
SRR1766445.3464120 chr2 60467296 N chr2 60467598 N DUP 12
SRR1766474.7532084 chr2 60467296 N chr2 60467598 N DUP 20
SRR1766446.4705664 chr2 60467408 N chr2 60467617 N DUP 16
SRR1766480.4112742 chr2 60467297 N chr2 60467611 N DUP 21
SRR1766460.11092820 chr2 60467402 N chr2 60467605 N DUP 17
SRR1766465.2042980 chr2 60467297 N chr2 60467755 N DUP 18
SRR1766463.5695715 chr2 60467467 N chr2 60468083 N DEL 5
SRR1766458.1886098 chr2 60467291 N chr2 60467530 N DUP 20
SRR1766478.11860608 chr2 60467311 N chr2 60467744 N DEL 10
SRR1766450.4600800 chr2 60467335 N chr2 60467765 N DEL 12
SRR1766445.7527810 chr2 60467353 N chr2 60467825 N DEL 15
SRR1766459.3303569 chr2 60467347 N chr2 60467879 N DEL 23
SRR1766464.5980845 chr2 60467297 N chr2 60467920 N DUP 19
SRR1766458.1886098 chr2 60467335 N chr2 60467888 N DEL 7
SRR1766445.10213320 chr2 60467331 N chr2 60467893 N DEL 29
SRR1766458.3329846 chr2 60467869 N chr2 60468117 N DUP 5
SRR1766461.4846002 chr2 60467242 N chr2 60467879 N DEL 17
SRR1766481.10885226 chr2 60467555 N chr2 60467874 N DEL 10
SRR1766442.3002635 chr2 60467226 N chr2 60467966 N DUP 23
SRR1766459.7325521 chr2 60467275 N chr2 60467816 N DEL 15
SRR1766483.5691955 chr2 60467286 N chr2 60468019 N DEL 10
SRR1766452.7151758 chr2 60467332 N chr2 60468056 N DEL 18
SRR1766478.8676184 chr2 60467221 N chr2 60468156 N DUP 16
SRR1766442.3002635 chr2 60467938 N chr2 60468174 N DUP 8
SRR1766459.890083 chr2 60467244 N chr2 60468199 N DEL 10
SRR1766442.30954513 chr2 60467242 N chr2 60468227 N DEL 14
SRR1766443.7941489 chr2 60467314 N chr2 60468227 N DEL 10
SRR1766450.4837751 chr2 60467314 N chr2 60468272 N DEL 15
SRR1766482.10514975 chr2 60468190 N chr2 60468242 N DEL 13
SRR1766455.9636460 chr2 60467346 N chr2 60468262 N DEL 20
SRR1766465.7484885 chr2 60468192 N chr2 60468262 N DEL 15
SRR1766466.1387877 chr2 60467284 N chr2 60468293 N DEL 7
SRR1766485.3801890 chr2 60467256 N chr2 60468262 N DEL 10
SRR1766459.4304213 chr2 60467331 N chr2 60468271 N DEL 16
SRR1766443.871209 chr2 60467306 N chr2 60468261 N DEL 15
SRR1766484.770940 chr2 60467244 N chr2 60468271 N DEL 18
SRR1766455.3902386 chr2 60467241 N chr2 60468271 N DEL 15
SRR1766467.899119 chr2 60467313 N chr2 60468271 N DEL 15
SRR1766484.10722202 chr2 60467241 N chr2 60468271 N DEL 15
SRR1766461.4443736 chr2 60467268 N chr2 60468271 N DEL 10
SRR1766476.6936973 chr2 60467235 N chr2 60468280 N DEL 5
SRR1766466.4855412 chr2 60467237 N chr2 60468288 N DEL 5
SRR1766478.1923593 chr9 129339964 N chr9 129340017 N DEL 10
SRR1766465.1120521 chr17 402016 N chr17 402092 N DUP 4
SRR1766462.10869470 chr17 402031 N chr17 402137 N DEL 4
SRR1766480.2776584 chr17 402226 N chr17 402302 N DUP 21
SRR1766467.5644062 chr17 402067 N chr17 402276 N DUP 7
SRR1766457.1002041 chr17 402226 N chr17 402302 N DUP 12
SRR1766444.2198687 chr17 402226 N chr17 402302 N DUP 10
SRR1766477.1418828 chr17 402226 N chr17 402302 N DUP 12
SRR1766455.8706326 chr17 402226 N chr17 402302 N DUP 13
SRR1766442.31412096 chr17 402226 N chr17 402302 N DUP 5
SRR1766468.2771315 chr17 402032 N chr17 402215 N DEL 1
SRR1766454.1685749 chr17 402100 N chr17 402234 N DEL 5
SRR1766471.5429379 chr17 402105 N chr17 402239 N DEL 2
SRR1766476.1272960 chr17 402032 N chr17 402292 N DEL 1
SRR1766480.7803243 chr1 24804533 N chr1 24804663 N DEL 1
SRR1766450.6008615 chr1 24804506 N chr1 24804579 N DUP 5
SRR1766475.6046822 chr5 117993527 N chr5 117993580 N DEL 9
SRR1766480.219519 chr5 117993527 N chr5 117993580 N DEL 12
SRR1766446.1599666 chr5 117993527 N chr5 117993580 N DEL 13
SRR1766442.11850697 chr5 117993528 N chr5 117993579 N DUP 5
SRR1766482.11208196 chr5 117993528 N chr5 117993579 N DUP 5
SRR1766474.1092769 chr5 117993518 N chr5 117993589 N DUP 5
SRR1766475.10193603 chr5 117993542 N chr5 117993595 N DEL 5
SRR1766467.3757217 chr5 117993545 N chr5 117993598 N DEL 5
SRR1766452.4998773 chr5 117993533 N chr5 117993606 N DEL 2
SRR1766448.10222591 chr5 117993534 N chr5 117993607 N DEL 1
SRR1766448.3767833 chr12 120021332 N chr12 120021636 N DEL 18
SRR1766472.9005505 chr12 120021648 N chr12 120021967 N DEL 7
SRR1766442.47140745 chr12 120021396 N chr12 120021698 N DUP 5
SRR1766447.5736528 chr12 120021396 N chr12 120021698 N DUP 10
SRR1766461.520360 chr12 120021719 N chr12 120022038 N DEL 19
SRR1766469.6940271 chr12 120021794 N chr12 120021933 N DUP 5
SRR1766442.4211080 chr22 26736381 N chr22 26736598 N DEL 15
SRR1766442.4273459 chr22 26736302 N chr22 26736483 N DUP 7
SRR1766442.36074868 chr22 26736264 N chr22 26736315 N DEL 3
SRR1766445.10291832 chr22 26736384 N chr22 26736611 N DEL 2
SRR1766470.9377049 chr1 83013698 N chr1 83013789 N DEL 2
SRR1766449.7094048 chr1 83013731 N chr1 83013787 N DEL 10
SRR1766445.8204391 chr1 83013731 N chr1 83013787 N DEL 11
SRR1766461.2771859 chr1 83013731 N chr1 83013787 N DEL 17
SRR1766476.3864456 chr1 83013731 N chr1 83013787 N DEL 19
SRR1766479.8992341 chr1 83013731 N chr1 83013787 N DEL 16
SRR1766470.2374739 chr1 83013736 N chr1 83013787 N DEL 10
SRR1766446.372013 chr1 83013731 N chr1 83013787 N DEL 10
SRR1766453.9248675 chr1 83013731 N chr1 83013787 N DEL 10
SRR1766443.4637349 chr1 83013726 N chr1 83013787 N DEL 10
SRR1766460.158631 chr1 83013698 N chr1 83013789 N DEL 29
SRR1766483.9963672 chr1 83013698 N chr1 83013789 N DEL 22
SRR1766485.11030020 chr1 83013698 N chr1 83013789 N DEL 15
SRR1766459.10635134 chr1 83013696 N chr1 83013787 N DEL 10
SRR1766469.8401615 chr1 83013698 N chr1 83013789 N DEL 15
SRR1766445.4701610 chr1 83013699 N chr1 83013790 N DEL 14
SRR1766443.8533574 chr1 83013700 N chr1 83013791 N DEL 13
SRR1766447.7463113 chr1 83013692 N chr1 83013793 N DEL 9
SRR1766459.365250 chr1 83013702 N chr1 83013793 N DEL 11
SRR1766474.11263734 chr1 83013693 N chr1 83013794 N DEL 8
SRR1766474.5462463 chr1 83013691 N chr1 83013797 N DEL 5
SRR1766456.1324571 chr1 83013710 N chr1 83013801 N DEL 3
SRR1766479.4409 chr1 83013707 N chr1 83013798 N DEL 6
SRR1766481.7009359 chr1 83013705 N chr1 83013796 N DEL 8
SRR1766454.7842111 chr1 83013708 N chr1 83013799 N DEL 5
SRR1766481.8605274 chrY 11011510 N chrY 11012053 N DUP 9
SRR1766474.570502 chrY 11011521 N chrY 11011657 N DUP 4
SRR1766472.6607448 chr21 8594954 N chr21 8595147 N DEL 11
SRR1766469.3974505 chr21 8594830 N chr21 8594974 N DUP 5
SRR1766470.7905476 chr21 8595217 N chr21 8595535 N DUP 5
SRR1766483.10467820 chr20 60764300 N chr20 60764515 N DUP 7
SRR1766468.820543 chr20 60764378 N chr20 60764457 N DUP 5
SRR1766460.9789388 chr20 60764457 N chr20 60764538 N DEL 5
SRR1766461.8666817 chr20 60764457 N chr20 60764538 N DEL 5
SRR1766462.1890756 chr20 60764457 N chr20 60764538 N DEL 5
SRR1766450.8603136 chr20 60764373 N chr20 60764482 N DUP 3
SRR1766460.2096389 chr20 60764436 N chr20 60764519 N DEL 7
SRR1766474.9122601 chr20 60764417 N chr20 60764498 N DEL 4
SRR1766483.12242794 chr8 64541138 N chr8 64541252 N DUP 5
SRR1766466.7092978 chr3 180459351 N chr3 180459494 N DEL 14
SRR1766482.8331568 chr3 180459367 N chr3 180459488 N DEL 3
SRR1766472.5473560 chr3 180459367 N chr3 180459488 N DEL 5
SRR1766479.4414614 chr3 180459415 N chr3 180459474 N DUP 5
SRR1766453.10264664 chr3 180459385 N chr3 180459444 N DUP 5
SRR1766442.30257483 chr1 15036449 N chr1 15036530 N DEL 5
SRR1766462.1179863 chr18 21967845 N chr18 21967997 N DUP 2
SRR1766442.39549658 chr6 158156913 N chr6 158156992 N DUP 7
SRR1766472.3220974 chr6 158157004 N chr6 158157065 N DEL 5
SRR1766442.10052923 chr6 158157004 N chr6 158157065 N DEL 5
SRR1766464.2046669 chr6 158157029 N chr6 158157108 N DUP 27
SRR1766486.11838286 chr6 158157049 N chr6 158157128 N DUP 5
SRR1766479.2483755 chr4 174294811 N chr4 174294895 N DEL 5
SRR1766473.9689996 chr15 33794366 N chr15 33794465 N DUP 6
SRR1766482.10136339 chr11 1628484 N chr11 1628549 N DUP 5
SRR1766443.9991109 chr11 1628484 N chr11 1628549 N DUP 5
SRR1766482.8865151 chr11 1628507 N chr11 1628574 N DEL 5
SRR1766461.7677152 chr11 1628535 N chr11 1628602 N DEL 5
SRR1766486.1635450 chr11 1628543 N chr11 1628610 N DEL 4
SRR1766466.10561535 chr19 50592961 N chr19 50593124 N DUP 5
SRR1766481.3727346 chr19 50593037 N chr19 50593094 N DEL 5
SRR1766442.22539105 chr19 40648112 N chr19 40648416 N DEL 5
SRR1766468.6285405 chr19 40648112 N chr19 40648416 N DEL 5
SRR1766482.8956078 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766484.5274196 chr19 40648120 N chr19 40648248 N DEL 5
SRR1766477.8015887 chr19 40648275 N chr19 40648450 N DUP 8
SRR1766451.8007667 chr19 40648154 N chr19 40648281 N DEL 7
SRR1766485.8338926 chr19 40648405 N chr19 40648502 N DEL 1
SRR1766455.6815717 chr19 40648121 N chr19 40648423 N DUP 3
SRR1766483.852367 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766452.588469 chr19 40648121 N chr19 40648423 N DUP 4
SRR1766447.9964384 chr19 40648114 N chr19 40648416 N DUP 5
SRR1766451.4827711 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766442.22467875 chr19 40648154 N chr19 40648409 N DEL 10
SRR1766456.6473153 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766467.2760437 chr19 40648189 N chr19 40648395 N DEL 7
SRR1766479.7727327 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766456.4561087 chr19 40648148 N chr19 40648450 N DUP 7
SRR1766478.5219336 chr19 40648113 N chr19 40648464 N DUP 6
SRR1766469.1686096 chr19 40648188 N chr19 40648394 N DEL 10
SRR1766482.6107492 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766459.4715714 chr19 40648404 N chr19 40648454 N DUP 14
SRR1766458.8205420 chr19 40648188 N chr19 40648394 N DEL 8
SRR1766451.3828811 chr19 40648404 N chr19 40648453 N DUP 16
SRR1766452.6100915 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766480.5028797 chr19 40648367 N chr19 40648464 N DUP 4
SRR1766484.11505551 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766463.9590277 chr19 40648139 N chr19 40648394 N DEL 5
SRR1766442.10186378 chr19 40648144 N chr19 40648399 N DEL 5
SRR1766442.34330807 chr19 40648145 N chr19 40648400 N DEL 5
SRR1766482.7207997 chr21 31843707 N chr21 31843762 N DUP 6
SRR1766483.10682850 chr21 31843707 N chr21 31843762 N DUP 3
SRR1766485.747262 chr21 31843707 N chr21 31843864 N DUP 3
SRR1766486.11170137 chr21 31843773 N chr21 31843860 N DUP 2
SRR1766477.11245934 chr21 31843841 N chr21 31843900 N DEL 2
SRR1766444.439063 chr12 122164137 N chr12 122164432 N DEL 10
SRR1766454.5677670 chr12 122163820 N chr12 122164123 N DEL 25
SRR1766450.7478382 chr12 122163811 N chr12 122164114 N DEL 4
SRR1766442.23317080 chr12 122164225 N chr12 122164823 N DEL 5
SRR1766479.2295405 chr12 122163738 N chr12 122164347 N DEL 1
SRR1766472.9684518 chr12 122163894 N chr12 122164489 N DUP 5
SRR1766462.3675853 chr12 122163894 N chr12 122164489 N DUP 5
SRR1766481.4009502 chr12 122163921 N chr12 122164518 N DEL 5
SRR1766478.10481426 chr12 122163922 N chr12 122164519 N DEL 5
SRR1766453.4354999 chr12 122163923 N chr12 122164520 N DEL 5
SRR1766454.8471312 chr12 122163934 N chr12 122164531 N DEL 2
SRR1766467.6344911 chr12 122164356 N chr12 122164659 N DEL 5
SRR1766465.9132301 chr12 122164357 N chr12 122164660 N DEL 5
SRR1766465.11018805 chr12 122164148 N chr12 122164746 N DEL 15
SRR1766479.6732906 chr12 122164200 N chr12 122164798 N DEL 20
SRR1766479.2414300 chr12 122164485 N chr12 122164789 N DEL 3
SRR1766482.4763780 chr12 122164493 N chr12 122164797 N DEL 5
SRR1766484.6868641 chr12 122163921 N chr12 122164821 N DEL 5
SRR1766442.32874286 chr12 122164617 N chr12 122164921 N DEL 5
SRR1766475.7100167 chr9 9845155 N chr9 9845230 N DEL 24
SRR1766486.3963338 chr9 9845197 N chr9 9845270 N DEL 12
SRR1766465.9503357 chr9 9845167 N chr9 9845242 N DEL 27
SRR1766483.9943874 chr9 9845197 N chr9 9845270 N DEL 16
SRR1766445.1971641 chr9 9845167 N chr9 9845230 N DEL 53
SRR1766476.8604135 chr9 9845211 N chr9 9845282 N DUP 17
SRR1766444.4430820 chr19 2973963 N chr19 2974261 N DEL 15
SRR1766443.8289955 chr19 2974030 N chr19 2974328 N DEL 5
SRR1766442.44837182 chr19 2974059 N chr19 2974357 N DEL 10
SRR1766486.7149952 chr6 78554152 N chr6 78554238 N DEL 1
SRR1766457.6197943 chr6 78554080 N chr6 78554135 N DEL 15
SRR1766477.1164122 chr6 78554069 N chr6 78554201 N DEL 6
SRR1766470.5203252 chr6 78554078 N chr6 78554200 N DEL 10
SRR1766483.11966298 chr6 78554078 N chr6 78554200 N DEL 10
SRR1766458.3102470 chr1 143225344 N chr1 143225462 N DEL 2
SRR1766479.13507727 chr7 34129758 N chr7 34129809 N DEL 22
SRR1766479.9531288 chr12 14179718 N chr12 14179847 N DEL 11
SRR1766484.17580 chr12 14179718 N chr12 14179847 N DEL 13
SRR1766457.5758255 chr12 14179718 N chr12 14179847 N DEL 13
SRR1766471.11701813 chr12 14179718 N chr12 14179847 N DEL 16
SRR1766446.5787655 chr12 14179718 N chr12 14179927 N DEL 17
SRR1766481.11031130 chr12 14179718 N chr12 14179927 N DEL 17
SRR1766475.5335324 chr12 14179718 N chr12 14179927 N DEL 17
SRR1766459.2640871 chr12 14179710 N chr12 14179759 N DUP 5
SRR1766461.8184172 chr12 14179711 N chr12 14179760 N DUP 4
SRR1766471.5341137 chr12 14179750 N chr12 14179989 N DUP 24
SRR1766470.1907208 chr12 14179750 N chr12 14179989 N DUP 24
SRR1766443.1479011 chr12 14179750 N chr12 14179989 N DUP 24
SRR1766454.8804235 chr12 14179674 N chr12 14179763 N DEL 2
SRR1766476.5757908 chr12 14179674 N chr12 14179763 N DEL 2
SRR1766465.2315672 chr12 14179675 N chr12 14179764 N DEL 1
SRR1766442.36783829 chr12 14179755 N chr12 14179873 N DUP 10
SRR1766481.1898537 chr12 14179756 N chr12 14179874 N DUP 9
SRR1766454.5363561 chr12 14179673 N chr12 14179879 N DEL 9
SRR1766442.28786137 chr22 48535707 N chr22 48535944 N DEL 5
SRR1766455.4348564 chr22 48535736 N chr22 48535841 N DUP 5
SRR1766475.10600698 chr12 132644816 N chr12 132644926 N DEL 5
SRR1766481.4181059 chr12 132644816 N chr12 132645089 N DEL 5
SRR1766450.7327889 chr12 132644836 N chr12 132645109 N DEL 3
SRR1766472.4310454 chr12 132645438 N chr12 132645498 N DEL 5
SRR1766463.9554293 chr15 97641268 N chr15 97641333 N DUP 28
SRR1766464.1175433 chr15 97641268 N chr15 97641333 N DUP 34
SRR1766471.8616447 chr15 97641149 N chr15 97641281 N DEL 7
SRR1766461.10816161 chr15 97641268 N chr15 97641333 N DUP 28
SRR1766459.5931635 chr15 97641268 N chr15 97641333 N DUP 30
SRR1766442.22567980 chr15 97641268 N chr15 97641333 N DUP 29
SRR1766460.9014412 chr7 67850050 N chr7 67850103 N DEL 10
SRR1766448.2491011 chr16 65855214 N chr16 65855269 N DEL 9
SRR1766464.477532 chr16 65855210 N chr16 65855270 N DEL 9
SRR1766454.6465392 chr6 82306852 N chr6 82306941 N DUP 11
SRR1766468.2679719 chr6 82306901 N chr6 82306964 N DUP 4
SRR1766481.11944599 chr6 82306901 N chr6 82306964 N DUP 5
SRR1766476.4807001 chr6 82306901 N chr6 82306964 N DUP 5
SRR1766451.3054501 chr6 82306901 N chr6 82306964 N DUP 7
SRR1766446.9773451 chr6 82306901 N chr6 82306964 N DUP 7
SRR1766447.8341173 chr6 82306901 N chr6 82306964 N DUP 7
SRR1766442.9173826 chr6 82306888 N chr6 82307003 N DUP 6
SRR1766454.3230512 chr6 82306920 N chr6 82306999 N DEL 12
SRR1766476.262797 chr6 82306886 N chr6 82306979 N DEL 1
SRR1766444.1225838 chr6 82306996 N chr6 82307055 N DEL 24
SRR1766442.22455973 chr6 82306996 N chr6 82307055 N DEL 21
SRR1766458.6858572 chr6 82306996 N chr6 82307055 N DEL 17
SRR1766478.11040264 chr6 82306996 N chr6 82307055 N DEL 17
SRR1766459.11232537 chr6 82306998 N chr6 82307077 N DEL 22
SRR1766448.10210807 chr6 82306998 N chr6 82307077 N DEL 22
SRR1766450.10261164 chr6 82306998 N chr6 82307077 N DEL 16
SRR1766460.3745333 chr6 82306998 N chr6 82307077 N DEL 15
SRR1766458.3474171 chr6 82306998 N chr6 82307077 N DEL 15
SRR1766486.6220893 chr6 82306998 N chr6 82307077 N DEL 15
SRR1766463.5288650 chr6 82306998 N chr6 82307077 N DEL 15
SRR1766442.2917627 chr6 82306934 N chr6 82307077 N DEL 9
SRR1766482.1897071 chr6 82306870 N chr6 82307081 N DEL 9
SRR1766466.7120217 chr6 82306930 N chr6 82307085 N DEL 7
SRR1766483.2360211 chr6 82306930 N chr6 82307085 N DEL 7
SRR1766471.10027172 chr6 82306934 N chr6 82307089 N DEL 3
SRR1766458.121812 chr12 131327152 N chr12 131327394 N DEL 5
SRR1766480.2123825 chr12 131327152 N chr12 131327394 N DEL 20
SRR1766478.2037580 chr12 131327103 N chr12 131327197 N DUP 22
SRR1766442.10665047 chr12 131327200 N chr12 131327347 N DEL 25
SRR1766442.80768 chr12 131327113 N chr12 131327181 N DEL 12
SRR1766448.1114047 chr12 131327259 N chr12 131327412 N DUP 5
SRR1766442.40634523 chr12 131327259 N chr12 131327412 N DUP 5
SRR1766462.5869521 chr12 131327259 N chr12 131327412 N DUP 5
SRR1766471.11102652 chr12 131327259 N chr12 131327412 N DUP 7
SRR1766445.10269501 chr12 131327259 N chr12 131327412 N DUP 6
SRR1766462.4630555 chr12 131327262 N chr12 131327415 N DUP 5
SRR1766473.6267181 chr12 131327265 N chr12 131327509 N DUP 5
SRR1766476.5047474 chr12 131327273 N chr12 131327438 N DUP 1
SRR1766475.5524825 chr12 131327116 N chr12 131327283 N DEL 1
SRR1766464.9519003 chr12 131327322 N chr12 131327392 N DUP 10
SRR1766476.7566276 chr12 131327117 N chr12 131327347 N DEL 13
SRR1766479.7246577 chr12 131327115 N chr12 131327345 N DEL 11
SRR1766460.2898581 chr13 106570669 N chr13 106570798 N DEL 9
SRR1766481.10731177 chr13 106570720 N chr13 106570783 N DUP 12
SRR1766444.5142341 chr13 106570861 N chr13 106570926 N DEL 5
SRR1766486.1896406 chr12 132518400 N chr12 132519012 N DEL 16
SRR1766442.42557153 chr12 132518423 N chr12 132518984 N DEL 5
SRR1766484.838480 chr12 132518452 N chr12 132519081 N DEL 1
SRR1766448.5784507 chr12 132518545 N chr12 132519123 N DEL 6
SRR1766466.37776 chr12 132518545 N chr12 132519123 N DEL 2
SRR1766473.8056729 chr12 132518367 N chr12 132518618 N DUP 5
SRR1766476.9916818 chr12 132518635 N chr12 132518727 N DEL 15
SRR1766465.8884821 chr12 132518428 N chr12 132518559 N DEL 36
SRR1766466.8381570 chr12 132518425 N chr12 132518568 N DEL 5
SRR1766475.8014597 chr12 132518611 N chr12 132518697 N DUP 1
SRR1766442.28993338 chr12 132518366 N chr12 132518764 N DUP 5
SRR1766461.10326392 chr12 132518787 N chr12 132519035 N DEL 5
SRR1766462.730940 chr12 132518680 N chr12 132518803 N DUP 10
SRR1766445.1105087 chr12 132518791 N chr12 132519123 N DEL 3
SRR1766480.5461433 chr12 132518402 N chr12 132518825 N DUP 5
SRR1766474.1106232 chr12 132518845 N chr12 132518938 N DEL 5
SRR1766459.9457135 chr12 132518845 N chr12 132518938 N DEL 1
SRR1766467.1551428 chr12 132518888 N chr12 132519040 N DEL 2
SRR1766469.11181550 chr12 132518772 N chr12 132518919 N DUP 1
SRR1766480.5461433 chr12 132518382 N chr12 132519053 N DEL 2
SRR1766449.7997128 chr12 132518990 N chr12 132519078 N DEL 1
SRR1766450.6598247 chr12 132518554 N chr12 132519092 N DEL 6
SRR1766442.43092106 chr12 132518614 N chr12 132519081 N DEL 5
SRR1766471.8389706 chr12 132518554 N chr12 132519092 N DEL 5
SRR1766462.745909 chr12 132518381 N chr12 132519100 N DEL 5
SRR1766453.8694160 chr12 132518383 N chr12 132519102 N DEL 5
SRR1766459.9457135 chr12 132518383 N chr12 132519102 N DEL 5
SRR1766482.8161618 chr12 132518966 N chr12 132519110 N DEL 10
SRR1766464.7669897 chr12 132518429 N chr12 132519117 N DEL 2
SRR1766467.10119278 chr2 236491181 N chr2 236491278 N DUP 10
SRR1766484.159036 chr2 236491181 N chr2 236491278 N DUP 11
SRR1766463.1122541 chr2 236491181 N chr2 236491278 N DUP 15
SRR1766469.5767519 chr2 236491181 N chr2 236491278 N DUP 15
SRR1766449.8201656 chr2 236491182 N chr2 236491296 N DUP 9
SRR1766464.2476334 chrX 98534232 N chrX 98534439 N DUP 11
SRR1766453.8252410 chrX 98534236 N chrX 98534439 N DUP 16
SRR1766462.2133312 chrX 98534246 N chrX 98534427 N DEL 1
SRR1766446.5815091 chrX 98534246 N chrX 98534423 N DEL 5
SRR1766458.879567 chrX 98534246 N chrX 98534425 N DEL 3
SRR1766465.10704363 chr8 55767151 N chr8 55767254 N DEL 1
SRR1766446.333761 chr8 55767151 N chr8 55767254 N DEL 1
SRR1766470.2058358 chr8 55767151 N chr8 55767254 N DEL 7
SRR1766485.2906837 chr8 55767151 N chr8 55767254 N DEL 9
SRR1766476.3342286 chr8 55767151 N chr8 55767254 N DEL 9
SRR1766442.10833203 chr8 55767151 N chr8 55767254 N DEL 10
SRR1766476.1719770 chr8 55767157 N chr8 55767260 N DEL 9
SRR1766442.35291346 chr8 55767163 N chr8 55767266 N DEL 3
SRR1766449.1460827 chr8 55767162 N chr8 55767265 N DEL 4
SRR1766468.3036859 chr8 55767159 N chr8 55767262 N DEL 7
SRR1766485.10372490 chr8 55767153 N chr8 55767256 N DEL 13
SRR1766472.4325818 chr9 15456010 N chr9 15456322 N DEL 1
SRR1766452.10646644 chrX 121079468 N chrX 121079768 N DEL 30
SRR1766479.11126714 chr9 135261561 N chr9 135261730 N DEL 1
SRR1766451.5205665 chr9 135261540 N chr9 135261781 N DUP 8
SRR1766458.7750060 chr9 135261540 N chr9 135261799 N DUP 10
SRR1766457.3518584 chr9 135261530 N chr9 135261799 N DUP 16
SRR1766447.8367222 chr9 135261476 N chr9 135261695 N DEL 2
SRR1766484.810925 chr9 135261535 N chr9 135261724 N DEL 12
SRR1766474.6905791 chr9 135261557 N chr9 135261726 N DEL 13
SRR1766442.9227022 chr9 135261732 N chr9 135261901 N DUP 7
SRR1766457.1617167 chr9 135261730 N chr9 135261805 N DUP 13
SRR1766455.2612109 chr9 135261730 N chr9 135261805 N DUP 13
SRR1766482.2305095 chr9 135261785 N chr9 135261944 N DUP 10
SRR1766455.8088660 chr9 135261474 N chr9 135261805 N DEL 10
SRR1766442.22325825 chr9 135261789 N chr9 135261866 N DEL 5
SRR1766468.6985064 chr9 135261811 N chr9 135261926 N DEL 53
SRR1766466.6729179 chr8 142674091 N chr8 142674285 N DEL 5
SRR1766445.10085021 chr8 142674091 N chr8 142674349 N DEL 5
SRR1766471.7128650 chr8 142674091 N chr8 142674349 N DEL 5
SRR1766442.11925313 chr8 142674091 N chr8 142674285 N DEL 15
SRR1766485.10405025 chr8 142674142 N chr8 142674336 N DEL 5
SRR1766481.6060086 chr8 142674285 N chr8 142674476 N DUP 5
SRR1766448.8912749 chr8 142674043 N chr8 142674364 N DUP 5
SRR1766442.45888971 chr8 142674152 N chr8 142674410 N DEL 5
SRR1766471.7142470 chr8 142674126 N chr8 142674578 N DEL 5
SRR1766442.7315077 chr3 15163457 N chr3 15163578 N DEL 5
SRR1766458.9032698 chr3 15163738 N chr3 15163893 N DUP 10
SRR1766456.4792546 chr3 1642982 N chr3 1643037 N DEL 4
SRR1766466.9172648 chr3 1642982 N chr3 1643037 N DEL 4
SRR1766478.7631287 chr16 30232047 N chr16 30232357 N DEL 6
SRR1766442.46811603 chr7 36939434 N chr7 36939517 N DEL 15
SRR1766455.2933259 chr7 36939434 N chr7 36939517 N DEL 15
SRR1766446.2478883 chr7 36939434 N chr7 36939517 N DEL 15
SRR1766477.4994065 chr7 36939434 N chr7 36939517 N DEL 15
SRR1766450.5949375 chr7 36939437 N chr7 36939520 N DEL 12
SRR1766481.3332250 chr1 53502840 N chr1 53503219 N DUP 5
SRR1766443.3145251 chr3 180873619 N chr3 180873942 N DEL 5
SRR1766483.259294 chr3 180873904 N chr3 180874227 N DEL 20
SRR1766473.1629757 chr3 180873639 N chr3 180873955 N DEL 2
SRR1766465.7642744 chr14 57333969 N chr14 57334144 N DUP 1
SRR1766446.8867870 chr14 57333976 N chr14 57334199 N DUP 6
SRR1766467.8369505 chr14 57333977 N chr14 57334200 N DUP 7
SRR1766484.8893371 chr14 57333977 N chr14 57334200 N DUP 7
SRR1766446.2655250 chr14 57333977 N chr14 57334200 N DUP 7
SRR1766467.10259265 chr14 57333977 N chr14 57334200 N DUP 2
SRR1766460.1828266 chr14 57333977 N chr14 57334200 N DUP 7
SRR1766465.3412747 chr14 57333982 N chr14 57334159 N DEL 1
SRR1766459.2299868 chr14 57334001 N chr14 57334225 N DEL 7
SRR1766486.7469457 chr14 57334001 N chr14 57334225 N DEL 7
SRR1766464.7255279 chr14 57334004 N chr14 57334228 N DEL 7
SRR1766465.6489570 chr14 57334004 N chr14 57334228 N DEL 7
SRR1766448.7773376 chr14 57333966 N chr14 57334239 N DEL 1
SRR1766467.3163924 chr14 57334029 N chr14 57334302 N DEL 5
SRR1766473.5188916 chr14 57333986 N chr14 57334259 N DEL 5
SRR1766474.10249534 chr14 57334041 N chr14 57334361 N DUP 5
SRR1766463.8689934 chr14 57334029 N chr14 57334302 N DEL 5
SRR1766479.9832079 chr14 57333992 N chr14 57334314 N DEL 5
SRR1766457.3896388 chr11 70411321 N chr11 70411372 N DEL 5
SRR1766445.8306148 chr11 70411459 N chr11 70411558 N DUP 5
SRR1766443.1539947 chr17 5015511 N chr17 5015826 N DEL 5
SRR1766486.1814027 chr17 5015644 N chr17 5015957 N DEL 4
SRR1766462.2569474 chr22 23381270 N chr22 23381411 N DEL 15
SRR1766445.8498237 chr22 23381269 N chr22 23381413 N DEL 12
SRR1766447.2477157 chr22 23381269 N chr22 23381422 N DEL 8
SRR1766479.12909996 chr1 1056468 N chr1 1056549 N DUP 2
SRR1766485.7849889 chr1 1056492 N chr1 1056581 N DEL 11
SRR1766454.2754508 chr10 41755895 N chr10 41756753 N DEL 17
SRR1766477.2790073 chr10 41755791 N chr10 41756475 N DUP 9
SRR1766476.8508302 chr10 41755533 N chr10 41756390 N DEL 10
SRR1766442.42184993 chr7 14471315 N chr7 14471407 N DEL 13
SRR1766471.6389135 chr7 14471315 N chr7 14471407 N DEL 20
SRR1766476.4369637 chr7 14471315 N chr7 14471407 N DEL 21
SRR1766459.2282115 chr7 14471315 N chr7 14471407 N DEL 26
SRR1766449.8432411 chr7 14471315 N chr7 14471469 N DEL 28
SRR1766454.1892234 chr7 14471315 N chr7 14471407 N DEL 25
SRR1766472.6711196 chr7 14471315 N chr7 14471407 N DEL 28
SRR1766442.12888009 chr7 14471315 N chr7 14471407 N DEL 24
SRR1766465.5927457 chr7 14471315 N chr7 14471407 N DEL 24
SRR1766450.3889651 chr7 14471315 N chr7 14471407 N DEL 24
SRR1766449.7626711 chr7 14471405 N chr7 14471530 N DUP 13
SRR1766460.11116178 chr7 14471405 N chr7 14471530 N DUP 8
SRR1766452.4210058 chr7 14471363 N chr7 14471488 N DUP 5
SRR1766454.5217581 chr7 14471363 N chr7 14471488 N DUP 5
SRR1766462.3678965 chr7 14471363 N chr7 14471488 N DUP 5
SRR1766471.4483334 chr7 14471363 N chr7 14471488 N DUP 5
SRR1766478.10394420 chr7 14471363 N chr7 14471488 N DUP 9
SRR1766443.3601825 chr7 14471363 N chr7 14471488 N DUP 9
SRR1766477.6030305 chr7 14471363 N chr7 14471488 N DUP 9
SRR1766462.10289493 chr7 14471334 N chr7 14471484 N DUP 9
SRR1766469.4150726 chr7 14471405 N chr7 14471530 N DUP 14
SRR1766481.12693527 chr7 14471405 N chr7 14471530 N DUP 14
SRR1766442.15588503 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766442.37713788 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766449.1240833 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766464.10588109 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766442.40180803 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766483.78704 chr7 14471405 N chr7 14471530 N DUP 12
SRR1766448.7831943 chr7 14471405 N chr7 14471530 N DUP 11
SRR1766454.5217581 chr7 14471405 N chr7 14471530 N DUP 11
SRR1766468.2715767 chr7 14471405 N chr7 14471530 N DUP 11
SRR1766443.8829054 chr7 14471405 N chr7 14471530 N DUP 8
SRR1766442.24603183 chr7 14471405 N chr7 14471530 N DUP 7
SRR1766476.4369637 chr7 14471405 N chr7 14471530 N DUP 7
SRR1766481.5736519 chr7 14471405 N chr7 14471530 N DUP 6
SRR1766442.6617803 chr7 14471405 N chr7 14471530 N DUP 6
SRR1766454.1927364 chr7 14471405 N chr7 14471530 N DUP 6
SRR1766469.4150726 chr7 14471405 N chr7 14471530 N DUP 6
SRR1766474.6478355 chr7 14471405 N chr7 14471530 N DUP 6
SRR1766479.4962057 chr7 14471405 N chr7 14471530 N DUP 6
SRR1766442.38380606 chr7 14471405 N chr7 14471530 N DUP 9
SRR1766452.2303670 chr7 14471405 N chr7 14471530 N DUP 9
SRR1766455.8519310 chr7 14471405 N chr7 14471530 N DUP 10
SRR1766467.7874942 chr7 14471405 N chr7 14471530 N DUP 9
SRR1766442.9179734 chr7 14471405 N chr7 14471530 N DUP 10
SRR1766449.7626711 chr7 14471405 N chr7 14471530 N DUP 10
SRR1766482.2760425 chr7 14471405 N chr7 14471530 N DUP 10
SRR1766450.4623313 chr7 14471363 N chr7 14471519 N DUP 4
SRR1766453.7653212 chr7 14471363 N chr7 14471519 N DUP 4
SRR1766467.1006666 chr7 14471363 N chr7 14471519 N DUP 4
SRR1766442.31177757 chr7 14471363 N chr7 14471519 N DUP 4
SRR1766464.7190733 chr7 14471363 N chr7 14471488 N DUP 5
SRR1766478.2508733 chr7 14471363 N chr7 14471488 N DUP 5
SRR1766479.7195450 chr7 14471363 N chr7 14471488 N DUP 5
SRR1766465.668370 chr7 14471363 N chr7 14471488 N DUP 6
SRR1766445.5485293 chr7 14471363 N chr7 14471488 N DUP 7
SRR1766449.10057302 chr7 14471363 N chr7 14471488 N DUP 7
SRR1766452.9180670 chr7 14471363 N chr7 14471488 N DUP 8
SRR1766461.1746745 chr7 14471363 N chr7 14471488 N DUP 7
SRR1766469.354700 chr7 14471363 N chr7 14471488 N DUP 7
SRR1766458.1643637 chr7 14471363 N chr7 14471488 N DUP 7
SRR1766466.9488781 chr7 14471363 N chr7 14471488 N DUP 7
SRR1766472.4514954 chr7 14471363 N chr7 14471488 N DUP 8
SRR1766442.37686586 chr7 14471363 N chr7 14471488 N DUP 8
SRR1766454.1827730 chr7 14471333 N chr7 14471483 N DUP 9
SRR1766449.7449003 chr7 14471405 N chr7 14471466 N DUP 18
SRR1766467.11600466 chr7 14471405 N chr7 14471466 N DUP 18
SRR1766446.4336791 chr7 14471405 N chr7 14471466 N DUP 18
SRR1766486.11271527 chr7 14471405 N chr7 14471466 N DUP 18
SRR1766465.6965993 chr7 14471405 N chr7 14471466 N DUP 17
SRR1766442.4927756 chr7 14471405 N chr7 14471466 N DUP 17
SRR1766443.211294 chr7 14471405 N chr7 14471466 N DUP 17
SRR1766442.233973 chr7 14471405 N chr7 14471466 N DUP 19
SRR1766450.5102090 chr7 14471405 N chr7 14471466 N DUP 19
SRR1766451.3264428 chr7 14471388 N chr7 14471482 N DUP 3
SRR1766478.1819822 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766445.7708660 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766446.3770641 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766471.5303173 chr7 14471405 N chr7 14471466 N DUP 19
SRR1766471.7149905 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766477.9785768 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766442.44498754 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766450.1169239 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766447.8222869 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766448.9387396 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766442.2648806 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766462.5752283 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766479.9203479 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766442.12253223 chr7 14471409 N chr7 14471470 N DUP 10
SRR1766442.33750572 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766471.8974421 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766481.10609624 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766453.1051164 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766471.3005635 chr7 14471405 N chr7 14471530 N DUP 13
SRR1766472.4514954 chr7 14471405 N chr7 14471530 N DUP 13
SRR1766472.389000 chr7 14471405 N chr7 14471530 N DUP 11
SRR1766478.5212267 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766457.6265077 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766471.7205843 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766457.6265077 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766470.9529769 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766466.37817 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766442.25108929 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766443.6083702 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766458.7578535 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766466.8820409 chr7 14471410 N chr7 14471502 N DUP 4
SRR1766482.10852768 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766442.6585063 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766456.2489751 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766451.9708365 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766445.2585395 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766480.566338 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766459.1216777 chr7 14471405 N chr7 14471466 N DUP 14
SRR1766475.2836113 chr7 14471405 N chr7 14471466 N DUP 15
SRR1766444.1066160 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766464.709269 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766447.8222869 chr7 14471405 N chr7 14471466 N DUP 16
SRR1766474.3356550 chr7 14471405 N chr7 14471466 N DUP 17
SRR1766442.19631537 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766464.3823515 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766442.19519932 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766483.1302022 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766445.5578674 chr7 14471405 N chr7 14471466 N DUP 20
SRR1766466.5525349 chr17 72948383 N chr17 72948456 N DEL 5
SRR1766456.3903884 chr17 72948351 N chr17 72948460 N DEL 10
SRR1766477.10058285 chr17 72948351 N chr17 72948460 N DEL 10
SRR1766445.6756708 chr17 72948430 N chr17 72948501 N DUP 15
SRR1766448.5056434 chr17 72948430 N chr17 72948501 N DUP 15
SRR1766455.6281613 chr17 72948430 N chr17 72948501 N DUP 15
SRR1766454.7345606 chr17 72948360 N chr17 72948433 N DEL 10
SRR1766481.4109840 chr17 72948357 N chr17 72948430 N DEL 10
SRR1766481.1686056 chr17 72948447 N chr17 72948554 N DUP 16
SRR1766486.7688914 chr17 72948351 N chr17 72948460 N DEL 5
SRR1766475.207492 chr17 72948423 N chr17 72948496 N DEL 5
SRR1766483.9495277 chr17 72948351 N chr17 72948496 N DEL 5
SRR1766451.8959237 chr21 6572866 N chr21 6573009 N DUP 1
SRR1766461.5395640 chr21 6572952 N chr21 6573054 N DUP 1
SRR1766452.3967246 chr21 6573044 N chr21 6573208 N DUP 12
SRR1766486.611663 chr12 78626155 N chr12 78626288 N DUP 4
SRR1766446.8604918 chr12 78626224 N chr12 78626295 N DUP 5
SRR1766449.10137744 chr12 78626224 N chr12 78626295 N DUP 8
SRR1766442.8095465 chr12 78626252 N chr12 78626307 N DUP 41
SRR1766442.12445560 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766450.3138475 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766472.1700060 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766442.8815642 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766445.9892531 chr12 78626252 N chr12 78626307 N DUP 40
SRR1766465.3333568 chr12 78626252 N chr12 78626307 N DUP 31
SRR1766457.96031 chr12 78626209 N chr12 78626281 N DEL 8
SRR1766458.9440262 chr12 78626209 N chr12 78626281 N DEL 8
SRR1766454.1997453 chr12 78626167 N chr12 78626302 N DEL 2
SRR1766445.6536061 chr17 18000173 N chr17 18000510 N DEL 27
SRR1766460.10087069 chr17 18000232 N chr17 18000507 N DEL 5
SRR1766486.10994695 chr17 18000232 N chr17 18000507 N DEL 5
SRR1766444.6355246 chr17 18000246 N chr17 18000409 N DUP 2
SRR1766455.4172804 chr17 18000207 N chr17 18000322 N DEL 2
SRR1766443.4725037 chr17 18000135 N chr17 18000400 N DEL 6
SRR1766449.10657426 chr17 18000165 N chr17 18000440 N DEL 8
SRR1766445.9003251 chr4 1026160 N chr4 1026221 N DUP 5
SRR1766446.2399663 chr17 891852 N chr17 892000 N DEL 5
SRR1766448.4302868 chr17 891844 N chr17 892359 N DEL 5
SRR1766446.2399663 chr17 891839 N chr17 892061 N DEL 21
SRR1766447.8441910 chr17 891869 N chr17 892347 N DEL 5
SRR1766477.4840604 chr17 891869 N chr17 892347 N DEL 5
SRR1766455.7714545 chr17 891874 N chr17 892059 N DEL 15
SRR1766472.6656346 chr17 891869 N chr17 892347 N DEL 10
SRR1766476.4696548 chr17 891893 N chr17 892225 N DEL 20
SRR1766449.3386904 chr17 891911 N chr17 892059 N DEL 5
SRR1766467.2065900 chr17 891913 N chr17 892171 N DEL 8
SRR1766444.259232 chr17 891857 N chr17 892298 N DUP 10
SRR1766446.8638380 chr17 891857 N chr17 892298 N DUP 17
SRR1766466.10502257 chr17 891904 N chr17 892234 N DUP 15
SRR1766469.2128702 chr17 891913 N chr17 892245 N DEL 14
SRR1766482.11089384 chr17 891874 N chr17 892206 N DEL 20
SRR1766479.2204105 chr17 891911 N chr17 892243 N DEL 13
SRR1766459.2193542 chr17 891904 N chr17 892234 N DUP 20
SRR1766456.2639566 chr17 891911 N chr17 892169 N DEL 12
SRR1766465.506976 chr17 891911 N chr17 892169 N DEL 12
SRR1766467.2065900 chr17 891911 N chr17 892169 N DEL 12
SRR1766450.2402753 chr17 891904 N chr17 892308 N DUP 10
SRR1766459.11362980 chr17 891904 N chr17 892308 N DUP 10
SRR1766464.4980319 chr17 892044 N chr17 892301 N DUP 10
SRR1766481.1777112 chr17 891904 N chr17 892087 N DUP 10
SRR1766457.6004435 chr17 891904 N chr17 892087 N DUP 5
SRR1766453.7408944 chr17 891904 N chr17 892087 N DUP 2
SRR1766454.1479710 chr17 892000 N chr17 892146 N DUP 10
SRR1766472.6656346 chr17 892022 N chr17 892388 N DUP 10
SRR1766469.9795142 chr17 891889 N chr17 892037 N DEL 14
SRR1766448.298804 chr17 891874 N chr17 892022 N DEL 5
SRR1766463.6155510 chr17 892126 N chr17 892275 N DEL 1
SRR1766458.2659553 chr17 891874 N chr17 892022 N DEL 5
SRR1766462.1593302 chr17 891963 N chr17 892037 N DEL 5
SRR1766457.1900164 chr17 891889 N chr17 892037 N DEL 10
SRR1766457.2518149 chr17 891889 N chr17 892037 N DEL 9
SRR1766453.1936841 chr17 892059 N chr17 892279 N DUP 10
SRR1766471.4387627 chr17 892059 N chr17 892279 N DUP 10
SRR1766447.3659235 chr17 891984 N chr17 892169 N DEL 5
SRR1766481.11640892 chr17 892153 N chr17 892300 N DUP 6
SRR1766458.3689918 chr17 891911 N chr17 892169 N DEL 20
SRR1766451.6151269 chr17 891904 N chr17 892234 N DUP 19
SRR1766486.2786602 chr17 891911 N chr17 892169 N DEL 20
SRR1766458.9460395 chr17 892169 N chr17 892279 N DUP 9
SRR1766457.1900164 chr17 891857 N chr17 892407 N DUP 12
SRR1766479.8993410 chr17 892169 N chr17 892279 N DUP 9
SRR1766451.6151269 chr17 891913 N chr17 892171 N DEL 16
SRR1766478.11126503 chr17 892169 N chr17 892279 N DUP 8
SRR1766483.545019 chr17 891969 N chr17 892043 N DEL 5
SRR1766450.6126923 chr17 891911 N chr17 892132 N DEL 7
SRR1766483.545019 chr17 891874 N chr17 892169 N DEL 5
SRR1766445.3118856 chr17 891911 N chr17 892169 N DEL 7
SRR1766453.10977745 chr17 892169 N chr17 892279 N DUP 10
SRR1766442.25512711 chr17 891911 N chr17 892169 N DEL 10
SRR1766461.1441231 chr17 891913 N chr17 892171 N DEL 14
SRR1766461.9527350 chr17 891913 N chr17 892171 N DEL 9
SRR1766464.7682659 chr17 891913 N chr17 892171 N DEL 10
SRR1766482.2243559 chr17 891913 N chr17 892208 N DEL 23
SRR1766470.447434 chr17 891904 N chr17 892234 N DUP 15
SRR1766449.1953732 chr17 891913 N chr17 892208 N DEL 20
SRR1766471.2982393 chr17 891893 N chr17 892188 N DEL 10
SRR1766456.1177652 chr17 891913 N chr17 892208 N DEL 20
SRR1766467.4831609 chr17 891913 N chr17 892208 N DEL 20
SRR1766476.4130494 chr17 892169 N chr17 892279 N DUP 10
SRR1766449.2820829 chr17 891913 N chr17 892208 N DEL 17
SRR1766450.10697150 chr17 891983 N chr17 892168 N DEL 5
SRR1766476.3253926 chr17 892169 N chr17 892279 N DUP 12
SRR1766448.10050972 chr17 892206 N chr17 892279 N DUP 5
SRR1766448.10068846 chr17 892169 N chr17 892279 N DUP 10
SRR1766456.1177652 chr17 891857 N chr17 892407 N DUP 10
SRR1766478.7375151 chr17 892247 N chr17 892357 N DEL 5
SRR1766485.7399758 chr17 891899 N chr17 892266 N DUP 12
SRR1766449.10754332 chr17 891845 N chr17 892395 N DUP 18
SRR1766475.2602459 chr17 891857 N chr17 892298 N DUP 15
SRR1766474.643074 chr17 891913 N chr17 892171 N DEL 17
SRR1766478.7375151 chr17 892153 N chr17 892300 N DUP 9
SRR1766485.1754467 chr17 892206 N chr17 892279 N DUP 7
SRR1766477.5614973 chr17 892028 N chr17 892321 N DUP 3
SRR1766458.6587337 chr17 891893 N chr17 892188 N DEL 10
SRR1766482.11089384 chr17 891886 N chr17 892218 N DEL 3
SRR1766458.9446698 chr17 891873 N chr17 892351 N DEL 9
SRR1766476.4130494 chr17 891873 N chr17 892351 N DEL 4
SRR1766460.10169943 chr4 11191938 N chr4 11192036 N DUP 20
SRR1766471.8245417 chr4 11191909 N chr4 11191969 N DEL 4
SRR1766484.11932817 chr22 36773321 N chr22 36773612 N DUP 5
SRR1766456.2239798 chr1 1099172 N chr1 1099705 N DEL 7
SRR1766474.10199119 chr1 1099268 N chr1 1099573 N DEL 5
SRR1766470.2749836 chr1 1099279 N chr1 1099584 N DEL 4
SRR1766451.5850922 chr1 1099437 N chr1 1099743 N DEL 5
SRR1766476.3066512 chr1 1099533 N chr1 1099688 N DEL 5
SRR1766454.8643206 chr1 1099547 N chr1 1099933 N DEL 15
SRR1766478.11491471 chr1 1099543 N chr1 1099698 N DEL 9
SRR1766442.41952013 chr1 1099543 N chr1 1099698 N DEL 15
SRR1766468.4969712 chr1 1099204 N chr1 1099583 N DEL 5
SRR1766461.5696299 chr1 1099215 N chr1 1099594 N DEL 5
SRR1766461.7236831 chr1 1099652 N chr1 1099805 N DUP 5
SRR1766451.4446064 chr1 1099723 N chr1 1099799 N DUP 5
SRR1766442.36666099 chr1 1099724 N chr1 1099954 N DUP 5
SRR1766479.13677176 chr1 1099495 N chr1 1099878 N DUP 5
SRR1766483.2020511 chr1 1099416 N chr1 1099800 N DEL 5
SRR1766481.557565 chr1 1099217 N chr1 1099827 N DEL 10
SRR1766442.3712138 chr1 1099471 N chr1 1099856 N DEL 7
SRR1766455.509015 chr1 1099737 N chr1 1099894 N DEL 6
SRR1766485.9160462 chr1 1099659 N chr1 1099893 N DEL 5
SRR1766443.4364131 chr1 1099214 N chr1 1099978 N DEL 2
SRR1766442.19993263 chr22 11019419 N chr22 11019688 N DEL 1
SRR1766472.2696023 chr22 11019376 N chr22 11019510 N DUP 4
SRR1766477.6546779 chr22 11019582 N chr22 11019716 N DEL 3
SRR1766479.8885286 chr22 11019449 N chr22 11019673 N DEL 3
SRR1766479.1068764 chr22 11019451 N chr22 11019720 N DEL 10
SRR1766459.2454077 chr22 11019586 N chr22 11019720 N DEL 5
SRR1766478.8169319 chr22 11019528 N chr22 11019840 N DUP 6
SRR1766455.1570977 chr22 11019507 N chr22 11019776 N DEL 6
SRR1766486.10067306 chr22 11019436 N chr22 11019795 N DEL 5
SRR1766466.7557129 chr22 11019501 N chr22 11019815 N DEL 10
SRR1766474.11247388 chr13 71552931 N chr13 71552996 N DEL 9
SRR1766480.1168746 chr10 60240183 N chr10 60240269 N DEL 1
SRR1766482.8864026 chr10 60240183 N chr10 60240269 N DEL 4
SRR1766477.7922198 chr10 60240183 N chr10 60240269 N DEL 5
SRR1766443.193253 chr10 60240259 N chr10 60240368 N DEL 1
SRR1766479.7995816 chr10 60240259 N chr10 60240368 N DEL 5
SRR1766486.1121972 chr10 60240259 N chr10 60240368 N DEL 13
SRR1766477.8986785 chr10 60240259 N chr10 60240368 N DEL 13
SRR1766447.460340 chr10 60240162 N chr10 60240282 N DUP 31
SRR1766457.6485003 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766461.10565373 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766451.8173222 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766444.5590973 chr10 60240258 N chr10 60240359 N DUP 5
SRR1766443.2558803 chr10 60240271 N chr10 60240402 N DUP 20
SRR1766451.10459403 chr10 60240271 N chr10 60240402 N DUP 13
SRR1766474.7729092 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766442.20425156 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766467.6718301 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766466.3883400 chr10 60240205 N chr10 60240303 N DEL 14
SRR1766482.7427773 chr10 60240205 N chr10 60240303 N DEL 13
SRR1766483.3981936 chr10 60240174 N chr10 60240314 N DEL 4
SRR1766477.8457743 chr10 60240352 N chr10 60240433 N DEL 7
SRR1766451.8156767 chr10 60240352 N chr10 60240433 N DEL 7
SRR1766486.498212 chr10 60240352 N chr10 60240433 N DEL 7
SRR1766458.242909 chr10 60240355 N chr10 60240436 N DEL 7
SRR1766458.9353275 chr6 84395673 N chr6 84395739 N DUP 5
SRR1766463.3848720 chr6 84395673 N chr6 84395751 N DUP 14
SRR1766474.8263643 chr6 84395673 N chr6 84395755 N DUP 16
SRR1766470.2023851 chr6 84395673 N chr6 84395755 N DUP 18
SRR1766445.3886393 chr6 84395676 N chr6 84395762 N DUP 16
SRR1766451.9177715 chr6 84395676 N chr6 84395762 N DUP 17
SRR1766469.151355 chr6 84395673 N chr6 84395763 N DUP 19
SRR1766442.32666096 chr6 84395673 N chr6 84395763 N DUP 21
SRR1766467.11104608 chr6 84395673 N chr6 84395755 N DUP 21
SRR1766457.6306110 chr6 84395688 N chr6 84395740 N DEL 7
SRR1766453.6018346 chr6 84395688 N chr6 84395740 N DEL 7
SRR1766460.2538248 chr4 189362690 N chr4 189362782 N DEL 5
SRR1766462.7304708 chr9 134977402 N chr9 134977531 N DEL 5
SRR1766450.5024073 chr9 134977402 N chr9 134977531 N DEL 5
SRR1766470.2929213 chr9 134977402 N chr9 134977531 N DEL 5
SRR1766480.8475885 chr9 134977402 N chr9 134977531 N DEL 5
SRR1766483.436591 chr9 134977404 N chr9 134977461 N DEL 6
SRR1766479.1138542 chr9 134977404 N chr9 134977461 N DEL 7
SRR1766483.9951045 chr9 134977404 N chr9 134977461 N DEL 14
SRR1766482.5753684 chr9 134977404 N chr9 134977461 N DEL 14
SRR1766442.27305789 chr9 134977404 N chr9 134977461 N DEL 14
SRR1766442.8032591 chr9 134977404 N chr9 134977461 N DEL 15
SRR1766467.1904545 chr9 134977404 N chr9 134977461 N DEL 15
SRR1766459.3045532 chr9 134977404 N chr9 134977461 N DEL 10
SRR1766476.4309473 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766442.38469052 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766484.3894179 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766456.4700733 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766472.3604016 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766477.10974077 chr9 134977407 N chr9 134977460 N DUP 12
SRR1766442.43984930 chr9 134977411 N chr9 134977646 N DUP 14
SRR1766454.10726972 chr9 134977433 N chr9 134977492 N DUP 19
SRR1766450.9781022 chr9 134977469 N chr9 134977596 N DUP 12
SRR1766476.10816124 chr9 134977469 N chr9 134977596 N DUP 12
SRR1766467.4816567 chr9 134977469 N chr9 134977596 N DUP 11
SRR1766442.36274519 chr9 134977469 N chr9 134977596 N DUP 9
SRR1766473.4806751 chr9 134977469 N chr9 134977596 N DUP 9
SRR1766479.4540809 chr9 134977469 N chr9 134977596 N DUP 10
SRR1766456.3413997 chr9 134977405 N chr9 134977530 N DUP 13
SRR1766443.10493125 chr9 134977367 N chr9 134977438 N DEL 2
SRR1766479.1138542 chr9 134977367 N chr9 134977438 N DEL 2
SRR1766444.2707604 chr9 134977364 N chr9 134977435 N DEL 5
SRR1766449.419393 chr9 134977411 N chr9 134977506 N DUP 12
SRR1766475.9121539 chr9 134977411 N chr9 134977506 N DUP 11
SRR1766461.3935249 chr9 134977463 N chr9 134977518 N DUP 12
SRR1766473.1244817 chr9 134977421 N chr9 134977492 N DUP 15
SRR1766477.11513909 chr9 134977421 N chr9 134977492 N DUP 15
SRR1766472.5761640 chr9 134977463 N chr9 134977530 N DUP 9
SRR1766481.106377 chr9 134977523 N chr9 134977614 N DUP 10
SRR1766458.7090655 chr9 134977523 N chr9 134977614 N DUP 11
SRR1766442.9244279 chr9 134977523 N chr9 134977612 N DUP 14
SRR1766476.8526366 chr9 134977523 N chr9 134977614 N DUP 12
SRR1766471.1607677 chr9 134977523 N chr9 134977614 N DUP 12
SRR1766454.9679075 chr9 134977523 N chr9 134977614 N DUP 13
SRR1766450.6772662 chr9 134977523 N chr9 134977614 N DUP 16
SRR1766472.901242 chr9 134977487 N chr9 134977556 N DEL 8
SRR1766479.10286008 chr9 134977487 N chr9 134977556 N DEL 8
SRR1766458.6309674 chr9 134977517 N chr9 134977632 N DEL 26
SRR1766462.1830892 chr9 134977470 N chr9 134977543 N DEL 5
SRR1766451.8835524 chr9 134977472 N chr9 134977545 N DEL 3
SRR1766479.10617019 chr9 134977473 N chr9 134977546 N DEL 2
SRR1766457.3736435 chr9 134977474 N chr9 134977547 N DEL 1
SRR1766452.464242 chr9 134977411 N chr9 134977626 N DEL 12
SRR1766472.4740285 chr9 134977371 N chr9 134977656 N DEL 6
SRR1766453.5706830 chr9 134977369 N chr9 134977654 N DEL 8
SRR1766444.5978649 chr19 777117 N chr19 777428 N DEL 8
SRR1766470.3209460 chr19 777163 N chr19 777474 N DEL 7
SRR1766473.5794568 chrX 2426503 N chrX 2426597 N DUP 10
SRR1766481.8678663 chr13 46273699 N chr13 46274010 N DEL 5
SRR1766456.1717753 chr13 46273749 N chr13 46274059 N DEL 5
SRR1766443.1018008 chr13 46273755 N chr13 46274095 N DUP 4
SRR1766451.6830745 chr8 58301684 N chr8 58301733 N DUP 16
SRR1766442.14526898 chr8 58301684 N chr8 58301733 N DUP 20
SRR1766442.25935094 chr8 58301684 N chr8 58301733 N DUP 28
SRR1766448.3398217 chr8 58301684 N chr8 58301733 N DUP 28
SRR1766443.10652901 chr8 58301684 N chr8 58301733 N DUP 19
SRR1766480.1991184 chr7 77509639 N chr7 77509865 N DEL 5
SRR1766482.8928199 chr7 77509670 N chr7 77510072 N DEL 5
SRR1766449.3446824 chr7 77509527 N chr7 77509750 N DUP 6
SRR1766482.3660550 chr7 77509535 N chr7 77509758 N DUP 6
SRR1766447.2137512 chr7 77509655 N chr7 77509879 N DUP 3
SRR1766469.10863890 chr7 77509597 N chr7 77509772 N DUP 1
SRR1766477.10189725 chr7 77509785 N chr7 77509962 N DEL 5
SRR1766442.24163358 chr7 77509730 N chr7 77509954 N DUP 3
SRR1766445.6000549 chr7 77509785 N chr7 77509962 N DEL 5
SRR1766479.9885570 chr7 77509730 N chr7 77509954 N DUP 5
SRR1766473.7833850 chr7 77509564 N chr7 77509790 N DEL 5
SRR1766486.6686341 chr7 77509822 N chr7 77509999 N DEL 2
SRR1766481.2330565 chr7 77509614 N chr7 77509791 N DEL 5
SRR1766464.4347992 chr7 77509619 N chr7 77509796 N DEL 5
SRR1766470.3762676 chr7 77509575 N chr7 77509801 N DEL 4
SRR1766464.2183762 chr7 77509587 N chr7 77509813 N DEL 1
SRR1766465.8769954 chr7 77509620 N chr7 77509801 N DEL 3
SRR1766479.626894 chr7 77509939 N chr7 77510115 N DUP 12
SRR1766461.10855440 chr7 77509939 N chr7 77510117 N DUP 16
SRR1766482.3319426 chr7 77509927 N chr7 77510102 N DUP 5
SRR1766445.4718043 chr7 77509939 N chr7 77510115 N DUP 12
SRR1766476.7955973 chr7 77509939 N chr7 77510115 N DUP 12
SRR1766466.11084121 chr7 77509939 N chr7 77510115 N DUP 12
SRR1766449.2522181 chr7 77509615 N chr7 77509919 N DEL 5
SRR1766448.6608303 chr7 77509764 N chr7 77509941 N DEL 5
SRR1766467.1787340 chr7 77509763 N chr7 77509939 N DEL 12
SRR1766446.5200636 chr7 77509773 N chr7 77509948 N DUP 10
SRR1766452.4464855 chr7 77509577 N chr7 77509930 N DEL 2
SRR1766442.10292021 chr7 77509822 N chr7 77509997 N DUP 5
SRR1766464.5431306 chr7 77509822 N chr7 77509997 N DUP 5
SRR1766468.409704 chr7 77509783 N chr7 77510009 N DEL 5
SRR1766442.36807288 chr7 77509616 N chr7 77510018 N DEL 5
SRR1766476.9594236 chr7 77509618 N chr7 77510020 N DEL 5
SRR1766442.13327404 chr7 77509619 N chr7 77510021 N DEL 5
SRR1766469.632584 chr7 77509620 N chr7 77510022 N DEL 5
SRR1766476.9817073 chr7 77509624 N chr7 77510026 N DEL 4
SRR1766455.3347702 chr17 56898315 N chr17 56898373 N DEL 1
SRR1766486.6794350 chr17 56898315 N chr17 56898466 N DUP 1
SRR1766442.27260014 chr11 45588110 N chr11 45588167 N DEL 2
SRR1766459.8667019 chr11 45588113 N chr11 45588176 N DEL 9
SRR1766449.2303191 chr11 45588087 N chr11 45588184 N DEL 7
SRR1766484.330427 chr11 45588086 N chr11 45588183 N DEL 8
SRR1766486.544889 chr11 45588087 N chr11 45588188 N DEL 3
SRR1766479.2161934 chr11 45588082 N chr11 45588211 N DEL 3
SRR1766460.5931047 chr11 45588088 N chr11 45588225 N DEL 5
SRR1766467.7868723 chr20 61444434 N chr20 61444579 N DUP 15
SRR1766447.1403723 chr20 61444434 N chr20 61444579 N DUP 16
SRR1766442.37515660 chr20 61444633 N chr20 61444716 N DUP 12
SRR1766444.1083896 chr20 61444666 N chr20 61444795 N DUP 18
SRR1766471.336574 chr19 15896155 N chr19 15896233 N DEL 1
SRR1766466.9953406 chr12 51858512 N chr12 51858817 N DEL 35
SRR1766475.6592978 chr12 51858574 N chr12 51858879 N DEL 3
SRR1766477.8327567 chr12 51858574 N chr12 51858879 N DEL 9
SRR1766476.6227842 chr12 87486358 N chr12 87486539 N DUP 5
SRR1766445.2468416 chr12 87486378 N chr12 87486539 N DUP 5
SRR1766456.5230040 chr12 87486322 N chr12 87486497 N DEL 14
SRR1766480.7247295 chr12 87486623 N chr12 87486677 N DUP 2
SRR1766483.8940027 chr12 87486623 N chr12 87486677 N DUP 3
SRR1766473.7679145 chr12 87486623 N chr12 87486677 N DUP 5
SRR1766484.7758897 chr12 87486595 N chr12 87486699 N DUP 12
SRR1766483.1172379 chr12 87486595 N chr12 87486699 N DUP 14
SRR1766459.11229876 chr12 87486595 N chr12 87486699 N DUP 14
SRR1766478.10271732 chr17 76730846 N chr17 76730981 N DUP 5
SRR1766486.3784541 chr17 76730852 N chr17 76730987 N DUP 1
SRR1766478.6720795 chr17 76730882 N chr17 76731019 N DEL 5
SRR1766458.7245423 chr17 76730882 N chr17 76731019 N DEL 5
SRR1766484.8592923 chr17 76730882 N chr17 76731019 N DEL 5
SRR1766466.8102457 chr17 76730882 N chr17 76731019 N DEL 5
SRR1766473.6713226 chr17 76730882 N chr17 76731019 N DEL 5
SRR1766446.917799 chr17 117017 N chr17 117079 N DUP 1
SRR1766463.1025964 chr17 117017 N chr17 117079 N DUP 1
SRR1766472.585622 chr17 117026 N chr17 117088 N DUP 1
SRR1766442.7836089 chr17 117013 N chr17 117075 N DUP 5
SRR1766442.12307572 chr17 117016 N chr17 117078 N DUP 2
SRR1766442.26579927 chr17 117015 N chr17 117077 N DUP 3
SRR1766442.38429287 chr17 117021 N chr17 117083 N DUP 3
SRR1766442.43138181 chr17 117013 N chr17 117075 N DUP 5
SRR1766447.8646606 chr17 117014 N chr17 117076 N DUP 4
SRR1766448.4933956 chr17 117014 N chr17 117076 N DUP 4
SRR1766448.10548757 chr17 117013 N chr17 117075 N DUP 5
SRR1766449.3887275 chr17 117021 N chr17 117083 N DUP 3
SRR1766453.10031649 chr17 117014 N chr17 117076 N DUP 4
SRR1766469.1844224 chr17 117002 N chr17 117127 N DUP 5
SRR1766481.7421178 chr17 117014 N chr17 117076 N DUP 4
SRR1766485.4180038 chr17 117015 N chr17 117077 N DUP 3
SRR1766486.10958169 chr17 117014 N chr17 117076 N DUP 4
SRR1766450.10247396 chr17 117009 N chr17 117071 N DUP 9
SRR1766448.3667487 chr17 117002 N chr17 117064 N DUP 5
SRR1766446.708550 chr17 117002 N chr17 117127 N DUP 5
SRR1766486.9999513 chr17 117002 N chr17 117064 N DUP 5
SRR1766442.40423508 chr17 117016 N chr17 117078 N DUP 1
SRR1766450.1808541 chr17 117002 N chr17 117064 N DUP 5
SRR1766466.6696125 chr17 117002 N chr17 117127 N DUP 5
SRR1766480.616778 chr17 117002 N chr17 117064 N DUP 5
SRR1766466.3854198 chr17 117002 N chr17 117064 N DUP 5
SRR1766445.5830528 chr17 117002 N chr17 117127 N DUP 5
SRR1766455.7498866 chr17 117002 N chr17 117127 N DUP 5
SRR1766458.9120514 chr17 117041 N chr17 117166 N DUP 5
SRR1766455.8904017 chr17 117002 N chr17 117064 N DUP 5
SRR1766465.687207 chr17 117058 N chr17 117119 N DUP 6
SRR1766447.6125383 chr17 117002 N chr17 117064 N DUP 5
SRR1766469.8152124 chr17 117002 N chr17 117127 N DUP 5
SRR1766469.10739723 chr17 117002 N chr17 117127 N DUP 5
SRR1766442.6138361 chr17 117002 N chr17 117127 N DUP 5
SRR1766471.4863973 chr17 117002 N chr17 117064 N DUP 5
SRR1766461.7107936 chr17 117058 N chr17 117119 N DUP 6
SRR1766442.8690072 chr17 117002 N chr17 117127 N DUP 5
SRR1766479.11193786 chr17 117002 N chr17 117127 N DUP 5
SRR1766442.1078323 chr17 117005 N chr17 117067 N DUP 1
SRR1766442.27717286 chr17 117004 N chr17 117066 N DUP 1
SRR1766443.10460236 chr17 117002 N chr17 117127 N DUP 6
SRR1766450.2719519 chr17 117004 N chr17 117066 N DUP 1
SRR1766474.4643110 chr17 117012 N chr17 117074 N DUP 1
SRR1766451.296208 chr17 117003 N chr17 117065 N DUP 2
SRR1766454.3541988 chr17 117003 N chr17 117065 N DUP 2
SRR1766461.6733109 chr17 117002 N chr17 117064 N DUP 7
SRR1766467.3306149 chr17 117002 N chr17 117127 N DUP 7
SRR1766471.5886747 chr17 117003 N chr17 117065 N DUP 2
SRR1766473.3806109 chr17 117003 N chr17 117065 N DUP 2
SRR1766474.7519187 chr17 117003 N chr17 117065 N DUP 2
SRR1766474.9177738 chr17 117002 N chr17 117127 N DUP 7
SRR1766460.4589126 chr17 117005 N chr17 117067 N DUP 3
SRR1766478.8274980 chr17 117003 N chr17 117065 N DUP 4
SRR1766445.8632610 chr17 117003 N chr17 117065 N DUP 1
SRR1766461.7431562 chr17 117004 N chr17 117066 N DUP 5
SRR1766476.2581186 chr3 121313950 N chr3 121314338 N DUP 5
SRR1766443.8170998 chr3 121314047 N chr3 121314242 N DUP 1
SRR1766442.5518755 chr3 121314156 N chr3 121314313 N DEL 5
SRR1766447.9990920 chr3 121314222 N chr3 121314339 N DEL 5
SRR1766462.667741 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766460.6286345 chr5 59200731 N chr5 59200790 N DUP 6
SRR1766452.9972041 chr5 59200701 N chr5 59200790 N DUP 10
SRR1766443.7152936 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766475.10476939 chr5 59200731 N chr5 59200790 N DUP 9
SRR1766486.4593672 chr5 59200701 N chr5 59200790 N DUP 10
SRR1766461.8382651 chr5 59200701 N chr5 59200790 N DUP 10
SRR1766457.3375765 chr5 59200701 N chr5 59200790 N DUP 8
SRR1766462.1242708 chr5 59200701 N chr5 59200790 N DUP 8
SRR1766480.6926333 chr5 59200701 N chr5 59200790 N DUP 15
SRR1766463.4737383 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766447.5231820 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766482.11326733 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766451.2589525 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766448.7759843 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766480.546699 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766450.1008389 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766477.6197748 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766463.6770281 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766477.9405509 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766469.9516957 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766481.9091587 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766485.5767850 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766474.9484491 chr5 59200731 N chr5 59200790 N DUP 10
SRR1766442.39059137 chr5 59200731 N chr5 59200790 N DUP 7
SRR1766485.11871785 chr5 59200731 N chr5 59200790 N DUP 6
SRR1766442.20219007 chr5 59200731 N chr5 59200790 N DUP 6
SRR1766477.9111117 chr5 59200697 N chr5 59200820 N DEL 17
SRR1766480.4686596 chr5 59200697 N chr5 59200820 N DEL 17
SRR1766466.6670269 chr5 59200697 N chr5 59200820 N DEL 16
SRR1766469.1302346 chr5 59200760 N chr5 59200823 N DEL 7
SRR1766481.4230140 chr5 59200760 N chr5 59200823 N DEL 7
SRR1766455.3197651 chr5 59200761 N chr5 59200824 N DEL 6
SRR1766449.8115795 chr5 59200766 N chr5 59200829 N DEL 5
SRR1766481.5361701 chr12 32563453 N chr12 32563610 N DEL 9
SRR1766455.554550 chr12 32563551 N chr12 32563748 N DEL 2
SRR1766468.473946 chr12 32563311 N chr12 32563583 N DUP 5
SRR1766442.44843422 chr12 32563440 N chr12 32563595 N DUP 9
SRR1766475.8209660 chr12 32563470 N chr12 32563704 N DEL 5
SRR1766457.1037828 chr12 32563348 N chr12 32563738 N DEL 2
SRR1766448.4408527 chr15 78040755 N chr15 78041014 N DEL 14
SRR1766472.1655674 chr15 78040755 N chr15 78041014 N DEL 14
SRR1766485.3376636 chr15 78040755 N chr15 78041014 N DEL 14
SRR1766455.4618863 chr15 78040778 N chr15 78041043 N DUP 10
SRR1766459.1953392 chr15 78040781 N chr15 78041046 N DUP 2
SRR1766446.5872316 chr15 78040841 N chr15 78041007 N DEL 5
SRR1766480.1329959 chr15 78040814 N chr15 78041009 N DEL 5
SRR1766460.917143 chr15 78040814 N chr15 78041009 N DEL 5
SRR1766442.2802308 chr15 78040936 N chr15 78041010 N DEL 5
SRR1766484.2222749 chr15 78040814 N chr15 78041017 N DEL 3
SRR1766485.1411607 chr15 78040842 N chr15 78041040 N DEL 10
SRR1766478.3815893 chr15 78040751 N chr15 78041046 N DEL 7
SRR1766469.4516228 chr1 232572826 N chr1 232572933 N DEL 5
SRR1766446.7288313 chr10 59696922 N chr10 59697003 N DEL 2
SRR1766468.2460452 chr10 59697159 N chr10 59697288 N DEL 1
SRR1766467.8985814 chr10 59697159 N chr10 59697288 N DEL 3
SRR1766468.2460452 chr10 59697192 N chr10 59697319 N DUP 5
SRR1766471.280476 chr3 21058621 N chr3 21058680 N DEL 7
SRR1766482.8309198 chr3 21058617 N chr3 21058680 N DEL 7
SRR1766479.10335913 chr3 21058612 N chr3 21058687 N DEL 7
SRR1766466.338198 chr3 21058613 N chr3 21058692 N DEL 3
SRR1766483.10833624 chr10 54332394 N chr10 54332467 N DEL 1
SRR1766462.3264366 chr10 54332394 N chr10 54332467 N DEL 4
SRR1766447.1311927 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766449.8249127 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766445.9434634 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766473.2895805 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766475.8405594 chr10 54332415 N chr10 54332481 N DUP 10
SRR1766484.353820 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766473.7372831 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766476.9797489 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766481.589331 chr10 54332395 N chr10 54332497 N DUP 28
SRR1766442.46601613 chr10 54332451 N chr10 54332517 N DUP 28
SRR1766443.5132830 chr10 54332451 N chr10 54332517 N DUP 28
SRR1766452.1402192 chr10 54332451 N chr10 54332517 N DUP 28
SRR1766463.1748149 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766464.6431826 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766465.5629767 chr10 54332447 N chr10 54332518 N DUP 18
SRR1766474.206051 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766477.11894468 chr10 54332415 N chr10 54332481 N DUP 38
SRR1766479.1053038 chr10 54332415 N chr10 54332481 N DUP 38
SRR1766485.3998464 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766451.4784982 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766454.6419540 chr10 54332415 N chr10 54332517 N DUP 24
SRR1766458.7801432 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766461.8011289 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766484.2908288 chr10 54332395 N chr10 54332502 N DUP 13
SRR1766473.10376766 chr10 54332415 N chr10 54332481 N DUP 12
SRR1766484.4795239 chr10 54332415 N chr10 54332517 N DUP 26
SRR1766462.7049217 chr10 54332395 N chr10 54332502 N DUP 17
SRR1766446.5320884 chr10 54332395 N chr10 54332502 N DUP 17
SRR1766476.9049963 chr10 54332415 N chr10 54332517 N DUP 12
SRR1766486.9902244 chr10 54332415 N chr10 54332481 N DUP 17
SRR1766466.5574371 chr10 54332395 N chr10 54332502 N DUP 20
SRR1766457.2433659 chr10 54332415 N chr10 54332517 N DUP 30
SRR1766445.2751006 chr10 54332395 N chr10 54332502 N DUP 10
SRR1766452.2995561 chr10 54332415 N chr10 54332481 N DUP 24
SRR1766456.4088960 chr10 54332415 N chr10 54332517 N DUP 23
SRR1766483.1231495 chr10 54332415 N chr10 54332517 N DUP 24
SRR1766450.9512239 chr10 54332415 N chr10 54332517 N DUP 25
SRR1766451.8621775 chr10 54332430 N chr10 54332508 N DEL 10
SRR1766470.5371781 chr10 54332420 N chr10 54332498 N DEL 10
SRR1766445.5636215 chr10 54332420 N chr10 54332498 N DEL 10
SRR1766456.961921 chr10 54332420 N chr10 54332498 N DEL 10
SRR1766452.10728406 chr10 54332425 N chr10 54332503 N DEL 10
SRR1766466.5574371 chr10 54332425 N chr10 54332503 N DEL 10
SRR1766478.4164181 chr10 54332426 N chr10 54332504 N DEL 9
SRR1766465.2268330 chr10 54332429 N chr10 54332507 N DEL 6
SRR1766465.9718384 chr7 29645319 N chr7 29645463 N DEL 5
SRR1766462.186963 chr7 29645319 N chr7 29645463 N DEL 5
SRR1766483.6686925 chr7 29645317 N chr7 29645463 N DEL 5
SRR1766463.5031867 chr7 29645319 N chr7 29645463 N DEL 5
SRR1766442.40955939 chr7 29645319 N chr7 29645463 N DEL 1
SRR1766442.25663924 chr7 29645319 N chr7 29645463 N DEL 5
SRR1766484.12079103 chr7 29645360 N chr7 29645468 N DEL 9
SRR1766475.8042433 chr7 29645332 N chr7 29645385 N DUP 6
SRR1766463.5292752 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766442.24575392 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766472.4590897 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766446.1722364 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766483.3084668 chr7 29645400 N chr7 29645498 N DUP 15
SRR1766470.7666158 chr7 29645401 N chr7 29645499 N DUP 15
SRR1766465.9718384 chr7 29645402 N chr7 29645500 N DUP 14
SRR1766453.295021 chr7 29645337 N chr7 29645388 N DEL 9
SRR1766449.3199308 chr7 29645337 N chr7 29645388 N DEL 9
SRR1766451.4509251 chr7 29645400 N chr7 29645496 N DUP 15
SRR1766484.11721869 chr7 29645400 N chr7 29645496 N DUP 15
SRR1766484.8909243 chr7 29645344 N chr7 29645409 N DEL 13
SRR1766465.9498306 chr7 29645344 N chr7 29645395 N DEL 8
SRR1766469.7612154 chr7 29645344 N chr7 29645395 N DEL 8
SRR1766449.1479476 chr7 29645344 N chr7 29645409 N DEL 11
SRR1766457.4701170 chr11 4569528 N chr11 4569590 N DEL 2
SRR1766453.6447787 chr11 4569379 N chr11 4569604 N DUP 5
SRR1766442.33723652 chrX 785313 N chrX 785453 N DUP 6
SRR1766485.3389116 chr6 170114191 N chr6 170114252 N DUP 8
SRR1766484.3072567 chr6 170114198 N chr6 170114301 N DUP 13
SRR1766459.3894899 chr6 170114189 N chr6 170114322 N DUP 12
SRR1766483.4372668 chr6 170114190 N chr6 170114323 N DUP 15
SRR1766459.1646041 chr6 170114229 N chr6 170114318 N DUP 24
SRR1766450.5150588 chr6 170114229 N chr6 170114318 N DUP 24
SRR1766473.1731086 chr6 170114229 N chr6 170114318 N DUP 23
SRR1766451.1404730 chrX 18418906 N chrX 18418979 N DEL 7
SRR1766464.1781835 chrX 18418906 N chrX 18418979 N DEL 8
SRR1766470.308385 chrX 18418846 N chrX 18418967 N DEL 2
SRR1766471.5555623 chr8 110927035 N chr8 110927128 N DUP 5
SRR1766485.11191357 chr15 101764166 N chr15 101764256 N DUP 3
SRR1766442.29793009 chr15 101764166 N chr15 101764256 N DUP 5
SRR1766462.9492241 chr15 101764166 N chr15 101764256 N DUP 5
SRR1766471.1857383 chr15 101764166 N chr15 101764256 N DUP 5
SRR1766452.2540848 chr15 101764225 N chr15 101764315 N DUP 5
SRR1766485.6905061 chr15 101764319 N chr15 101764411 N DEL 1
SRR1766467.4396470 chr15 101764166 N chr15 101764256 N DUP 5
SRR1766472.694450 chr15 101764224 N chr15 101764316 N DEL 5
SRR1766463.5511179 chr15 101764225 N chr15 101764315 N DUP 5
SRR1766447.3049962 chr15 101764166 N chr15 101764256 N DUP 5
SRR1766453.383796 chr15 101764166 N chr15 101764256 N DUP 5
SRR1766464.2163804 chr15 101764225 N chr15 101764315 N DUP 5
SRR1766451.4407656 chr15 101764227 N chr15 101764317 N DUP 5
SRR1766453.1733493 chr15 101764259 N chr15 101764693 N DUP 10
SRR1766455.4302704 chr15 101764319 N chr15 101764411 N DEL 10
SRR1766484.7666525 chr15 101764289 N chr15 101764634 N DEL 5
SRR1766458.1356069 chr15 101764237 N chr15 101764327 N DUP 3
SRR1766486.3609840 chr15 101764239 N chr15 101764329 N DUP 1
SRR1766460.123773 chr15 101764166 N chr15 101764347 N DUP 7
SRR1766483.4307986 chr15 101764279 N chr15 101764525 N DUP 5
SRR1766446.3617331 chr15 101764224 N chr15 101764316 N DEL 5
SRR1766453.10359876 chr15 101764224 N chr15 101764316 N DEL 5
SRR1766463.3417515 chr15 101764166 N chr15 101764347 N DUP 5
SRR1766473.2541099 chr15 101764224 N chr15 101764316 N DEL 5
SRR1766482.12207217 chr15 101764166 N chr15 101764347 N DUP 10
SRR1766446.9569808 chr15 101764226 N chr15 101764318 N DEL 5
SRR1766450.1604757 chr15 101764350 N chr15 101764693 N DUP 5
SRR1766457.7199974 chr15 101764237 N chr15 101764329 N DEL 2
SRR1766450.5800086 chr15 101764350 N chr15 101764693 N DUP 5
SRR1766475.1006834 chr15 101764402 N chr15 101764656 N DEL 5
SRR1766465.10950306 chr15 101764198 N chr15 101764634 N DEL 20
SRR1766480.8022948 chr15 101764220 N chr15 101764403 N DEL 5
SRR1766467.7537170 chr15 101764198 N chr15 101764634 N DEL 10
SRR1766472.4239090 chr15 101764402 N chr15 101764656 N DEL 5
SRR1766465.8653620 chr15 101764402 N chr15 101764656 N DEL 5
SRR1766467.2935707 chr15 101764220 N chr15 101764403 N DEL 5
SRR1766464.2496722 chr15 101764168 N chr15 101764505 N DUP 1
SRR1766458.7596497 chr15 101764168 N chr15 101764505 N DUP 1
SRR1766464.5071485 chr15 101764168 N chr15 101764505 N DUP 5
SRR1766448.9545282 chr15 101764168 N chr15 101764505 N DUP 5
SRR1766442.43907360 chr15 101764168 N chr15 101764505 N DUP 5
SRR1766448.4117458 chr15 101764168 N chr15 101764505 N DUP 5
SRR1766479.8518422 chr15 101764168 N chr15 101764505 N DUP 5
SRR1766483.11961352 chr15 101764445 N chr15 101764697 N DUP 4
SRR1766485.4017270 chr15 101764464 N chr15 101764716 N DUP 5
SRR1766471.4159492 chr15 101764588 N chr15 101764686 N DEL 5
SRR1766478.7284480 chr15 101764329 N chr15 101764486 N DEL 6
SRR1766479.1802390 chr15 101764199 N chr15 101764538 N DEL 3
SRR1766473.2541099 chr15 101764290 N chr15 101764633 N DUP 5
SRR1766463.10515371 chr15 101764434 N chr15 101764686 N DUP 5
SRR1766472.10453392 chr15 101764434 N chr15 101764686 N DUP 6
SRR1766486.10907114 chr22 47020038 N chr22 47020137 N DUP 5
SRR1766449.1790892 chr8 144601302 N chr8 144601493 N DUP 1
SRR1766463.9448856 chr8 144601367 N chr8 144601740 N DUP 5
SRR1766442.42699791 chr8 144601351 N chr8 144601724 N DUP 5
SRR1766448.3253553 chr8 144601422 N chr8 144601499 N DUP 5
SRR1766443.2825560 chr8 144601311 N chr8 144601466 N DEL 1
SRR1766486.4567720 chr8 144601621 N chr8 144601700 N DUP 8
SRR1766446.7613458 chr8 144601465 N chr8 144601646 N DEL 5
SRR1766477.11396242 chr11 70777034 N chr11 70777184 N DUP 6
SRR1766450.8103163 chr2 240812601 N chr2 240812862 N DUP 7
SRR1766454.5114430 chr2 240812796 N chr2 240812892 N DUP 6
SRR1766464.5226294 chr2 240812755 N chr2 240812906 N DUP 5
SRR1766459.2013915 chr2 240812755 N chr2 240812906 N DUP 5
SRR1766447.3045474 chr2 240812918 N chr2 240813065 N DUP 5
SRR1766459.2013915 chr2 240812903 N chr2 240813013 N DUP 1
SRR1766443.5895509 chr2 240813036 N chr2 240813113 N DEL 4
SRR1766477.775968 chr2 240813036 N chr2 240813113 N DEL 5
SRR1766455.7353378 chr2 240812882 N chr2 240813067 N DUP 5
SRR1766455.8309116 chr2 240813036 N chr2 240813168 N DUP 17
SRR1766470.10372775 chr2 240812711 N chr2 240812992 N DEL 3
SRR1766480.6824114 chr2 240813053 N chr2 240813109 N DUP 8
SRR1766462.8782756 chr2 240812862 N chr2 240813161 N DUP 22
SRR1766450.8103163 chr2 240813025 N chr2 240813176 N DUP 17
SRR1766467.426328 chr2 240813034 N chr2 240813185 N DUP 15
SRR1766442.17802355 chr2 240812914 N chr2 240813025 N DEL 15
SRR1766461.9781002 chr2 240813025 N chr2 240813081 N DUP 9
SRR1766445.5308104 chr2 240813034 N chr2 240813109 N DUP 12
SRR1766469.6886259 chr2 240813030 N chr2 240813181 N DUP 27
SRR1766469.4241378 chr2 240813029 N chr2 240813104 N DUP 10
SRR1766444.3285386 chr2 240812821 N chr2 240813123 N DUP 11
SRR1766478.1226564 chr2 240813034 N chr2 240813109 N DUP 12
SRR1766442.23769213 chr2 240813030 N chr2 240813105 N DUP 22
SRR1766442.6040113 chr2 240813025 N chr2 240813100 N DUP 17
SRR1766464.2540435 chr2 240813053 N chr2 240813185 N DUP 22
SRR1766446.4905422 chr2 240812886 N chr2 240813035 N DEL 12
SRR1766451.1171433 chr2 240812840 N chr2 240813030 N DEL 12
SRR1766480.6824114 chr2 240812838 N chr2 240813028 N DEL 7
SRR1766453.903357 chr2 240813025 N chr2 240813100 N DUP 10
SRR1766445.5308104 chr2 240812905 N chr2 240813035 N DEL 5
SRR1766467.3676091 chr2 240813025 N chr2 240813100 N DUP 13
SRR1766457.3026398 chr2 240812980 N chr2 240813092 N DUP 12
SRR1766460.7765759 chr2 240813030 N chr2 240813105 N DUP 21
SRR1766454.9323411 chr2 240813074 N chr2 240813149 N DUP 6
SRR1766470.1657817 chr2 240813049 N chr2 240813181 N DUP 17
SRR1766470.9988440 chr2 240813034 N chr2 240813109 N DUP 11
SRR1766454.8581403 chr2 240813030 N chr2 240813181 N DUP 8
SRR1766455.8309116 chr2 240812766 N chr2 240813048 N DEL 5
SRR1766442.2156248 chr2 240813025 N chr2 240813081 N DUP 6
SRR1766465.11194010 chr2 240813074 N chr2 240813168 N DUP 5
SRR1766474.11298971 chr2 240813074 N chr2 240813168 N DUP 5
SRR1766442.23769213 chr2 240813074 N chr2 240813149 N DUP 5
SRR1766467.4985569 chr2 240813054 N chr2 240813110 N DUP 10
SRR1766485.11826011 chr2 240813090 N chr2 240813165 N DUP 5
SRR1766458.5999729 chr2 240813074 N chr2 240813149 N DUP 5
SRR1766465.11194010 chr2 240813025 N chr2 240813100 N DUP 20
SRR1766451.5293117 chr2 240813025 N chr2 240813100 N DUP 17
SRR1766484.3223190 chr2 240813093 N chr2 240813149 N DUP 5
SRR1766457.7014094 chr2 240812906 N chr2 240813074 N DEL 5
SRR1766478.1226564 chr2 240813030 N chr2 240813105 N DUP 11
SRR1766475.8746701 chr2 240812908 N chr2 240813076 N DEL 5
SRR1766461.1982519 chr2 240812911 N chr2 240813079 N DEL 5
SRR1766479.7479122 chr2 240812898 N chr2 240813085 N DEL 4
SRR1766464.2317221 chr3 100503112 N chr3 100503177 N DUP 6
SRR1766480.4629870 chr6 121497528 N chr6 121497841 N DEL 32
SRR1766484.8618003 chr1 222138535 N chr1 222139069 N DEL 2
SRR1766458.617247 chr1 222138535 N chr1 222139069 N DEL 3
SRR1766462.4666856 chr1 222138535 N chr1 222139069 N DEL 5
SRR1766481.6370041 chr1 222138464 N chr1 222138541 N DUP 8
SRR1766474.4994567 chr1 222138549 N chr1 222138621 N DEL 7
SRR1766442.22887709 chr1 222138535 N chr1 222138607 N DEL 2
SRR1766478.7777456 chr1 222138535 N chr1 222138607 N DEL 2
SRR1766444.3627954 chr1 222138549 N chr1 222138621 N DEL 7
SRR1766465.7924496 chr1 222138549 N chr1 222138621 N DEL 7
SRR1766442.5293301 chr1 222138549 N chr1 222138621 N DEL 7
SRR1766478.10353635 chr1 222138549 N chr1 222138621 N DEL 7
SRR1766460.2170627 chr1 222138535 N chr1 222138607 N DEL 2
SRR1766479.4018808 chr1 222138566 N chr1 222139065 N DEL 2
SRR1766449.71745 chr1 222138566 N chr1 222139065 N DEL 3
SRR1766455.1677590 chr1 222138566 N chr1 222139065 N DEL 3
SRR1766466.4025446 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766479.9068596 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766454.4070858 chr1 222138464 N chr1 222138576 N DUP 12
SRR1766466.2815478 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766465.5134546 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766463.3102088 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766462.3957041 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766442.6740649 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766481.9479786 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766483.10093285 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766463.4946414 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766470.1619055 chr1 222138602 N chr1 222139065 N DEL 4
SRR1766455.738276 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766479.10421235 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766481.403046 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766457.3455908 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766482.6539943 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766466.5935024 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766455.981657 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766452.10344895 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766473.71052 chr1 222138535 N chr1 222138607 N DEL 7
SRR1766475.11536885 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766481.4222045 chr1 222138638 N chr1 222139065 N DEL 3
SRR1766480.726800 chr1 222138464 N chr1 222138648 N DUP 9
SRR1766472.12031612 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766471.10008279 chr1 222138464 N chr1 222138648 N DUP 10
SRR1766474.2819192 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766447.4359764 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766453.807811 chr1 222138480 N chr1 222138594 N DEL 10
SRR1766453.4410555 chr1 222138464 N chr1 222138720 N DUP 10
SRR1766457.7977743 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766481.8367044 chr1 222138594 N chr1 222139091 N DUP 5
SRR1766465.10286575 chr1 222138435 N chr1 222138593 N DEL 5
SRR1766448.7057918 chr1 222138590 N chr1 222139087 N DUP 5
SRR1766442.27964230 chr1 222138418 N chr1 222138592 N DEL 5
SRR1766477.3983293 chr1 222138593 N chr1 222139090 N DUP 5
SRR1766454.2408489 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766454.8490558 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766452.9703927 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766458.3284469 chr1 222138464 N chr1 222138720 N DUP 10
SRR1766449.9621529 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766457.1804210 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766474.8810035 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766453.9186822 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766483.6083413 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766449.246978 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766449.5873486 chr1 222138525 N chr1 222138621 N DEL 5
SRR1766463.7458923 chr1 222138525 N chr1 222138621 N DEL 5
SRR1766473.10501907 chr1 222138525 N chr1 222138621 N DEL 5
SRR1766475.6317486 chr1 222138590 N chr1 222139087 N DUP 5
SRR1766465.3358518 chr1 222138592 N chr1 222139089 N DUP 5
SRR1766450.6346618 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766449.9188503 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766461.7368103 chr1 222138549 N chr1 222138621 N DEL 11
SRR1766455.1427494 chr1 222138591 N chr1 222139088 N DUP 5
SRR1766458.6167105 chr1 222138621 N chr1 222138716 N DUP 17
SRR1766445.1444277 chr1 222138592 N chr1 222139089 N DUP 5
SRR1766472.9671242 chr1 222138593 N chr1 222139090 N DUP 5
SRR1766474.8810035 chr1 222138594 N chr1 222139091 N DUP 5
SRR1766480.3706325 chr1 222138594 N chr1 222139091 N DUP 5
SRR1766470.3907091 chr1 222138704 N chr1 222139093 N DUP 4
SRR1766470.730542 chr1 222138482 N chr1 222138704 N DEL 8
SRR1766464.8883538 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766474.4994567 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766480.3776867 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766460.6920778 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766443.8166889 chr1 222138621 N chr1 222138680 N DUP 17
SRR1766442.14631633 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766448.10707003 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766450.3388448 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766474.4741407 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766449.3131395 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766450.686287 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766466.2815478 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766443.247536 chr1 222138446 N chr1 222138614 N DEL 7
SRR1766456.740891 chr1 222138590 N chr1 222139087 N DUP 5
SRR1766464.4845557 chr1 222138594 N chr1 222139091 N DUP 5
SRR1766470.1619055 chr1 222138594 N chr1 222139091 N DUP 5
SRR1766483.10165478 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766457.7801531 chr1 222138621 N chr1 222138716 N DUP 17
SRR1766463.7371081 chr1 222138621 N chr1 222138716 N DUP 17
SRR1766446.8970471 chr1 222138549 N chr1 222138621 N DEL 12
SRR1766442.27392663 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766450.1538416 chr1 222138464 N chr1 222138720 N DUP 10
SRR1766470.191399 chr1 222138621 N chr1 222138836 N DUP 5
SRR1766455.2840841 chr1 222138681 N chr1 222138874 N DEL 17
SRR1766449.6015105 chr1 222138512 N chr1 222138814 N DEL 2
SRR1766459.10233140 chr1 222138645 N chr1 222138874 N DEL 17
SRR1766468.6207798 chr1 222138645 N chr1 222138874 N DEL 17
SRR1766460.6807251 chr1 222138645 N chr1 222138874 N DEL 17
SRR1766459.10191300 chr1 222138838 N chr1 222139083 N DUP 5
SRR1766472.10590882 chr1 222138551 N chr1 222138839 N DEL 5
SRR1766477.11406760 chr1 222138847 N chr1 222139092 N DUP 5
SRR1766479.12026076 chr1 222138849 N chr1 222139094 N DUP 4
SRR1766462.6454565 chr1 222138874 N chr1 222139083 N DUP 5
SRR1766461.4249118 chr1 222138551 N chr1 222138875 N DEL 5
SRR1766452.2453572 chr1 222138553 N chr1 222138877 N DEL 5
SRR1766467.2168407 chr1 222138883 N chr1 222139092 N DUP 5
SRR1766447.2156986 chr1 222138885 N chr1 222139094 N DUP 4
SRR1766470.1219278 chr1 222138935 N chr1 222138994 N DUP 12
SRR1766467.3963487 chr1 222138935 N chr1 222138994 N DUP 13
SRR1766485.6487619 chr1 222138935 N chr1 222138994 N DUP 13
SRR1766483.10199415 chr1 222138935 N chr1 222138994 N DUP 13
SRR1766461.9707072 chr1 222138910 N chr1 222139083 N DUP 5
SRR1766450.6139146 chr1 222138935 N chr1 222138994 N DUP 16
SRR1766467.8566483 chr1 222138935 N chr1 222138994 N DUP 16
SRR1766458.80854 chr1 222138553 N chr1 222138913 N DEL 5
SRR1766447.3679167 chr1 222138914 N chr1 222139087 N DUP 5
SRR1766464.8669415 chr1 222138942 N chr1 222139039 N DUP 22
SRR1766473.7230085 chr1 222138941 N chr1 222139038 N DUP 5
SRR1766475.7434629 chr1 222138944 N chr1 222139041 N DUP 2
SRR1766442.23570587 chr1 222138942 N chr1 222139039 N DUP 27
SRR1766475.1358042 chr1 222138977 N chr1 222139042 N DEL 23
SRR1766449.5092166 chr1 222138977 N chr1 222139042 N DEL 21
SRR1766481.6370041 chr1 222138977 N chr1 222139042 N DEL 19
SRR1766445.6910106 chr1 222138977 N chr1 222139042 N DEL 17
SRR1766453.6593069 chr1 222138413 N chr1 222139043 N DEL 10
SRR1766474.4741407 chr1 222138421 N chr1 222139053 N DEL 1
SRR1766460.4984969 chr1 222138966 N chr1 222139059 N DEL 6
SRR1766454.7958236 chr1 222138521 N chr1 222139055 N DEL 2
SRR1766473.10501907 chr1 222138521 N chr1 222139055 N DEL 2
SRR1766480.3776867 chr1 222138522 N chr1 222139056 N DEL 1
SRR1766472.6019506 chr19 28081857 N chr19 28082035 N DUP 1
SRR1766447.2504396 chr19 28081800 N chr19 28082049 N DEL 2
SRR1766474.4024607 chr20 59956962 N chr20 59957067 N DEL 13
SRR1766455.5887717 chr20 59956986 N chr20 59957167 N DEL 9
SRR1766479.1340934 chr20 59957091 N chr20 59957188 N DEL 1
SRR1766468.5624000 chr16 73349761 N chr16 73349892 N DEL 14
SRR1766442.26682763 chr16 73349787 N chr16 73349847 N DEL 5
SRR1766449.1820965 chr16 73349791 N chr16 73349847 N DEL 15
SRR1766462.8181061 chr16 73349787 N chr16 73349847 N DEL 40
SRR1766445.8897429 chr6 39845423 N chr6 39845513 N DUP 10
SRR1766451.419444 chr6 39845533 N chr6 39845634 N DUP 1
SRR1766477.9837302 chr7 136568138 N chr7 136568195 N DUP 5
SRR1766452.4992925 chr3 49148215 N chr3 49148378 N DUP 3
SRR1766461.2539640 chr22 21307853 N chr22 21307989 N DEL 10
SRR1766477.9376893 chr22 21307866 N chr22 21308002 N DEL 5
SRR1766446.757484 chr22 21307820 N chr22 21307873 N DUP 5
SRR1766477.8270310 chr7 374228 N chr7 374295 N DEL 9
SRR1766468.3734584 chr7 374231 N chr7 374298 N DEL 9
SRR1766467.11934303 chr18 57195534 N chr18 57195839 N DEL 1
SRR1766442.15321006 chr18 57195534 N chr18 57195839 N DEL 3
SRR1766475.1263481 chr18 57195534 N chr18 57195839 N DEL 5
SRR1766453.4366155 chr18 57195534 N chr18 57195839 N DEL 5
SRR1766468.1314171 chr18 57195534 N chr18 57195839 N DEL 5
SRR1766458.3310857 chr18 57195534 N chr18 57195839 N DEL 5
SRR1766455.3319618 chr18 57195534 N chr18 57195839 N DEL 5
SRR1766445.1227529 chr18 57195550 N chr18 57195851 N DEL 5
SRR1766468.935971 chr18 57195549 N chr18 57195870 N DEL 2
SRR1766472.9881375 chr18 57195549 N chr18 57195870 N DEL 2
SRR1766442.24342718 chr12 47633363 N chr12 47633428 N DEL 4
SRR1766481.9432372 chr12 47633365 N chr12 47633430 N DEL 2
SRR1766449.10040052 chr12 47633552 N chr12 47633701 N DUP 9
SRR1766475.7155758 chr12 47633336 N chr12 47633742 N DUP 2
SRR1766442.44968766 chr12 47633336 N chr12 47633742 N DUP 2
SRR1766442.42867642 chr14 105083462 N chr14 105083610 N DEL 5
SRR1766442.45672787 chr14 105083583 N chr14 105083738 N DEL 4
SRR1766468.6337788 chr16 24833622 N chr16 24833785 N DUP 6
SRR1766442.27489692 chr1 248671490 N chr1 248671644 N DEL 3
SRR1766485.5533042 chr1 248671523 N chr1 248671779 N DEL 3
SRR1766478.773293 chr1 248671513 N chr1 248671565 N DEL 10
SRR1766443.3378031 chr1 248671495 N chr1 248671545 N DUP 11
SRR1766481.5569726 chr1 248671537 N chr1 248671895 N DEL 24
SRR1766479.9642603 chr1 248671478 N chr1 248671528 N DUP 7
SRR1766485.6704924 chr1 248671591 N chr1 248672255 N DEL 5
SRR1766442.25282649 chr1 248671591 N chr1 248671643 N DEL 5
SRR1766460.4100720 chr1 248671597 N chr1 248671649 N DEL 15
SRR1766480.3023694 chr1 248671541 N chr1 248672154 N DEL 20
SRR1766466.4029576 chr1 248671615 N chr1 248671667 N DEL 5
SRR1766444.6626282 chr1 248671550 N chr1 248671600 N DUP 10
SRR1766485.670378 chr1 248671615 N chr1 248671667 N DEL 5
SRR1766461.1873620 chr1 248671591 N chr1 248671643 N DEL 5
SRR1766459.9088911 chr1 248671615 N chr1 248671667 N DEL 5
SRR1766464.1488881 chr1 248671615 N chr1 248671667 N DEL 5
SRR1766471.6123440 chr1 248671565 N chr1 248671666 N DUP 5
SRR1766473.10864160 chr1 248671694 N chr1 248671848 N DEL 9
SRR1766442.26904559 chr1 248671700 N chr1 248671752 N DEL 10
SRR1766444.2414775 chr1 248671617 N chr1 248671667 N DUP 10
SRR1766453.1743087 chr1 248671667 N chr1 248672278 N DUP 5
SRR1766477.1289963 chr1 248671690 N chr1 248672048 N DEL 5
SRR1766470.10764973 chr1 248671698 N chr1 248671750 N DEL 20
SRR1766477.7562770 chr1 248671698 N chr1 248671750 N DEL 20
SRR1766446.9745601 chr1 248671492 N chr1 248671697 N DEL 10
SRR1766444.3160027 chr1 248671700 N chr1 248671854 N DEL 25
SRR1766443.3378031 chr1 248671593 N chr1 248671747 N DEL 5
SRR1766444.2281295 chr1 248671500 N chr1 248671756 N DEL 5
SRR1766467.11232696 chr1 248671514 N chr1 248671770 N DEL 5
SRR1766475.3397961 chr1 248671690 N chr1 248671793 N DEL 15
SRR1766463.1988046 chr1 248671700 N chr1 248671854 N DEL 20
SRR1766442.15003947 chr1 248671676 N chr1 248671830 N DEL 5
SRR1766454.6453669 chr1 248671649 N chr1 248671854 N DEL 18
SRR1766442.46182949 chr1 248671649 N chr1 248671854 N DEL 17
SRR1766463.9172595 chr1 248671611 N chr1 248671867 N DEL 7
SRR1766453.7832241 chr1 248671649 N chr1 248671854 N DEL 16
SRR1766452.9269382 chr1 248671649 N chr1 248671854 N DEL 15
SRR1766479.2531538 chr1 248671518 N chr1 248671876 N DEL 5
SRR1766444.6554448 chr1 248671899 N chr1 248672051 N DUP 5
SRR1766475.3361687 chr1 248671679 N chr1 248671935 N DEL 6
SRR1766467.7817174 chr1 248671598 N chr1 248672109 N DEL 3
SRR1766444.3106193 chr1 248672050 N chr1 248672153 N DEL 5
SRR1766446.7852720 chr1 248672050 N chr1 248672153 N DEL 5
SRR1766471.2280111 chr1 248671502 N chr1 248672013 N DEL 5
SRR1766459.5820952 chr1 248671796 N chr1 248672052 N DEL 5
SRR1766481.11281124 chr1 248671518 N chr1 248672080 N DEL 5
SRR1766486.10368362 chr1 248671508 N chr1 248672121 N DEL 3
SRR1766474.5697147 chr1 248671795 N chr1 248672153 N DEL 5
SRR1766474.6249825 chr1 248671795 N chr1 248672153 N DEL 5
SRR1766458.6008101 chr1 248671795 N chr1 248672153 N DEL 5
SRR1766468.3889302 chr1 248672057 N chr1 248672160 N DEL 5
SRR1766451.9832788 chr1 248671517 N chr1 248672181 N DEL 11
SRR1766444.6626282 chr1 248671514 N chr1 248672229 N DEL 10
SRR1766452.7339732 chr1 248671591 N chr1 248672255 N DEL 5
SRR1766476.1492918 chr14 41808522 N chr14 41808709 N DUP 4
SRR1766451.2882279 chr14 41808513 N chr14 41808572 N DEL 1
SRR1766442.21176099 chr14 41808516 N chr14 41808713 N DEL 1
SRR1766480.1008855 chr10 39178401 N chr10 39178912 N DUP 6
SRR1766455.8088938 chr10 39178401 N chr10 39178912 N DUP 9
SRR1766454.4107566 chr10 39178416 N chr10 39178927 N DEL 9
SRR1766463.4326132 chr10 39178419 N chr10 39178930 N DEL 8
SRR1766474.11526135 chr10 39178420 N chr10 39178931 N DEL 7
SRR1766466.11209878 chr18 49848423 N chr18 49848495 N DEL 5
SRR1766456.724119 chr17 75872137 N chr17 75872435 N DEL 14
SRR1766482.436339 chr17 75871906 N chr17 75872205 N DEL 10
SRR1766479.9599377 chr14 82607343 N chr14 82607404 N DUP 10
SRR1766452.9045460 chr14 82607295 N chr14 82607348 N DEL 17
SRR1766474.7699060 chr3 79771249 N chr3 79771310 N DUP 6
SRR1766470.3626839 chr3 79771313 N chr3 79771366 N DEL 16
SRR1766457.2863696 chr3 79771313 N chr3 79771366 N DEL 16
SRR1766443.4299929 chr3 79771313 N chr3 79771366 N DEL 16
SRR1766442.42521545 chr3 79771313 N chr3 79771366 N DEL 16
SRR1766453.3847903 chr3 79771313 N chr3 79771366 N DEL 23
SRR1766452.10372461 chr3 79771313 N chr3 79771366 N DEL 28
SRR1766476.6189739 chr3 79771313 N chr3 79771366 N DEL 28
SRR1766478.11206097 chr3 79771269 N chr3 79771336 N DEL 2
SRR1766448.3725473 chr3 79771313 N chr3 79771366 N DEL 28
SRR1766480.4567817 chr3 79771313 N chr3 79771366 N DEL 14
SRR1766472.3445736 chr3 79771313 N chr3 79771366 N DEL 13
SRR1766446.9308234 chr3 79771313 N chr3 79771366 N DEL 10
SRR1766447.5268777 chr3 79771313 N chr3 79771366 N DEL 10
SRR1766447.9036611 chr3 79771313 N chr3 79771366 N DEL 10
SRR1766485.2913517 chr3 79771313 N chr3 79771366 N DEL 9
SRR1766465.5551019 chr3 79771314 N chr3 79771367 N DEL 9
SRR1766451.6874420 chr3 79771315 N chr3 79771368 N DEL 9
SRR1766447.10117963 chr3 79771334 N chr3 79771411 N DEL 3
SRR1766471.6029111 chr17 81809364 N chr17 81809421 N DEL 5
SRR1766472.6680002 chr17 81809331 N chr17 81809438 N DUP 7
SRR1766476.7007132 chr20 53657641 N chr20 53657691 N DUP 6
SRR1766457.5345770 chr18 72966204 N chr18 72966284 N DUP 7
SRR1766475.410540 chr14 73372455 N chr14 73372572 N DUP 11
SRR1766458.9505826 chr8 5137582 N chr8 5137638 N DEL 5
SRR1766442.30819934 chr3 185234638 N chr3 185234740 N DEL 1
SRR1766460.3575807 chr3 185234638 N chr3 185234740 N DEL 4
SRR1766470.3394762 chr3 185234638 N chr3 185234740 N DEL 5
SRR1766442.17851214 chr3 185234638 N chr3 185234740 N DEL 5
SRR1766442.23224411 chr3 185234638 N chr3 185234740 N DEL 5
SRR1766468.6695960 chr3 185234638 N chr3 185234740 N DEL 5
SRR1766454.4468928 chr3 185234642 N chr3 185234744 N DEL 10
SRR1766473.1042833 chr3 185234642 N chr3 185234744 N DEL 10
SRR1766477.379369 chr3 185234652 N chr3 185234754 N DEL 1
SRR1766442.13627180 chr3 185234648 N chr3 185234750 N DEL 5
SRR1766466.7910216 chr3 185234644 N chr3 185234746 N DEL 9
SRR1766471.10897347 chr3 185234648 N chr3 185234750 N DEL 5
SRR1766472.11113620 chr3 185234647 N chr3 185234749 N DEL 6
SRR1766483.10297726 chr3 185234650 N chr3 185234752 N DEL 3
SRR1766444.2785896 chr10 47500958 N chr10 47501119 N DEL 5
SRR1766480.7124154 chr10 47500918 N chr10 47501079 N DEL 50
SRR1766467.10174377 chr10 47500983 N chr10 47501144 N DEL 5
SRR1766460.6260554 chr5 113457760 N chr5 113457919 N DEL 1
SRR1766471.6355433 chr5 113457760 N chr5 113457919 N DEL 2
SRR1766463.23793 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766469.2967933 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766482.974488 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766455.1971677 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766442.47014451 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766460.1599166 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766466.126792 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766479.10157233 chr5 113457891 N chr5 113458048 N DUP 10
SRR1766469.7198026 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766443.3450670 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766442.38274130 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766479.11818483 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766449.5028117 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766478.7423482 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766451.10056006 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766472.2650627 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766457.3286361 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766470.10988022 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766462.9825491 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766451.1847370 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766478.2940952 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766443.3135601 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766474.10181054 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766481.9749085 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766460.935189 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766459.9025141 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766460.9731 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766462.3483180 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766451.9921350 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766463.4513314 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766450.3323057 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766483.3648948 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766485.8723972 chr5 113457884 N chr5 113458041 N DUP 5
SRR1766473.3034832 chr5 113457885 N chr5 113458042 N DUP 5
SRR1766484.1771972 chr5 113457886 N chr5 113458043 N DUP 5
SRR1766447.1272301 chr5 113457888 N chr5 113458045 N DUP 5
SRR1766463.6553965 chr5 113457766 N chr5 113457925 N DEL 9
SRR1766450.6993766 chr5 113457883 N chr5 113458042 N DEL 5
SRR1766465.4316727 chrX 129915132 N chrX 129915445 N DUP 15
SRR1766481.8563156 chr22 10852371 N chr22 10852764 N DEL 7
SRR1766466.10124973 chr22 10852371 N chr22 10852764 N DEL 8
SRR1766472.2097136 chr22 10852371 N chr22 10852764 N DEL 9
SRR1766484.9613249 chr22 10852268 N chr22 10852461 N DUP 10
SRR1766445.1142379 chr22 10852268 N chr22 10852461 N DUP 10
SRR1766443.3365446 chr22 10852385 N chr22 10852778 N DEL 1
SRR1766469.43910 chr22 10852301 N chr22 10852494 N DUP 5
SRR1766484.2905409 chr22 10852259 N chr22 10852454 N DEL 1
SRR1766478.8227075 chr22 10852306 N chr22 10852501 N DEL 2
SRR1766450.1225959 chr2 725677 N chr2 725846 N DEL 5
SRR1766483.5282975 chr18 47366969 N chr18 47367088 N DUP 11
SRR1766457.5688609 chr1 1109035 N chr1 1109127 N DUP 10
SRR1766444.3461233 chr1 1109017 N chr1 1109141 N DUP 5
SRR1766442.38086200 chr1 1109035 N chr1 1109127 N DUP 16
SRR1766468.114204 chr1 1109057 N chr1 1109186 N DEL 8
SRR1766467.10013687 chr3 11605270 N chr3 11605449 N DEL 4
SRR1766469.6198993 chr9 41772921 N chr9 41773012 N DEL 5
SRR1766447.2076169 chr9 41772980 N chr9 41773101 N DEL 1
SRR1766485.3660307 chr9 41772872 N chr9 41772993 N DEL 10
SRR1766459.8409490 chr17 82386500 N chr17 82386569 N DUP 15
SRR1766462.9749659 chr17 82386500 N chr17 82386569 N DUP 6
SRR1766465.1688822 chr17 82386500 N chr17 82386569 N DUP 5
SRR1766470.5713670 chr17 82386538 N chr17 82386588 N DUP 9
SRR1766464.4382881 chr17 82386448 N chr17 82386519 N DEL 5
SRR1766465.7696133 chr17 82386453 N chr17 82386524 N DEL 5
SRR1766481.6552074 chr17 82386455 N chr17 82386526 N DEL 3
SRR1766476.8693519 chr17 82386582 N chr17 82386634 N DEL 5
SRR1766486.11731478 chr17 82386582 N chr17 82386634 N DEL 5
SRR1766482.10168135 chr17 82386451 N chr17 82386643 N DEL 5
SRR1766453.2055080 chr17 82386454 N chr17 82386646 N DEL 3
SRR1766475.42300 chr17 82386456 N chr17 82386648 N DEL 1
SRR1766482.4236878 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766443.556153 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766456.549974 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766442.42119236 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766443.2869696 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766442.15663745 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766442.32601120 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766469.6568722 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766461.10319547 chr21 41887630 N chr21 41887772 N DUP 5
SRR1766443.6471730 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766475.376015 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766483.10551491 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766449.3863223 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766460.9515969 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766474.1350636 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766454.10169443 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766484.9455887 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766470.11129279 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766472.2305390 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766479.81902 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766471.12080401 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766467.5426662 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766482.11807608 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766450.6968671 chr21 41887682 N chr21 41887776 N DUP 5
SRR1766484.1162010 chr6 52014664 N chr6 52014805 N DEL 5
SRR1766478.6257576 chr6 52014649 N chr6 52014851 N DEL 9
SRR1766470.1159129 chr6 52014651 N chr6 52014843 N DUP 5
SRR1766476.4971546 chr6 52014651 N chr6 52014843 N DUP 5
SRR1766462.5300438 chr6 52014651 N chr6 52014843 N DUP 5
SRR1766446.10385175 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766450.11060074 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766485.11909878 chr6 52014649 N chr6 52014943 N DEL 9
SRR1766463.8032437 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766472.4152114 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766462.10319172 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766445.8448833 chr6 52014649 N chr6 52014943 N DEL 9
SRR1766460.2284660 chr6 52014649 N chr6 52014943 N DEL 9
SRR1766460.9634889 chr6 52014653 N chr6 52014939 N DEL 13
SRR1766484.6897562 chr6 52014652 N chr6 52014946 N DEL 9
SRR1766478.6257576 chr6 52014655 N chr6 52014949 N DEL 4
SRR1766442.42094979 chr6 52014655 N chr6 52014941 N DEL 13
SRR1766484.11597001 chr6 52014655 N chr6 52014941 N DEL 13
SRR1766442.24946104 chr6 52014656 N chr6 52014950 N DEL 8
SRR1766468.8035034 chr6 52014658 N chr6 52014952 N DEL 6
SRR1766482.7343640 chr6 52014662 N chr6 52014956 N DEL 2
SRR1766466.837833 chr1 22755048 N chr1 22755110 N DUP 13
SRR1766451.4577843 chr1 22754984 N chr1 22755048 N DEL 10
SRR1766457.2714944 chr1 22754986 N chr1 22755050 N DEL 8
SRR1766476.8110657 chr4 180390369 N chr4 180391110 N DEL 3
SRR1766485.2212307 chr4 180390369 N chr4 180391110 N DEL 5
SRR1766484.12077800 chr4 180390369 N chr4 180391110 N DEL 5
SRR1766443.7069877 chr4 180390369 N chr4 180391110 N DEL 5
SRR1766466.6547283 chr4 180390391 N chr4 180390816 N DEL 5
SRR1766447.4244409 chr4 180390391 N chr4 180390816 N DEL 5
SRR1766449.8046268 chr4 180390391 N chr4 180390816 N DEL 5
SRR1766485.7153843 chr4 180390391 N chr4 180390816 N DEL 5
SRR1766479.1726308 chr4 180390392 N chr4 180391140 N DEL 5
SRR1766485.8312066 chr4 180390392 N chr4 180391140 N DEL 5
SRR1766445.463633 chr4 180390392 N chr4 180391140 N DEL 5
SRR1766455.3149196 chr4 180390367 N chr4 180390452 N DEL 2
SRR1766484.9313434 chr4 180390367 N chr4 180390452 N DEL 3
SRR1766444.928956 chr4 180390367 N chr4 180390452 N DEL 6
SRR1766445.1893402 chr4 180390367 N chr4 180390452 N DEL 7
SRR1766471.5261253 chr4 180390409 N chr4 180390936 N DEL 9
SRR1766484.12287193 chr4 180390409 N chr4 180390936 N DEL 11
SRR1766450.194875 chr4 180390409 N chr4 180390936 N DEL 12
SRR1766459.4419610 chr4 180390409 N chr4 180390936 N DEL 13
SRR1766471.7443098 chr4 180390409 N chr4 180390936 N DEL 12
SRR1766460.9806584 chr4 180390409 N chr4 180390936 N DEL 15
SRR1766452.9299665 chr4 180390409 N chr4 180390936 N DEL 15
SRR1766450.10652025 chr4 180390409 N chr4 180390936 N DEL 15
SRR1766479.139386 chr4 180390409 N chr4 180390936 N DEL 15
SRR1766472.3155088 chr4 180390444 N chr4 180390809 N DEL 14
SRR1766462.7069828 chr4 180390417 N chr4 180390886 N DEL 22
SRR1766459.4403780 chr4 180390452 N chr4 180390887 N DEL 19
SRR1766451.438492 chr4 180390414 N chr4 180391137 N DUP 11
SRR1766470.10014425 chr4 180390487 N chr4 180390586 N DEL 7
SRR1766442.17689936 chr4 180390487 N chr4 180390586 N DEL 7
SRR1766459.5624152 chr4 180390380 N chr4 180390533 N DUP 13
SRR1766483.6671724 chr4 180390380 N chr4 180390533 N DUP 13
SRR1766443.6654511 chr4 180390402 N chr4 180390477 N DUP 23
SRR1766478.11533604 chr4 180390374 N chr4 180390531 N DUP 9
SRR1766483.8177189 chr4 180390368 N chr4 180390497 N DUP 9
SRR1766453.944544 chr4 180390470 N chr4 180390925 N DEL 14
SRR1766477.1269157 chr4 180390393 N chr4 180390452 N DEL 10
SRR1766484.11443669 chr4 180390382 N chr4 180390453 N DEL 9
SRR1766442.1455741 chr4 180390383 N chr4 180390454 N DEL 9
SRR1766448.4970352 chr4 180390385 N chr4 180390456 N DEL 9
SRR1766474.7871701 chr4 180390393 N chr4 180390464 N DEL 9
SRR1766463.7852344 chr4 180390554 N chr4 180390971 N DUP 12
SRR1766482.10433225 chr4 180390391 N chr4 180390466 N DEL 7
SRR1766479.5240832 chr4 180390393 N chr4 180390464 N DEL 9
SRR1766443.6654511 chr4 180390428 N chr4 180390575 N DUP 8
SRR1766442.28328481 chr4 180390393 N chr4 180390464 N DEL 9
SRR1766452.7536901 chr4 180390425 N chr4 180390488 N DEL 5
SRR1766453.175560 chr4 180390563 N chr4 180391010 N DEL 17
SRR1766464.5492340 chr4 180390565 N chr4 180391028 N DEL 10
SRR1766463.10119812 chr4 180390380 N chr4 180390577 N DUP 13
SRR1766463.2829584 chr4 180390531 N chr4 180390598 N DEL 19
SRR1766476.542262 chr4 180390413 N chr4 180390488 N DEL 11
SRR1766464.10665890 chr4 180390425 N chr4 180390488 N DEL 10
SRR1766467.2050280 chr4 180390500 N chr4 180390607 N DUP 8
SRR1766447.4650057 chr4 180390505 N chr4 180391050 N DUP 16
SRR1766473.4308230 chr4 180390544 N chr4 180390617 N DUP 14
SRR1766484.7957851 chr4 180390530 N chr4 180391208 N DUP 20
SRR1766485.2214726 chr4 180390474 N chr4 180390550 N DUP 7
SRR1766445.2808920 chr4 180390521 N chr4 180390608 N DEL 12
SRR1766444.2556506 chr4 180390576 N chr4 180390639 N DUP 21
SRR1766442.15525373 chr4 180390582 N chr4 180390651 N DUP 19
SRR1766459.11342664 chr4 180390454 N chr4 180390553 N DUP 9
SRR1766463.10231352 chr4 180390544 N chr4 180390617 N DUP 14
SRR1766445.1266894 chr4 180390416 N chr4 180390585 N DUP 5
SRR1766453.9285961 chr4 180390416 N chr4 180390585 N DUP 5
SRR1766447.7975053 chr4 180390416 N chr4 180390585 N DUP 6
SRR1766442.7375522 chr4 180390474 N chr4 180390550 N DUP 8
SRR1766466.4311964 chr4 180390390 N chr4 180390584 N DUP 9
SRR1766475.9099197 chr4 180390454 N chr4 180390553 N DUP 4
SRR1766465.5096490 chr4 180390522 N chr4 180391031 N DUP 16
SRR1766453.8198161 chr4 180390554 N chr4 180390663 N DUP 16
SRR1766457.3492504 chr4 180390454 N chr4 180390553 N DUP 4
SRR1766447.4244409 chr4 180390522 N chr4 180391031 N DUP 15
SRR1766484.1149727 chr4 180390500 N chr4 180390575 N DUP 5
SRR1766462.7298785 chr4 180390410 N chr4 180390506 N DEL 15
SRR1766443.2526497 chr4 180390585 N chr4 180390654 N DUP 19
SRR1766459.5463201 chr4 180390522 N chr4 180391031 N DUP 13
SRR1766472.6517602 chr4 180390544 N chr4 180390637 N DUP 14
SRR1766463.10231352 chr4 180390401 N chr4 180390500 N DEL 10
SRR1766455.341676 chr4 180390496 N chr4 180390561 N DUP 7
SRR1766462.5206312 chr4 180390532 N chr4 180390597 N DUP 10
SRR1766467.9349849 chr4 180390575 N chr4 180390646 N DUP 17
SRR1766451.8325002 chr4 180390454 N chr4 180390607 N DUP 8
SRR1766467.9349849 chr4 180390557 N chr4 180390658 N DUP 19
SRR1766443.3998687 chr4 180390598 N chr4 180391109 N DUP 11
SRR1766476.10044986 chr4 180390532 N chr4 180390597 N DUP 10
SRR1766448.8151012 chr4 180390627 N chr4 180390816 N DEL 9
SRR1766448.6423808 chr4 180390627 N chr4 180390816 N DEL 10
SRR1766464.2668361 chr4 180390544 N chr4 180390637 N DUP 14
SRR1766456.4045381 chr4 180390530 N chr4 180391208 N DUP 19
SRR1766474.9021775 chr4 180390454 N chr4 180390669 N DUP 15
SRR1766447.8760417 chr4 180390576 N chr4 180391031 N DUP 22
SRR1766470.8122318 chr4 180390376 N chr4 180390626 N DUP 15
SRR1766475.3706410 chr4 180390425 N chr4 180390544 N DEL 10
SRR1766461.6673320 chr4 180390576 N chr4 180390639 N DUP 16
SRR1766469.6715686 chr4 180390428 N chr4 180390627 N DUP 2
SRR1766451.379061 chr4 180390564 N chr4 180391210 N DUP 12
SRR1766484.828261 chr4 180390474 N chr4 180390595 N DUP 16
SRR1766445.2102350 chr4 180390407 N chr4 180390498 N DEL 11
SRR1766466.5507101 chr4 180390510 N chr4 180390839 N DUP 11
SRR1766457.4507058 chr4 180390598 N chr4 180391059 N DUP 18
SRR1766446.30308 chr4 180390401 N chr4 180390534 N DEL 10
SRR1766467.10523921 chr4 180390544 N chr4 180390595 N DUP 14
SRR1766473.8686144 chr4 180390544 N chr4 180390595 N DUP 14
SRR1766453.989434 chr4 180390428 N chr4 180390569 N DEL 10
SRR1766442.37506877 chr4 180390532 N chr4 180390619 N DUP 13
SRR1766466.1386725 chr4 180390548 N chr4 180390805 N DUP 8
SRR1766461.11144720 chr4 180390600 N chr4 180391029 N DUP 15
SRR1766483.1096213 chr4 180390569 N chr4 180391050 N DUP 17
SRR1766452.2302878 chr4 180390575 N chr4 180390646 N DUP 2
SRR1766455.53868 chr4 180390530 N chr4 180390773 N DUP 8
SRR1766483.2267552 chr4 180390575 N chr4 180390646 N DUP 3
SRR1766449.2156050 chr4 180390649 N chr4 180391161 N DEL 2
SRR1766484.8345527 chr4 180390575 N chr4 180390646 N DUP 5
SRR1766458.3466092 chr4 180390500 N chr4 180390563 N DUP 6
SRR1766475.5697602 chr4 180390376 N chr4 180390626 N DUP 16
SRR1766452.2108395 chr4 180390607 N chr4 180391036 N DUP 17
SRR1766475.11510260 chr4 180390546 N chr4 180390649 N DUP 7
SRR1766479.139386 chr4 180390522 N chr4 180390607 N DUP 20
SRR1766453.10347114 chr4 180390668 N chr4 180390807 N DEL 8
SRR1766454.5424402 chr4 180390604 N chr4 180390994 N DEL 18
SRR1766476.8110657 chr4 180390544 N chr4 180390637 N DUP 15
SRR1766445.463633 chr4 180390575 N chr4 180390644 N DUP 18
SRR1766472.1079366 chr4 180390646 N chr4 180390994 N DEL 12
SRR1766458.2769907 chr4 180390544 N chr4 180390627 N DUP 15
SRR1766442.11889975 chr4 180390505 N chr4 180391050 N DUP 16
SRR1766453.53516 chr4 180390638 N chr4 180390745 N DUP 29
SRR1766453.11134061 chr4 180390545 N chr4 180390638 N DUP 20
SRR1766484.11305872 chr4 180390598 N chr4 180390875 N DUP 10
SRR1766458.6553799 chr4 180390538 N chr4 180390646 N DUP 19
SRR1766466.7114130 chr4 180390522 N chr4 180390733 N DUP 14
SRR1766477.4294853 chr4 180390505 N chr4 180390738 N DUP 15
SRR1766461.3163747 chr4 180390538 N chr4 180390646 N DUP 21
SRR1766449.9336359 chr4 180390676 N chr4 180391146 N DEL 22
SRR1766472.3801090 chr4 180390538 N chr4 180390646 N DUP 22
SRR1766471.5533460 chr4 180390538 N chr4 180390646 N DUP 22
SRR1766442.2995494 chr4 180390609 N chr4 180390660 N DEL 18
SRR1766455.6728830 chr4 180390372 N chr4 180390713 N DUP 5
SRR1766463.9271647 chr4 180390454 N chr4 180390541 N DUP 10
SRR1766442.568999 chr4 180390547 N chr4 180390736 N DUP 5
SRR1766481.12960831 chr4 180390549 N chr4 180390738 N DUP 5
SRR1766446.3164411 chr4 180390618 N chr4 180390691 N DUP 14
SRR1766472.8600641 chr4 180390551 N chr4 180391066 N DUP 17
SRR1766460.2011715 chr4 180390393 N chr4 180390650 N DEL 3
SRR1766448.5019961 chr4 180390551 N chr4 180391066 N DUP 17
SRR1766467.10246740 chr4 180390551 N chr4 180391066 N DUP 17
SRR1766455.8286378 chr4 180390640 N chr4 180390735 N DUP 20
SRR1766442.42794430 chr4 180390640 N chr4 180390735 N DUP 20
SRR1766478.1118388 chr4 180390628 N chr4 180390691 N DUP 14
SRR1766477.9996967 chr4 180390554 N chr4 180390745 N DUP 17
SRR1766471.5188130 chr4 180390554 N chr4 180390745 N DUP 14
SRR1766455.7549782 chr4 180390595 N chr4 180390866 N DEL 15
SRR1766481.7475507 chr4 180390893 N chr4 180390979 N DUP 16
SRR1766482.9747182 chr4 180390893 N chr4 180390979 N DUP 16
SRR1766481.6054022 chr4 180390556 N chr4 180391077 N DUP 12
SRR1766476.10967478 chr4 180390556 N chr4 180391077 N DUP 13
SRR1766453.944544 chr4 180390468 N chr4 180391067 N DUP 11
SRR1766466.4819193 chr4 180390680 N chr4 180390943 N DEL 6
SRR1766471.7783539 chr4 180390637 N chr4 180391012 N DEL 25
SRR1766443.6415213 chr4 180390595 N chr4 180391012 N DEL 18
SRR1766476.9582469 chr4 180390628 N chr4 180390691 N DUP 14
SRR1766483.12416279 chr4 180390973 N chr4 180391024 N DUP 16
SRR1766463.8309583 chr4 180390942 N chr4 180391027 N DUP 13
SRR1766463.9279167 chr4 180390935 N chr4 180391050 N DUP 15
SRR1766481.13197869 chr4 180390538 N chr4 180391051 N DUP 15
SRR1766466.1952421 chr4 180390390 N chr4 180390973 N DEL 8
SRR1766470.3960076 chr4 180390546 N chr4 180391109 N DUP 13
SRR1766469.1276665 chr4 180390838 N chr4 180390980 N DEL 12
SRR1766454.532033 chr4 180390562 N chr4 180391095 N DUP 9
SRR1766479.8971394 chr4 180390936 N chr4 180391103 N DUP 11
SRR1766484.6153647 chr4 180390804 N chr4 180390945 N DEL 2
SRR1766451.6369990 chr4 180390804 N chr4 180390995 N DEL 2
SRR1766470.2566927 chr4 180390574 N chr4 180391087 N DUP 9
SRR1766483.1263045 chr4 180390804 N chr4 180390995 N DEL 2
SRR1766442.33295538 chr4 180390988 N chr4 180391087 N DUP 18
SRR1766454.7691693 chr4 180390574 N chr4 180391087 N DUP 10
SRR1766448.9780384 chr4 180390599 N chr4 180391004 N DEL 6
SRR1766453.10166399 chr4 180390599 N chr4 180391004 N DEL 6
SRR1766486.6814917 chr4 180390988 N chr4 180391087 N DUP 15
SRR1766478.2978765 chr4 180390502 N chr4 180391089 N DUP 13
SRR1766468.6005559 chr4 180390981 N chr4 180391068 N DUP 14
SRR1766469.8261919 chr4 180391005 N chr4 180391094 N DUP 17
SRR1766475.6965280 chr4 180391005 N chr4 180391094 N DUP 17
SRR1766484.2489579 chr4 180390685 N chr4 180391169 N DEL 12
SRR1766449.1749899 chr4 180390591 N chr4 180391050 N DUP 21
SRR1766454.6360892 chr4 180390935 N chr4 180391050 N DUP 21
SRR1766478.5627240 chr4 180390553 N chr4 180391181 N DEL 17
SRR1766464.9414523 chr4 180390608 N chr4 180391214 N DEL 28
SRR1766449.1214453 chr4 180391059 N chr4 180391181 N DEL 29
SRR1766442.47067820 chr4 180390615 N chr4 180391224 N DEL 37
SRR1766445.7827924 chr4 180390615 N chr4 180391224 N DEL 42
SRR1766482.5674698 chr4 180390607 N chr4 180391213 N DEL 23
SRR1766454.5424402 chr4 180390615 N chr4 180391224 N DEL 41
SRR1766473.8686144 chr4 180390607 N chr4 180391213 N DEL 23
SRR1766467.1808429 chr4 180390607 N chr4 180391213 N DEL 22
SRR1766454.6324027 chr4 180390615 N chr4 180391224 N DEL 34
SRR1766449.1749899 chr4 180390615 N chr4 180391224 N DEL 34
SRR1766442.26071044 chr4 180390615 N chr4 180391224 N DEL 33
SRR1766460.7594419 chr4 180390607 N chr4 180391213 N DEL 20
SRR1766442.46293936 chr4 180390413 N chr4 180391213 N DEL 10
SRR1766469.2793875 chr4 180390421 N chr4 180391224 N DEL 23
SRR1766458.4247491 chr4 180390421 N chr4 180391224 N DEL 23
SRR1766453.10166399 chr4 180390421 N chr4 180391224 N DEL 23
SRR1766474.4166687 chr4 180390413 N chr4 180391213 N DEL 10
SRR1766442.33369200 chr4 180390413 N chr4 180391213 N DEL 10
SRR1766458.6553799 chr4 180390413 N chr4 180391213 N DEL 10
SRR1766454.3828767 chr4 180390387 N chr4 180391224 N DEL 15
SRR1766450.2182247 chr2 2750311 N chr2 2750440 N DUP 18
SRR1766449.380163 chr2 2750317 N chr2 2750414 N DUP 4
SRR1766443.6652909 chr2 2750288 N chr2 2750417 N DUP 5
SRR1766474.3865549 chr2 2750299 N chr2 2750539 N DUP 6
SRR1766475.5825530 chr2 2750301 N chr2 2750541 N DUP 2
SRR1766464.5719430 chr2 2750301 N chr2 2750541 N DUP 8
SRR1766483.3248156 chr2 2750547 N chr2 2750603 N DEL 15
SRR1766466.9420768 chr2 2750547 N chr2 2750603 N DEL 17
SRR1766453.356498 chr2 2750547 N chr2 2750603 N DEL 17
SRR1766442.22281966 chr2 2750547 N chr2 2750603 N DEL 17
SRR1766472.10192678 chr2 2750547 N chr2 2750603 N DEL 17
SRR1766479.13543375 chr2 2750418 N chr2 2750579 N DUP 8
SRR1766485.4408538 chr11 17545663 N chr11 17545714 N DEL 5
SRR1766442.5946897 chr17 79701261 N chr17 79701317 N DEL 5
SRR1766463.10329068 chr17 79701428 N chr17 79701565 N DEL 19
SRR1766466.5002608 chr17 79701731 N chr17 79701823 N DEL 6
SRR1766474.3026621 chr17 79701355 N chr17 79701823 N DEL 6
SRR1766465.6622716 chr17 79701377 N chr17 79701898 N DEL 10
SRR1766460.8405020 chr17 79701362 N chr17 79701883 N DEL 5
SRR1766454.3506115 chr17 79701363 N chr17 79701884 N DEL 5
SRR1766478.6264161 chr6 162010661 N chr6 162010762 N DEL 28
SRR1766476.7743555 chr6 162010663 N chr6 162010726 N DEL 32
SRR1766461.2921576 chr6 162010639 N chr6 162010715 N DUP 10
SRR1766454.376527 chr6 162010639 N chr6 162010715 N DUP 10
SRR1766479.4048513 chr6 162010690 N chr6 162011085 N DUP 11
SRR1766486.11476199 chr6 162010682 N chr6 162010753 N DUP 7
SRR1766483.5142264 chr6 162010662 N chr6 162010756 N DEL 9
SRR1766448.3475578 chr6 162010638 N chr6 162010721 N DUP 19
SRR1766469.8231917 chr6 162010640 N chr6 162010809 N DUP 23
SRR1766464.10151878 chr6 162010742 N chr6 162010859 N DUP 15
SRR1766472.2579692 chr6 162010726 N chr6 162010863 N DUP 16
SRR1766461.5979337 chr6 162010736 N chr6 162011095 N DUP 11
SRR1766459.2315868 chr6 162010729 N chr6 162010806 N DUP 17
SRR1766458.6783959 chr6 162010730 N chr6 162010929 N DUP 16
SRR1766442.24017496 chr6 162011193 N chr6 162011641 N DUP 17
SRR1766465.7360623 chr6 162011300 N chr6 162011378 N DUP 34
SRR1766469.10602117 chr6 162011300 N chr6 162011378 N DUP 34
SRR1766452.5136227 chr6 162011290 N chr6 162011365 N DUP 23
SRR1766452.15055 chr6 162011200 N chr6 162011285 N DEL 14
SRR1766477.11353208 chr6 162010442 N chr6 162011459 N DUP 9
SRR1766464.9320101 chr6 162011079 N chr6 162011387 N DEL 2
SRR1766442.25714311 chr6 162011471 N chr6 162011656 N DEL 51
SRR1766444.6190508 chr6 162011471 N chr6 162011656 N DEL 51
SRR1766448.4306549 chr6 162011471 N chr6 162011656 N DEL 30
SRR1766463.1801395 chr6 162011471 N chr6 162011656 N DEL 27
SRR1766480.7989608 chr6 162011471 N chr6 162011656 N DEL 27
SRR1766449.9442248 chr6 162011431 N chr6 162011656 N DEL 21
SRR1766480.7891343 chr6 162011205 N chr6 162011663 N DEL 1
SRR1766483.322228 chr6 162010420 N chr6 162011677 N DEL 5
SRR1766462.5368872 chr10 133443894 N chr10 133443957 N DEL 1
SRR1766442.31307446 chr10 133443933 N chr10 133443994 N DUP 5
SRR1766460.10551259 chr10 133443996 N chr10 133444115 N DUP 5
SRR1766473.1548829 chr21 44592070 N chr21 44592428 N DEL 6
SRR1766444.5972280 chr21 44591841 N chr21 44591968 N DEL 4
SRR1766443.10049907 chr21 44592020 N chr21 44592376 N DUP 35
SRR1766471.8305933 chr21 44592020 N chr21 44592376 N DUP 35
SRR1766485.10431269 chr21 44592020 N chr21 44592376 N DUP 25
SRR1766474.3024844 chr21 44591992 N chr21 44592348 N DUP 5
SRR1766449.4765488 chr21 44592020 N chr21 44592376 N DUP 24
SRR1766476.4651601 chr21 44592020 N chr21 44592376 N DUP 10
SRR1766483.8148887 chr21 44592020 N chr21 44592376 N DUP 10
SRR1766472.9101274 chr21 44592020 N chr21 44592376 N DUP 10
SRR1766483.5298277 chr21 44592020 N chr21 44592376 N DUP 10
SRR1766450.985912 chr21 44592023 N chr21 44592379 N DUP 10
SRR1766474.9009850 chr21 44592029 N chr21 44592385 N DUP 5
SRR1766482.6040281 chr21 44592152 N chr21 44592244 N DUP 5
SRR1766470.8655630 chr21 44592152 N chr21 44592244 N DUP 5
SRR1766460.1594864 chr21 44592020 N chr21 44592376 N DUP 3
SRR1766466.6902338 chr21 44592020 N chr21 44592376 N DUP 3
SRR1766471.2235854 chr21 44592020 N chr21 44592376 N DUP 4
SRR1766442.35438280 chr21 44592020 N chr21 44592376 N DUP 30
SRR1766464.9726640 chr10 62370098 N chr10 62370151 N DUP 7
SRR1766454.7696305 chr10 62370207 N chr10 62370322 N DEL 5
SRR1766470.3248882 chr10 62370207 N chr10 62370322 N DEL 7
SRR1766445.7761047 chr10 62370105 N chr10 62370384 N DUP 7
SRR1766463.10410612 chr10 62370207 N chr10 62370322 N DEL 7
SRR1766475.1414942 chr10 62370098 N chr10 62370179 N DUP 7
SRR1766444.6192668 chr10 62370179 N chr10 62370322 N DEL 7
SRR1766480.5960956 chr10 62370207 N chr10 62370322 N DEL 3
SRR1766479.2383398 chr10 62370207 N chr10 62370322 N DEL 6
SRR1766451.3564425 chr10 62370098 N chr10 62370151 N DUP 7
SRR1766479.5282877 chr10 62370207 N chr10 62370322 N DEL 7
SRR1766479.2836380 chr10 62370207 N chr10 62370322 N DEL 7
SRR1766470.2909655 chr10 62370098 N chr10 62370151 N DUP 7
SRR1766451.4145670 chr10 62370207 N chr10 62370322 N DEL 7
SRR1766472.2214094 chr10 62370207 N chr10 62370322 N DEL 7
SRR1766465.9662192 chr10 62370179 N chr10 62370324 N DEL 9
SRR1766470.5109988 chr10 62370179 N chr10 62370324 N DEL 9
SRR1766471.11923041 chr10 62370179 N chr10 62370324 N DEL 9
SRR1766471.1752403 chr10 62370179 N chr10 62370322 N DEL 7
SRR1766458.479807 chr10 62370179 N chr10 62370324 N DEL 9
SRR1766448.5719136 chr10 62370179 N chr10 62370322 N DEL 7
SRR1766443.10118154 chr10 62370179 N chr10 62370324 N DEL 9
SRR1766461.9839282 chr10 62370179 N chr10 62370324 N DEL 9
SRR1766474.4000908 chr10 62370151 N chr10 62370322 N DEL 7
SRR1766457.8636531 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766485.6071582 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766449.7172061 chr10 62370151 N chr10 62370322 N DEL 7
SRR1766485.11791759 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766471.8908687 chr10 62370151 N chr10 62370322 N DEL 7
SRR1766454.4909792 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766466.9069368 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766458.1924551 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766469.10779747 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766458.1924551 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766486.5019417 chr10 62370151 N chr10 62370324 N DEL 9
SRR1766468.1645065 chr10 62370123 N chr10 62370324 N DEL 9
SRR1766478.9624923 chr10 62370123 N chr10 62370322 N DEL 7
SRR1766442.32678365 chr10 62370104 N chr10 62370331 N DEL 6
SRR1766457.9228327 chr10 62370106 N chr10 62370333 N DEL 4
SRR1766473.8103408 chr10 62370442 N chr10 62371227 N DEL 18
SRR1766474.9835975 chr10 62370456 N chr10 62370520 N DEL 14
SRR1766483.1161636 chr10 62370456 N chr10 62370520 N DEL 14
SRR1766442.10435810 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766482.4763274 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766442.44983845 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766472.6901547 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766481.11281261 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766479.5205598 chr10 62370442 N chr10 62370816 N DEL 14
SRR1766458.2540289 chr10 62370492 N chr10 62371252 N DEL 5
SRR1766482.2569140 chr10 62370492 N chr10 62371252 N DEL 5
SRR1766465.1358823 chr10 62370476 N chr10 62370609 N DEL 25
SRR1766444.5133737 chr10 62370456 N chr10 62370578 N DEL 31
SRR1766481.5667546 chr10 62370448 N chr10 62370628 N DEL 33
SRR1766483.2472541 chr10 62370448 N chr10 62370628 N DEL 36
SRR1766468.4425924 chr10 62370487 N chr10 62370602 N DEL 35
SRR1766453.8332201 chr10 62370419 N chr10 62370548 N DUP 4
SRR1766453.437737 chr10 62370419 N chr10 62370548 N DUP 4
SRR1766451.6475581 chr10 62370459 N chr10 62371349 N DUP 13
SRR1766454.5464023 chr10 62370472 N chr10 62370556 N DUP 12
SRR1766472.7780208 chr10 62370472 N chr10 62370556 N DUP 12
SRR1766486.1035245 chr10 62370472 N chr10 62370536 N DUP 4
SRR1766469.9363987 chr10 62370439 N chr10 62370606 N DUP 10
SRR1766472.6668756 chr10 62370509 N chr10 62370575 N DUP 5
SRR1766476.5322532 chr10 62370607 N chr10 62371260 N DUP 31
SRR1766465.9662192 chr10 62370667 N chr10 62371215 N DEL 4
SRR1766461.856574 chr10 62370667 N chr10 62371215 N DEL 5
SRR1766473.2857913 chr10 62370584 N chr10 62371255 N DUP 26
SRR1766468.4165849 chr10 62370628 N chr10 62370685 N DUP 16
SRR1766486.2026388 chr10 62370607 N chr10 62371260 N DUP 18
SRR1766465.9426169 chr10 62370394 N chr10 62370735 N DUP 5
SRR1766446.2021540 chr10 62370773 N chr10 62370824 N DEL 3
SRR1766483.7509108 chr10 62370489 N chr10 62370689 N DEL 14
SRR1766463.2283060 chr10 62370489 N chr10 62370689 N DEL 14
SRR1766450.4901618 chr10 62370489 N chr10 62370689 N DEL 13
SRR1766467.11907405 chr10 62370791 N chr10 62370869 N DEL 11
SRR1766460.6498764 chr10 62370791 N chr10 62370869 N DEL 12
SRR1766449.408250 chr10 62370791 N chr10 62370869 N DEL 12
SRR1766483.3007261 chr10 62370707 N chr10 62370801 N DUP 13
SRR1766446.8689418 chr10 62370707 N chr10 62370801 N DUP 13
SRR1766475.3600823 chr10 62370707 N chr10 62370801 N DUP 13
SRR1766471.9827554 chr10 62370750 N chr10 62370828 N DUP 22
SRR1766475.1761349 chr10 62370750 N chr10 62370828 N DUP 24
SRR1766453.874456 chr10 62370750 N chr10 62370828 N DUP 25
SRR1766477.3191317 chr10 62371045 N chr10 62371435 N DUP 27
SRR1766460.3236897 chr10 62370997 N chr10 62371319 N DUP 14
SRR1766477.7288064 chr10 62370997 N chr10 62371319 N DUP 14
SRR1766478.9704075 chr10 62370998 N chr10 62371320 N DUP 13
SRR1766450.6102635 chr10 62371037 N chr10 62371190 N DUP 25
SRR1766477.3191317 chr10 62371041 N chr10 62371122 N DUP 6
SRR1766483.4505711 chr10 62370439 N chr10 62371077 N DEL 9
SRR1766474.1030344 chr10 62371134 N chr10 62371189 N DUP 17
SRR1766449.9409974 chr10 62371128 N chr10 62371264 N DUP 29
SRR1766466.8289641 chr10 62371128 N chr10 62371264 N DUP 28
SRR1766455.4451455 chr10 62371128 N chr10 62371264 N DUP 25
SRR1766472.10783213 chr10 62371208 N chr10 62371297 N DUP 17
SRR1766442.38681972 chr10 62371208 N chr10 62371297 N DUP 16
SRR1766458.2012467 chr10 62370572 N chr10 62371128 N DEL 17
SRR1766462.11124359 chr10 62371209 N chr10 62371293 N DUP 36
SRR1766464.7645344 chr10 62371128 N chr10 62371264 N DUP 34
SRR1766450.2799415 chr10 62371128 N chr10 62371264 N DUP 33
SRR1766460.3236897 chr10 62371200 N chr10 62371302 N DUP 26
SRR1766460.11272820 chr10 62371209 N chr10 62371293 N DUP 35
SRR1766465.4221373 chr10 62371209 N chr10 62371293 N DUP 35
SRR1766456.1453839 chr10 62370472 N chr10 62371160 N DEL 3
SRR1766460.4981163 chr10 62370544 N chr10 62371226 N DEL 11
SRR1766442.10057080 chr10 62370472 N chr10 62371160 N DEL 3
SRR1766447.2680118 chr10 62370544 N chr10 62371226 N DEL 11
SRR1766459.5340769 chr10 62371035 N chr10 62371289 N DUP 11
SRR1766458.386574 chr10 62371209 N chr10 62371293 N DUP 35
SRR1766447.1331450 chr10 62371209 N chr10 62371293 N DUP 36
SRR1766473.8585888 chr10 62370440 N chr10 62371324 N DUP 4
SRR1766449.9354824 chr10 62370574 N chr10 62371227 N DEL 15
SRR1766474.6230009 chr10 62370641 N chr10 62371350 N DUP 5
SRR1766442.36098140 chr10 62370641 N chr10 62371350 N DUP 8
SRR1766459.5912398 chr10 62370641 N chr10 62371350 N DUP 9
SRR1766474.7089512 chr10 62370641 N chr10 62371350 N DUP 9
SRR1766463.9309583 chr10 62370641 N chr10 62371350 N DUP 10
SRR1766472.1990295 chr10 62370641 N chr10 62371350 N DUP 10
SRR1766442.23639227 chr10 62370661 N chr10 62371350 N DUP 12
SRR1766459.7640060 chr10 62370661 N chr10 62371350 N DUP 13
SRR1766468.7101019 chr10 62370661 N chr10 62371350 N DUP 15
SRR1766447.3273557 chr10 62370661 N chr10 62371350 N DUP 16
SRR1766470.4571153 chr10 62370661 N chr10 62371350 N DUP 18
SRR1766475.6643257 chr10 62370463 N chr10 62371362 N DUP 14
SRR1766442.16091078 chr10 62370463 N chr10 62371362 N DUP 16
SRR1766457.5323815 chr10 62371330 N chr10 62371438 N DUP 4
SRR1766463.2059416 chr10 62370659 N chr10 62371381 N DEL 20
SRR1766472.100128 chr10 62371441 N chr10 62371531 N DUP 17
SRR1766449.1569407 chr10 62371147 N chr10 62371401 N DEL 11
SRR1766472.2210632 chr10 62371147 N chr10 62371401 N DEL 12
SRR1766471.10937371 chr10 62371227 N chr10 62371449 N DUP 27
SRR1766476.10880071 chr10 62371227 N chr10 62371449 N DUP 27
SRR1766481.5366256 chr10 62371419 N chr10 62371509 N DUP 20
SRR1766442.35009943 chr10 62371342 N chr10 62371419 N DEL 17
SRR1766483.8121208 chr10 62370450 N chr10 62371423 N DEL 11
SRR1766450.2799415 chr10 62371362 N chr10 62371499 N DEL 9
SRR1766472.2765911 chr10 62371349 N chr10 62371426 N DEL 8
SRR1766485.6959853 chr10 62371419 N chr10 62371509 N DUP 25
SRR1766468.7101019 chr10 62370711 N chr10 62371431 N DEL 3
SRR1766474.4442024 chr10 62370537 N chr10 62371440 N DEL 9
SRR1766479.844802 chr10 62370538 N chr10 62371441 N DEL 9
SRR1766470.4571153 chr10 62371362 N chr10 62371499 N DEL 14
SRR1766443.3644545 chr10 62371362 N chr10 62371499 N DEL 11
SRR1766474.6714397 chr10 62371343 N chr10 62371453 N DEL 1
SRR1766459.5912398 chr10 62371400 N chr10 62371468 N DEL 9
SRR1766481.1999257 chr10 62370483 N chr10 62371471 N DEL 9
SRR1766472.4502727 chr10 62370389 N chr10 62371471 N DEL 12
SRR1766475.9920196 chr10 62371477 N chr10 62371540 N DUP 6
SRR1766466.186680 chr10 62371362 N chr10 62371499 N DEL 20
SRR1766485.6747037 chr10 62371362 N chr10 62371499 N DEL 19
SRR1766446.2942575 chr10 62371362 N chr10 62371499 N DEL 19
SRR1766473.389348 chr10 62371367 N chr10 62371522 N DEL 21
SRR1766442.35009943 chr10 62371367 N chr10 62371522 N DEL 21
SRR1766460.11272820 chr10 62371367 N chr10 62371522 N DEL 21
SRR1766444.3315944 chr10 62371368 N chr10 62371523 N DEL 21
SRR1766456.5460621 chr10 62370536 N chr10 62371499 N DEL 16
SRR1766446.9787988 chr10 62371365 N chr10 62371520 N DEL 19
SRR1766463.9309583 chr10 62371365 N chr10 62371520 N DEL 19
SRR1766450.8728826 chr10 62371343 N chr10 62371520 N DEL 13
SRR1766447.3718226 chr10 62370457 N chr10 62371521 N DEL 12
SRR1766476.10094059 chr10 62370458 N chr10 62371522 N DEL 12
SRR1766462.6477231 chr10 62370450 N chr10 62371523 N DEL 11
SRR1766457.6641208 chr9 89254409 N chr9 89254828 N DEL 5
SRR1766478.3632890 chr9 89254390 N chr9 89254628 N DUP 16
SRR1766457.924407 chr9 89254362 N chr9 89254418 N DUP 9
SRR1766471.1406341 chr9 89254362 N chr9 89254418 N DUP 10
SRR1766481.7223719 chr9 89254380 N chr9 89254445 N DUP 5
SRR1766470.5150812 chr9 89254378 N chr9 89254665 N DUP 1
SRR1766442.13338086 chr9 89254496 N chr9 89254617 N DEL 20
SRR1766474.1220066 chr9 89254491 N chr9 89254612 N DEL 20
SRR1766447.5453694 chr9 89254527 N chr9 89254761 N DEL 6
SRR1766457.1922693 chr9 89254379 N chr9 89254530 N DUP 8
SRR1766444.525149 chr9 89254425 N chr9 89254483 N DEL 20
SRR1766471.11312798 chr9 89254135 N chr9 89254628 N DUP 12
SRR1766446.1680281 chr9 89254515 N chr9 89254600 N DEL 5
SRR1766477.9737244 chr9 89254418 N chr9 89254660 N DEL 30
SRR1766444.3368329 chr9 89254391 N chr9 89254640 N DEL 12
SRR1766464.8671432 chr9 89254332 N chr9 89254813 N DEL 10
SRR1766443.4524061 chr9 89254382 N chr9 89254847 N DEL 9
SRR1766460.4310361 chr9 89254386 N chr9 89254847 N DEL 5
SRR1766482.2135009 chr9 89254771 N chr9 89254853 N DEL 9
SRR1766473.1880943 chr9 89254771 N chr9 89254877 N DEL 4
SRR1766477.1721813 chr9 89254202 N chr9 89254861 N DEL 3
SRR1766484.11829728 chr9 89254761 N chr9 89254867 N DEL 5
SRR1766442.10966655 chr2 121138920 N chr2 121138977 N DEL 2
SRR1766476.923467 chr2 121138920 N chr2 121138977 N DEL 2
SRR1766472.10934985 chr1 42385988 N chr1 42386039 N DEL 3
SRR1766476.3522553 chr1 42385883 N chr1 42386055 N DEL 5
SRR1766445.2715382 chr3 101891468 N chr3 101891711 N DEL 5
SRR1766468.4967917 chr3 101891496 N chr3 101891710 N DEL 27
SRR1766445.2576012 chr3 101891503 N chr3 101891782 N DUP 1
SRR1766461.1309879 chr3 101891807 N chr3 101891957 N DEL 5
SRR1766459.7433179 chr3 101891807 N chr3 101891957 N DEL 5
SRR1766442.40296750 chr3 101891541 N chr3 101891822 N DEL 5
SRR1766457.5412595 chr3 101891541 N chr3 101891822 N DEL 5
SRR1766486.3460673 chr3 101891541 N chr3 101891822 N DEL 5
SRR1766474.5053015 chr3 101891541 N chr3 101891822 N DEL 5
SRR1766485.10920699 chr3 101891485 N chr3 101891822 N DEL 5
SRR1766447.8131578 chr3 101891485 N chr3 101891822 N DEL 5
SRR1766447.98876 chr3 101891412 N chr3 101891829 N DEL 5
SRR1766468.4967917 chr3 101891569 N chr3 101891836 N DEL 1
SRR1766462.11183524 chr9 86463042 N chr9 86463123 N DUP 2
SRR1766453.10640705 chr9 86463042 N chr9 86463123 N DUP 4
SRR1766473.8416303 chr9 86463042 N chr9 86463123 N DUP 11
SRR1766448.4580055 chr9 86463210 N chr9 86463275 N DEL 6
SRR1766465.543609 chr9 86463063 N chr9 86463130 N DEL 17
SRR1766474.722261 chr9 86463063 N chr9 86463130 N DEL 17
SRR1766442.30482406 chr9 86463063 N chr9 86463130 N DEL 16
SRR1766479.6879434 chr9 86463065 N chr9 86463132 N DEL 11
SRR1766459.9487662 chr9 86463062 N chr9 86463133 N DEL 11
SRR1766463.2603338 chr9 86463065 N chr9 86463171 N DEL 1
SRR1766446.7599462 chr9 86463064 N chr9 86463170 N DEL 2
SRR1766481.9277817 chr9 86463064 N chr9 86463170 N DEL 2
SRR1766460.1377064 chr9 86462997 N chr9 86463175 N DEL 6
SRR1766486.4446054 chr9 86463084 N chr9 86463220 N DEL 7
SRR1766477.11059651 chr9 86463084 N chr9 86463220 N DEL 7
SRR1766476.6189344 chr9 86463084 N chr9 86463220 N DEL 7
SRR1766482.5325297 chr9 86463080 N chr9 86463220 N DEL 7
SRR1766463.5412444 chr9 86463063 N chr9 86463223 N DEL 7
SRR1766481.1412109 chr9 86463226 N chr9 86463290 N DUP 7
SRR1766470.2736025 chrX 42286098 N chrX 42286173 N DUP 4
SRR1766473.11056231 chr3 48839035 N chr3 48839340 N DEL 5
SRR1766471.12164032 chr13 83380655 N chr13 83380712 N DUP 2
SRR1766466.2151266 chr13 83380699 N chr13 83380754 N DEL 3
SRR1766471.4290421 chr13 83380731 N chr13 83380782 N DEL 21
SRR1766463.9696539 chr13 83380731 N chr13 83380782 N DEL 27
SRR1766477.9032097 chr13 83380677 N chr13 83380782 N DEL 11
SRR1766443.1149649 chr13 83380667 N chr13 83380832 N DEL 5
SRR1766481.12524624 chr13 83380656 N chr13 83380865 N DEL 10
SRR1766460.10782732 chr21 41806374 N chr21 41806690 N DEL 11
SRR1766442.4372818 chr21 41806210 N chr21 41806290 N DUP 10
SRR1766482.13240996 chr21 41806383 N chr21 41806454 N DEL 17
SRR1766470.5985547 chr21 41806140 N chr21 41806228 N DEL 5
SRR1766478.5641816 chr21 41805924 N chr21 41806061 N DUP 5
SRR1766481.8927194 chr21 41806151 N chr21 41806327 N DUP 17
SRR1766470.11074115 chr21 41806223 N chr21 41806318 N DUP 1
SRR1766469.9926387 chr21 41806325 N chr21 41806417 N DEL 16
SRR1766473.8889776 chr21 41806489 N chr21 41806547 N DEL 18
SRR1766484.1831171 chr21 41806228 N chr21 41806665 N DUP 27
SRR1766445.566274 chr21 41806307 N chr21 41806426 N DEL 16
SRR1766447.6306350 chr21 41806152 N chr21 41806584 N DUP 7
SRR1766476.3703027 chr21 41806186 N chr21 41806242 N DUP 17
SRR1766476.7958269 chr21 41806210 N chr21 41806546 N DUP 16
SRR1766444.611543 chr21 41806183 N chr21 41806238 N DEL 12
SRR1766484.2166193 chr21 41806323 N chr21 41806639 N DEL 18
SRR1766452.9152131 chr21 41806263 N chr21 41806334 N DUP 14
SRR1766459.2739168 chr21 41805931 N chr21 41806155 N DEL 6
SRR1766445.1901079 chr21 41806288 N chr21 41806362 N DUP 19
SRR1766442.44317868 chr21 41806255 N chr21 41806727 N DUP 12
SRR1766458.7000275 chr21 41806187 N chr21 41806544 N DUP 8
SRR1766479.9912411 chr21 41806230 N chr21 41806837 N DUP 2
SRR1766442.31815950 chr21 41806169 N chr21 41806331 N DUP 14
SRR1766458.7756977 chr21 41806161 N chr21 41806216 N DEL 5
SRR1766474.10598312 chr21 41806169 N chr21 41806239 N DEL 11
SRR1766446.2582196 chr21 41806135 N chr21 41806253 N DEL 10
SRR1766479.4774370 chr21 41806214 N chr21 41806282 N DUP 10
SRR1766470.8640975 chr21 41806195 N chr21 41806585 N DUP 13
SRR1766461.10308705 chr21 41806169 N chr21 41806331 N DUP 14
SRR1766452.1363878 chr21 41806198 N chr21 41806383 N DUP 3
SRR1766473.41245 chr21 41805892 N chr21 41806188 N DEL 5
SRR1766446.8352937 chr21 41806246 N chr21 41806302 N DUP 13
SRR1766474.6163715 chr21 41806182 N chr21 41806343 N DUP 10
SRR1766480.3595308 chr21 41806222 N chr21 41806443 N DEL 16
SRR1766471.6681576 chr21 41806351 N chr21 41806403 N DEL 4
SRR1766456.2850148 chr21 41806381 N chr21 41806437 N DEL 5
SRR1766456.5892728 chr21 41806210 N chr21 41806495 N DUP 10
SRR1766482.360597 chr21 41806361 N chr21 41806541 N DUP 21
SRR1766463.9678769 chr21 41806210 N chr21 41806350 N DUP 12
SRR1766472.1682337 chr21 41806279 N chr21 41806692 N DUP 8
SRR1766447.8793223 chr21 41806275 N chr21 41806636 N DEL 6
SRR1766447.6731503 chr21 41805852 N chr21 41806266 N DUP 1
SRR1766466.9286961 chr21 41806151 N chr21 41806767 N DUP 8
SRR1766462.507819 chr21 41806216 N chr21 41806329 N DUP 13
SRR1766460.5737883 chr21 41806331 N chr21 41806536 N DEL 19
SRR1766451.6119418 chr21 41806207 N chr21 41806323 N DUP 19
SRR1766451.1777787 chr21 41806230 N chr21 41806599 N DUP 20
SRR1766456.1235504 chr21 41806316 N chr21 41806549 N DEL 8
SRR1766453.5408994 chr21 41806302 N chr21 41806454 N DEL 22
SRR1766446.4924919 chr21 41806344 N chr21 41806636 N DEL 4
SRR1766479.4774370 chr21 41806360 N chr21 41806753 N DEL 10
SRR1766472.1682337 chr21 41806284 N chr21 41806482 N DUP 6
SRR1766442.19177731 chr21 41806140 N chr21 41806544 N DEL 12
SRR1766447.2611677 chr21 41806314 N chr21 41806460 N DEL 9
SRR1766448.10061173 chr21 41806141 N chr21 41806383 N DUP 6
SRR1766454.8150005 chr21 41806161 N chr21 41806255 N DEL 5
SRR1766442.35918755 chr21 41806152 N chr21 41806306 N DEL 12
SRR1766462.8138703 chr21 41806138 N chr21 41806558 N DUP 6
SRR1766473.11226221 chr21 41806140 N chr21 41806255 N DEL 4
SRR1766461.6400848 chr21 41806239 N chr21 41806694 N DUP 10
SRR1766442.19970808 chr21 41806165 N chr21 41806403 N DEL 2
SRR1766486.3566662 chr21 41806135 N chr21 41806253 N DEL 12
SRR1766455.5441746 chr21 41806195 N chr21 41806368 N DUP 17
SRR1766454.9188359 chr21 41806337 N chr21 41806417 N DEL 19
SRR1766467.2469423 chr21 41806222 N chr21 41806775 N DUP 15
SRR1766471.7782337 chr21 41806216 N chr21 41806329 N DUP 13
SRR1766462.507819 chr21 41805867 N chr21 41806232 N DEL 6
SRR1766452.5411341 chr21 41806228 N chr21 41806320 N DUP 15
SRR1766467.6093453 chr21 41806462 N chr21 41806581 N DUP 12
SRR1766452.4513262 chr21 41806195 N chr21 41806293 N DUP 14
SRR1766483.6090902 chr21 41806284 N chr21 41806764 N DEL 18
SRR1766447.7925912 chr21 41806198 N chr21 41806683 N DUP 10
SRR1766455.504532 chr21 41806201 N chr21 41806365 N DUP 12
SRR1766484.182936 chr21 41806135 N chr21 41806253 N DEL 3
SRR1766449.1067258 chr21 41806161 N chr21 41806228 N DEL 12
SRR1766455.5792477 chr21 41806243 N chr21 41806308 N DUP 10
SRR1766447.2395898 chr21 41806194 N chr21 41806752 N DEL 14
SRR1766467.7745823 chr21 41805975 N chr21 41806350 N DUP 8
SRR1766472.1854614 chr21 41806202 N chr21 41806342 N DUP 8
SRR1766465.3093147 chr21 41805944 N chr21 41806285 N DEL 6
SRR1766442.16985810 chr21 41806333 N chr21 41806521 N DEL 21
SRR1766485.6322990 chr21 41806240 N chr21 41806380 N DUP 12
SRR1766481.4157761 chr21 41806162 N chr21 41806380 N DUP 10
SRR1766449.3083375 chr21 41806168 N chr21 41806317 N DUP 26
SRR1766470.4625374 chr21 41806196 N chr21 41806720 N DUP 10
SRR1766456.3360709 chr21 41806237 N chr21 41806323 N DUP 12
SRR1766462.6370980 chr21 41806181 N chr21 41806303 N DUP 12
SRR1766479.12294387 chr21 41806150 N chr21 41806772 N DUP 13
SRR1766445.5013700 chr21 41806277 N chr21 41806719 N DUP 5
SRR1766474.5784086 chr21 41806254 N chr21 41806448 N DEL 12
SRR1766442.39351101 chr21 41806222 N chr21 41806392 N DUP 11
SRR1766442.3101599 chr21 41806209 N chr21 41806593 N DUP 13
SRR1766473.2361154 chr21 41806195 N chr21 41806329 N DUP 18
SRR1766448.5043384 chr21 41806351 N chr21 41806521 N DEL 17
SRR1766473.9285030 chr21 41806421 N chr21 41806814 N DUP 20
SRR1766470.7485156 chr21 41806248 N chr21 41806316 N DUP 1
SRR1766483.2245272 chr21 41806143 N chr21 41806228 N DEL 16
SRR1766470.7074814 chr21 41806136 N chr21 41806336 N DUP 17
SRR1766464.1708541 chr21 41806363 N chr21 41806446 N DEL 5
SRR1766474.5784086 chr21 41806164 N chr21 41806216 N DEL 5
SRR1766458.4548608 chr21 41806289 N chr21 41806339 N DUP 9
SRR1766465.8040727 chr21 41806341 N chr21 41806454 N DEL 20
SRR1766442.12570152 chr21 41806241 N chr21 41806757 N DEL 13
SRR1766464.5726126 chr21 41806291 N chr21 41806683 N DUP 13
SRR1766457.6040645 chr21 41806136 N chr21 41806282 N DUP 7
SRR1766457.9369004 chr21 41806490 N chr21 41806564 N DUP 17
SRR1766460.650262 chr21 41806213 N chr21 41806719 N DUP 13
SRR1766447.1323725 chr21 41806182 N chr21 41806343 N DUP 13
SRR1766463.7942114 chr21 41806145 N chr21 41806222 N DUP 6
SRR1766481.13029015 chr21 41805943 N chr21 41806263 N DEL 6
SRR1766465.922917 chr21 41806282 N chr21 41806637 N DEL 8
SRR1766448.9185457 chr21 41806198 N chr21 41806359 N DUP 14
SRR1766442.43917223 chr21 41806306 N chr21 41806829 N DUP 16
SRR1766466.6208572 chr21 41806155 N chr21 41806235 N DUP 12
SRR1766454.8334503 chr21 41806246 N chr21 41806634 N DEL 11
SRR1766469.7286902 chr21 41806159 N chr21 41806227 N DUP 12
SRR1766478.3901595 chr21 41806265 N chr21 41806517 N DUP 7
SRR1766443.3255838 chr21 41806418 N chr21 41806769 N DUP 11
SRR1766473.11579232 chr21 41806182 N chr21 41806667 N DUP 10
SRR1766459.2526939 chr21 41806258 N chr21 41806323 N DUP 12
SRR1766451.1701559 chr21 41806144 N chr21 41806338 N DUP 4
SRR1766470.8640975 chr21 41806220 N chr21 41806693 N DUP 18
SRR1766450.1600464 chr21 41806218 N chr21 41806288 N DEL 20
SRR1766452.10527393 chr21 41806140 N chr21 41806544 N DEL 12
SRR1766442.44763926 chr21 41806246 N chr21 41806561 N DUP 10
SRR1766442.21669087 chr21 41806147 N chr21 41806477 N DUP 8
SRR1766467.6563996 chr21 41806396 N chr21 41806753 N DEL 23
SRR1766451.1906347 chr21 41806354 N chr21 41806524 N DEL 13
SRR1766449.5210184 chr21 41806182 N chr21 41806283 N DUP 16
SRR1766458.1991 chr21 41806138 N chr21 41806383 N DUP 8
SRR1766463.8505495 chr21 41806186 N chr21 41806305 N DUP 10
SRR1766466.8986444 chr21 41806379 N chr21 41806644 N DEL 13
SRR1766442.4372818 chr21 41806234 N chr21 41806659 N DUP 6
SRR1766444.580946 chr1 77870717 N chr1 77870794 N DEL 5
SRR1766474.706275 chr1 207617649 N chr1 207617708 N DUP 2
SRR1766469.1186929 chr21 41689406 N chr21 41689463 N DEL 5
SRR1766468.1457788 chr21 41689406 N chr21 41689463 N DEL 5
SRR1766478.4338504 chr21 41689406 N chr21 41689463 N DEL 6
SRR1766474.9304335 chr21 41689406 N chr21 41689463 N DEL 6
SRR1766454.7733584 chr21 41689406 N chr21 41689463 N DEL 12
SRR1766447.4972719 chr21 41689406 N chr21 41689463 N DEL 17
SRR1766473.11526555 chr21 41689406 N chr21 41689463 N DEL 23
SRR1766448.2749749 chr21 41689413 N chr21 41689470 N DEL 30
SRR1766454.7733584 chr21 41689406 N chr21 41689463 N DEL 30
SRR1766485.3656635 chr21 41689452 N chr21 41689507 N DUP 1
SRR1766461.2009814 chr21 41689406 N chr21 41689463 N DEL 19
SRR1766474.10444562 chr21 41689406 N chr21 41689463 N DEL 15
SRR1766480.2775272 chr21 41689289 N chr21 41689514 N DEL 4
SRR1766483.12274304 chr21 41689466 N chr21 41689551 N DEL 5
SRR1766473.3761607 chr21 41689444 N chr21 41689585 N DEL 4
SRR1766467.48576 chr21 41689407 N chr21 41689632 N DEL 5
SRR1766463.8545920 chr21 41689372 N chr21 41689653 N DEL 5
SRR1766484.1995272 chr21 41689405 N chr21 41689658 N DEL 5
SRR1766466.3037715 chr21 41689407 N chr21 41689660 N DEL 5
SRR1766455.467584 chr21 41689414 N chr21 41689667 N DEL 1
SRR1766477.8706893 chr1 24799246 N chr1 24799406 N DEL 5
SRR1766445.8144050 chr1 24799301 N chr1 24799659 N DEL 2
SRR1766442.3883391 chr1 24799262 N chr1 24799420 N DUP 5
SRR1766475.1735405 chr1 24799263 N chr1 24799421 N DUP 5
SRR1766443.1630092 chr1 24799591 N chr1 24799672 N DEL 7
SRR1766470.278842 chr1 24799751 N chr1 24799850 N DUP 1
SRR1766460.10388209 chr2 237213142 N chr2 237213318 N DUP 5
SRR1766449.1325271 chr2 237213041 N chr2 237213221 N DUP 1
SRR1766461.668789 chr2 237213041 N chr2 237213221 N DUP 3
SRR1766458.4421562 chr2 237213041 N chr2 237213221 N DUP 5
SRR1766452.6830529 chr2 237213041 N chr2 237213221 N DUP 5
SRR1766455.8405496 chr2 237213041 N chr2 237213221 N DUP 5
SRR1766445.494189 chr2 237213041 N chr2 237213221 N DUP 5
SRR1766459.1391696 chr2 237213041 N chr2 237213221 N DUP 5
SRR1766469.8130379 chr2 237213055 N chr2 237213184 N DEL 5
SRR1766455.3368279 chr2 237213222 N chr2 237213400 N DUP 5
SRR1766451.10269866 chr2 237213089 N chr2 237213271 N DEL 15
SRR1766462.2859043 chr2 237213089 N chr2 237213271 N DEL 10
SRR1766448.3789745 chr2 237213089 N chr2 237213271 N DEL 5
SRR1766442.6969715 chr2 237213099 N chr2 237213281 N DEL 5
SRR1766442.25444463 chr2 237213248 N chr2 237213426 N DUP 5
SRR1766443.9223970 chr2 237213099 N chr2 237213281 N DEL 5
SRR1766476.10129682 chr2 237213119 N chr2 237213255 N DEL 1
SRR1766442.40288973 chr2 237213099 N chr2 237213281 N DEL 5
SRR1766486.6699266 chr2 237213119 N chr2 237213246 N DEL 5
SRR1766450.5588772 chr2 237213089 N chr2 237213271 N DEL 5
SRR1766458.9360887 chr2 237213104 N chr2 237213286 N DEL 5
SRR1766482.8195867 chr2 237213089 N chr2 237213271 N DEL 5
SRR1766442.4228028 chr2 237213089 N chr2 237213271 N DEL 5
SRR1766446.148849 chr2 237213089 N chr2 237213271 N DEL 5
SRR1766442.6774635 chr2 237213089 N chr2 237213271 N DEL 5
SRR1766465.2231821 chr2 237213094 N chr2 237213276 N DEL 5
SRR1766471.1094131 chr2 237213052 N chr2 237213278 N DEL 5
SRR1766464.2769925 chr2 237213101 N chr2 237213283 N DEL 3
SRR1766447.10055837 chr2 237213102 N chr2 237213313 N DEL 5
SRR1766446.5283487 chr2 237213055 N chr2 237213363 N DEL 5
SRR1766483.5364740 chr12 129136984 N chr12 129137040 N DUP 15
SRR1766483.1407132 chr12 129136981 N chr12 129137194 N DUP 5
SRR1766486.5897967 chr12 129136944 N chr12 129137034 N DEL 14
SRR1766466.8294429 chr12 129137128 N chr12 129137346 N DEL 14
SRR1766465.4551593 chr12 129136882 N chr12 129137263 N DEL 1
SRR1766469.8107112 chr12 129136933 N chr12 129137266 N DEL 5
SRR1766462.8529724 chr12 129137305 N chr12 129137373 N DUP 13
SRR1766464.2355358 chr12 129136935 N chr12 129137322 N DEL 4
SRR1766452.7941670 chr12 129136936 N chr12 129137323 N DEL 3
SRR1766446.6281644 chr12 129136789 N chr12 129137346 N DEL 5
SRR1766442.45144305 chr12 129136962 N chr12 129137355 N DEL 1
SRR1766459.9443173 chr9 29018197 N chr9 29018263 N DUP 13
SRR1766484.3136401 chr16 8612801 N chr16 8612914 N DUP 5
SRR1766465.5140907 chr16 8612801 N chr16 8612914 N DUP 5
SRR1766470.9207133 chr16 8612801 N chr16 8612914 N DUP 5
SRR1766480.3249239 chr16 8612801 N chr16 8612914 N DUP 5
SRR1766442.3398025 chr16 8612801 N chr16 8612914 N DUP 5
SRR1766444.6187894 chr16 8612801 N chr16 8612914 N DUP 5
SRR1766442.38550696 chr16 8612801 N chr16 8612914 N DUP 5
SRR1766450.766250 chr16 69478630 N chr16 69478679 N DUP 10
SRR1766446.3775312 chr1 143252731 N chr1 143252807 N DEL 5
SRR1766477.10538957 chr1 143252720 N chr1 143252940 N DUP 5
SRR1766456.1154243 chr1 143252720 N chr1 143252940 N DUP 3
SRR1766474.1805383 chr1 143252720 N chr1 143252940 N DUP 3
SRR1766453.2237855 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766486.4798208 chr1 143252851 N chr1 143252944 N DUP 7
SRR1766449.8723641 chr1 143252837 N chr1 143252956 N DUP 13
SRR1766453.7633560 chr1 143252731 N chr1 143252807 N DEL 5
SRR1766462.7850877 chr1 143252815 N chr1 143252889 N DUP 5
SRR1766485.5199237 chr1 143252720 N chr1 143252940 N DUP 2
SRR1766459.2001175 chr1 143252720 N chr1 143252940 N DUP 2
SRR1766451.2995187 chr1 143252720 N chr1 143252940 N DUP 2
SRR1766473.10371123 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766442.30394635 chr1 143252731 N chr1 143252807 N DEL 5
SRR1766483.6043079 chr1 143252740 N chr1 143252816 N DEL 7
SRR1766447.2681208 chr1 143252720 N chr1 143252940 N DUP 3
SRR1766471.10087879 chr1 143252731 N chr1 143252807 N DEL 5
SRR1766458.5447060 chr1 143252720 N chr1 143252940 N DUP 2
SRR1766476.5538837 chr1 143252720 N chr1 143252940 N DUP 3
SRR1766476.8280623 chr1 143252731 N chr1 143252807 N DEL 5
SRR1766463.4979657 chr1 143252851 N chr1 143252944 N DUP 8
SRR1766450.3976154 chr1 143252720 N chr1 143252940 N DUP 4
SRR1766442.282241 chr1 143252720 N chr1 143252940 N DUP 4
SRR1766463.8544135 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766465.11248058 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766442.29266828 chr1 143252863 N chr1 143252933 N DUP 31
SRR1766459.2069306 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766442.19942282 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766484.754501 chr1 143252720 N chr1 143252940 N DUP 4
SRR1766457.5623702 chr1 143252867 N chr1 143252960 N DUP 4
SRR1766469.2100488 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766442.42165973 chr1 143252732 N chr1 143252808 N DEL 5
SRR1766485.9716711 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766484.10529205 chr1 143252727 N chr1 143252947 N DUP 3
SRR1766466.7102231 chr1 143252720 N chr1 143252940 N DUP 3
SRR1766479.6963010 chr1 143252731 N chr1 143252807 N DEL 5
SRR1766467.9192236 chr1 143252795 N chr1 143252874 N DEL 4
SRR1766473.448722 chr1 143252815 N chr1 143252937 N DUP 3
SRR1766450.2231097 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766479.7061322 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766469.1651792 chr1 143252720 N chr1 143252940 N DUP 5
SRR1766455.1125063 chr1 143252720 N chr1 143252940 N DUP 4
SRR1766443.7275706 chr1 143252732 N chr1 143252808 N DEL 5
SRR1766459.11190465 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766466.478038 chr1 143252748 N chr1 143252876 N DEL 2
SRR1766448.9436169 chr1 143252720 N chr1 143252940 N DUP 3
SRR1766481.276861 chr1 143252720 N chr1 143252940 N DUP 3
SRR1766463.5212223 chr1 143252720 N chr1 143252940 N DUP 1
SRR1766462.4075909 chr1 143252732 N chr1 143252808 N DEL 5
SRR1766465.8273340 chr1 143252732 N chr1 143252808 N DEL 5
SRR1766442.1487754 chr1 143252816 N chr1 143252890 N DUP 2
SRR1766452.10088354 chr1 143252802 N chr1 143252855 N DEL 10
SRR1766469.2803978 chr16 572789 N chr16 572898 N DUP 5
SRR1766454.1677753 chr16 572819 N chr16 572873 N DUP 2
SRR1766462.7977576 chr16 572742 N chr16 572853 N DEL 6
SRR1766467.10876389 chr16 572855 N chr16 572964 N DUP 4
SRR1766469.2610054 chr16 572884 N chr16 572993 N DUP 5
SRR1766486.11107469 chr16 572745 N chr16 572911 N DEL 5
SRR1766471.5903303 chr1 48227376 N chr1 48227776 N DEL 2
SRR1766482.7535552 chr1 48227437 N chr1 48227719 N DEL 12
SRR1766468.4008914 chr1 48227352 N chr1 48227748 N DUP 10
SRR1766484.10413642 chr1 48227352 N chr1 48227748 N DUP 10
SRR1766458.7365467 chr1 48227439 N chr1 48227670 N DEL 12
SRR1766477.7245553 chr1 48227324 N chr1 48227433 N DEL 6
SRR1766473.4958510 chr1 48227385 N chr1 48227451 N DEL 6
SRR1766452.7903858 chr1 48227371 N chr1 48227592 N DUP 9
SRR1766469.2729490 chr1 48227371 N chr1 48227592 N DUP 9
SRR1766478.3658996 chr1 48227431 N chr1 48227544 N DEL 3
SRR1766442.27452924 chr1 48227439 N chr1 48227603 N DEL 14
SRR1766472.9722936 chr1 48227439 N chr1 48227603 N DEL 11
SRR1766481.7906636 chr1 48227439 N chr1 48227603 N DEL 9
SRR1766457.8538438 chr1 48227452 N chr1 48227616 N DEL 10
SRR1766472.1687981 chr1 48227480 N chr1 48227642 N DEL 1
SRR1766447.5758758 chr1 48227442 N chr1 48227606 N DEL 7
SRR1766442.15365569 chr1 48227324 N chr1 48227718 N DUP 5
SRR1766479.5882255 chr1 48227324 N chr1 48227663 N DEL 5
SRR1766453.40431 chr9 43348023 N chr9 43348194 N DEL 4
SRR1766462.5102165 chr9 43348011 N chr9 43348108 N DUP 5
SRR1766463.6850786 chr9 43347921 N chr9 43348023 N DEL 8
SRR1766458.4516773 chr9 43348090 N chr9 43348259 N DUP 10
SRR1766445.1553709 chr13 64512251 N chr13 64512319 N DEL 5
SRR1766474.10559403 chr13 64512251 N chr13 64512319 N DEL 5
SRR1766466.3206846 chr13 64512251 N chr13 64512319 N DEL 5
SRR1766481.220567 chr13 64512251 N chr13 64512319 N DEL 5
SRR1766442.19884481 chr13 64512251 N chr13 64512319 N DEL 5
SRR1766475.1633431 chr13 64512251 N chr13 64512319 N DEL 9
SRR1766449.5439652 chr13 64512251 N chr13 64512319 N DEL 10
SRR1766474.9958923 chr13 64512282 N chr13 64512348 N DUP 5
SRR1766477.5727403 chr13 64512282 N chr13 64512348 N DUP 5
SRR1766452.6196879 chr13 64512282 N chr13 64512348 N DUP 10
SRR1766445.10110973 chr13 64512282 N chr13 64512348 N DUP 6
SRR1766442.7701048 chr13 64512282 N chr13 64512348 N DUP 5
SRR1766456.5544593 chr13 64512282 N chr13 64512348 N DUP 5
SRR1766467.3054642 chr13 64512282 N chr13 64512348 N DUP 5
SRR1766453.8458317 chr13 64512282 N chr13 64512348 N DUP 5
SRR1766473.9068340 chr5 43031885 N chr5 43032301 N DEL 7
SRR1766442.26892609 chr5 43032002 N chr5 43032408 N DEL 8
SRR1766451.4218689 chr5 43032104 N chr5 43032319 N DEL 3
SRR1766459.10711430 chr5 43032211 N chr5 43032270 N DEL 8
SRR1766450.1640922 chr5 43031960 N chr5 43032079 N DEL 14
SRR1766479.2922720 chr5 43032078 N chr5 43032199 N DUP 30
SRR1766448.7722582 chr5 43032027 N chr5 43032211 N DUP 30
SRR1766463.9215058 chr5 43032090 N chr5 43032148 N DEL 27
SRR1766450.10915952 chr5 43032027 N chr5 43032211 N DUP 31
SRR1766469.6876778 chr5 43032027 N chr5 43032211 N DUP 31
SRR1766453.1629404 chr5 43032027 N chr5 43032211 N DUP 33
SRR1766483.7341588 chr5 43032027 N chr5 43032211 N DUP 33
SRR1766485.10285801 chr5 43032261 N chr5 43032366 N DEL 9
SRR1766445.2880406 chr5 43031941 N chr5 43032262 N DUP 10
SRR1766485.9416488 chr5 43032123 N chr5 43032195 N DEL 19
SRR1766473.4245758 chr5 43031941 N chr5 43032262 N DUP 15
SRR1766448.2870126 chr5 43031941 N chr5 43032262 N DUP 16
SRR1766473.9068340 chr5 43031941 N chr5 43032262 N DUP 16
SRR1766478.10334282 chr5 43032078 N chr5 43032199 N DUP 19
SRR1766446.8876971 chr5 43032189 N chr5 43032295 N DUP 27
SRR1766448.10120210 chr5 43032181 N chr5 43032262 N DUP 21
SRR1766486.8988579 chr5 43032181 N chr5 43032262 N DUP 18
SRR1766453.6605225 chr5 43032181 N chr5 43032262 N DUP 18
SRR1766449.6650428 chr5 43032189 N chr5 43032295 N DUP 24
SRR1766461.8829494 chr5 43032189 N chr5 43032295 N DUP 29
SRR1766475.7592665 chr5 43032181 N chr5 43032262 N DUP 23
SRR1766481.6751386 chr5 43032078 N chr5 43032199 N DUP 16
SRR1766443.9126058 chr5 43031968 N chr5 43032194 N DEL 8
SRR1766479.8454088 chr5 43032407 N chr5 43032458 N DEL 29
SRR1766473.7931566 chr5 43032407 N chr5 43032458 N DEL 31
SRR1766476.5470935 chr5 43032407 N chr5 43032458 N DEL 31
SRR1766448.3464580 chr5 43032166 N chr5 43032447 N DUP 24
SRR1766476.3704795 chr5 43032125 N chr5 43032414 N DUP 29
SRR1766442.4235579 chr5 43031926 N chr5 43032389 N DEL 10
SRR1766457.3913274 chr5 43031900 N chr5 43032391 N DEL 10
SRR1766448.4974782 chr5 43031902 N chr5 43032393 N DEL 9
SRR1766453.3669188 chr5 43032367 N chr5 43032450 N DEL 32
SRR1766479.11598357 chr5 43032462 N chr5 43032526 N DUP 35
SRR1766474.191719 chr5 43032462 N chr5 43032526 N DUP 29
SRR1766480.978193 chr5 43032180 N chr5 43032449 N DEL 5
SRR1766450.1640922 chr5 43032367 N chr5 43032450 N DEL 16
SRR1766446.8876971 chr5 43032454 N chr5 43032516 N DUP 11
SRR1766463.5462795 chr22 18369679 N chr22 18370310 N DEL 1
SRR1766443.4607614 chr22 18369679 N chr22 18370310 N DEL 15
SRR1766460.5151530 chr22 18369691 N chr22 18370007 N DEL 5
SRR1766469.8144003 chr22 18369869 N chr22 18370500 N DEL 1
SRR1766455.383445 chr22 18369907 N chr22 18370223 N DEL 2
SRR1766471.6793136 chr22 18369593 N chr22 18369907 N DUP 5
SRR1766469.10435273 chr22 18369593 N chr22 18369907 N DUP 5
SRR1766461.315178 chr22 18369686 N chr22 18370002 N DEL 5
SRR1766455.6097918 chr22 18369686 N chr22 18370002 N DEL 5
SRR1766465.1647216 chr22 18369686 N chr22 18370002 N DEL 5
SRR1766445.3232673 chr22 18369739 N chr22 18370368 N DUP 5
SRR1766455.2608701 chr22 18369749 N chr22 18370378 N DUP 5
SRR1766461.2692580 chr22 18369734 N chr22 18370363 N DUP 5
SRR1766453.6845333 chr22 18369763 N chr22 18370392 N DUP 13
SRR1766477.10486013 chr22 18369763 N chr22 18370392 N DUP 15
SRR1766486.1986731 chr22 18369768 N chr22 18370397 N DUP 8
SRR1766480.4704091 chr22 18369829 N chr22 18370460 N DEL 10
SRR1766465.5453104 chr22 18369773 N chr22 18370402 N DUP 5
SRR1766485.11657075 chr22 18369907 N chr22 18370223 N DEL 5
SRR1766476.2307356 chr22 18369907 N chr22 18370223 N DEL 5
SRR1766460.5151530 chr22 18369907 N chr22 18370223 N DEL 5
SRR1766453.6845333 chr22 18369908 N chr22 18370224 N DEL 5
SRR1766480.4550064 chr22 18369807 N chr22 18370227 N DEL 5
SRR1766455.3697294 chr22 18369735 N chr22 18370364 N DUP 5
SRR1766455.3697294 chr22 18369679 N chr22 18370310 N DEL 5
SRR1766478.6593647 chr22 18369679 N chr22 18370310 N DEL 5
SRR1766480.4550064 chr22 18369679 N chr22 18370310 N DEL 5
SRR1766476.3471834 chr22 18369763 N chr22 18370392 N DUP 10
SRR1766454.430473 chr22 18369829 N chr22 18370460 N DEL 10
SRR1766485.2670937 chr22 18369829 N chr22 18370460 N DEL 5
SRR1766462.8216893 chr22 18369829 N chr22 18370460 N DEL 5
SRR1766460.6710395 chr22 10527116 N chr22 10527206 N DUP 5
SRR1766480.8142036 chr18 57510089 N chr18 57510405 N DEL 4
SRR1766450.9031329 chr18 57510089 N chr18 57510405 N DEL 5
SRR1766457.5978257 chr18 57510089 N chr18 57510405 N DEL 5
SRR1766464.9424044 chr18 57510089 N chr18 57510405 N DEL 5
SRR1766474.10590673 chr18 57510089 N chr18 57510405 N DEL 5
SRR1766457.4185471 chr18 57510089 N chr18 57510405 N DEL 6
SRR1766459.2612625 chr18 57510089 N chr18 57510405 N DEL 8
SRR1766451.10079258 chr18 57510089 N chr18 57510405 N DEL 11
SRR1766457.3096592 chr18 57510089 N chr18 57510405 N DEL 11
SRR1766470.3025904 chr18 57510089 N chr18 57510405 N DEL 15
SRR1766449.10607714 chr18 57510107 N chr18 57510423 N DEL 19
SRR1766454.10361147 chr18 57510089 N chr18 57510405 N DEL 25
SRR1766482.3349832 chr18 57510089 N chr18 57510405 N DEL 25
SRR1766442.27638210 chr18 57510089 N chr18 57510405 N DEL 25
SRR1766449.8983745 chr18 57510089 N chr18 57510405 N DEL 25
SRR1766450.646054 chr18 57510102 N chr18 57510418 N DEL 29
SRR1766467.5930255 chr18 57510089 N chr18 57510405 N DEL 30
SRR1766485.3130853 chr18 57510089 N chr18 57510405 N DEL 31
SRR1766455.4905559 chr18 57510089 N chr18 57510405 N DEL 38
SRR1766456.1169560 chr18 57510168 N chr18 57510482 N DUP 5
SRR1766467.1129899 chr18 57510309 N chr18 57510940 N DEL 6
SRR1766481.6960857 chr18 57510313 N chr18 57510944 N DEL 10
SRR1766451.2995563 chr18 57510338 N chr18 57510969 N DEL 5
SRR1766486.7595106 chr18 57510101 N chr18 57510417 N DEL 3
SRR1766466.6177915 chr18 57510102 N chr18 57510418 N DEL 2
SRR1766484.11364550 chr18 57510099 N chr18 57510415 N DEL 5
SRR1766465.7042304 chr18 57510352 N chr18 57510978 N DUP 1
SRR1766457.4582137 chr18 57510359 N chr18 57510991 N DEL 4
SRR1766482.3349832 chr18 57510363 N chr18 57510993 N DEL 1
SRR1766476.4927544 chr4 1828658 N chr4 1829142 N DEL 5
SRR1766459.2202818 chr4 1828666 N chr4 1828920 N DEL 10
SRR1766484.12098173 chr4 1828538 N chr4 1828668 N DUP 5
SRR1766480.1877353 chr4 1828648 N chr4 1828701 N DEL 17
SRR1766442.21132551 chr4 1828648 N chr4 1828701 N DEL 27
SRR1766481.2319602 chr4 1828664 N chr4 1829379 N DUP 5
SRR1766458.6712066 chr4 1828648 N chr4 1828701 N DEL 14
SRR1766460.6051148 chr4 1828648 N chr4 1828701 N DEL 12
SRR1766442.16185263 chr4 1828701 N chr4 1828827 N DUP 5
SRR1766461.5491812 chr4 1828661 N chr4 1828714 N DEL 2
SRR1766458.2454561 chr4 1828797 N chr4 1829281 N DEL 1
SRR1766454.8781160 chr4 1828632 N chr4 1828938 N DUP 1
SRR1766448.6661967 chr4 1828623 N chr4 1828929 N DUP 2
SRR1766467.7997487 chr4 1828859 N chr4 1829570 N DUP 5
SRR1766462.4568999 chr4 1828928 N chr4 1828978 N DUP 5
SRR1766460.10397151 chr4 1828931 N chr4 1829110 N DEL 7
SRR1766451.4217898 chr4 1828688 N chr4 1828991 N DUP 2
SRR1766459.2202818 chr4 1828705 N chr4 1828959 N DEL 5
SRR1766485.8645800 chr4 1828524 N chr4 1829008 N DUP 5
SRR1766467.11156364 chr4 1828524 N chr4 1829008 N DUP 5
SRR1766486.6919240 chr4 1828704 N chr4 1829009 N DEL 5
SRR1766453.2825784 chr4 1828531 N chr4 1829015 N DUP 5
SRR1766483.9636836 chr4 1828677 N chr4 1829031 N DEL 1
SRR1766475.10731124 chr4 1828930 N chr4 1829107 N DUP 6
SRR1766454.9614146 chr4 1829140 N chr4 1829371 N DEL 7
SRR1766453.1783894 chr4 1829142 N chr4 1829322 N DEL 7
SRR1766476.2999925 chr4 1828653 N chr4 1829187 N DUP 6
SRR1766463.2272550 chr4 1829190 N chr4 1829371 N DEL 5
SRR1766442.33257968 chr4 1828888 N chr4 1829243 N DUP 1
SRR1766461.5491812 chr4 1828667 N chr4 1829153 N DEL 5
SRR1766485.6098567 chr4 1828701 N chr4 1829133 N DEL 5
SRR1766442.1045601 chr4 1828532 N chr4 1829194 N DUP 5
SRR1766465.6480444 chr4 1828950 N chr4 1829181 N DEL 1
SRR1766461.7761117 chr4 1828804 N chr4 1829288 N DEL 5
SRR1766466.8776810 chr4 1828560 N chr4 1829224 N DEL 5
SRR1766453.6536708 chr4 1828557 N chr4 1829221 N DEL 5
SRR1766486.4873356 chr4 1828797 N chr4 1829281 N DEL 5
SRR1766457.7982100 chr4 1828929 N chr4 1829337 N DUP 5
SRR1766471.2680304 chr4 1828555 N chr4 1829219 N DEL 5
SRR1766442.11419759 chr4 1828648 N chr4 1828701 N DEL 21
SRR1766486.3832765 chr4 1828668 N chr4 1829332 N DEL 5
SRR1766460.9155440 chr4 1828903 N chr4 1829260 N DEL 1
SRR1766467.722773 chr4 1828668 N chr4 1829332 N DEL 5
SRR1766467.3652921 chr4 1828920 N chr4 1829377 N DUP 10
SRR1766461.1243451 chr4 1828664 N chr4 1829327 N DEL 2
SRR1766461.1243451 chr4 1828778 N chr4 1829403 N DUP 2
SRR1766467.735690 chr4 1828778 N chr4 1829403 N DUP 1
SRR1766479.6866267 chr4 1828665 N chr4 1829332 N DEL 8
SRR1766469.3650260 chr4 1828656 N chr4 1829323 N DEL 8
SRR1766468.1874683 chr4 1828706 N chr4 1829369 N DEL 5
SRR1766459.4695374 chr4 1829371 N chr4 1829497 N DUP 1
SRR1766480.8195504 chr4 1828536 N chr4 1829505 N DUP 1
SRR1766450.970903 chr4 1828797 N chr4 1829461 N DEL 5
SRR1766447.159061 chr4 1828797 N chr4 1829461 N DEL 5
SRR1766463.898930 chr4 1828887 N chr4 1829424 N DEL 5
SRR1766475.2742768 chr4 1828933 N chr4 1829470 N DEL 15
SRR1766452.8452279 chr4 1828662 N chr4 1829505 N DEL 3
SRR1766468.159034 chr17 2562384 N chr17 2562452 N DEL 9
SRR1766458.7233194 chr10 102666912 N chr10 102667518 N DEL 3
SRR1766482.3246480 chr10 102667080 N chr10 102667689 N DEL 3
SRR1766452.9664530 chr15 27313378 N chr15 27313443 N DUP 10
SRR1766447.6576208 chr15 27313377 N chr15 27313428 N DUP 10
SRR1766446.5127551 chr2 126174285 N chr2 126174422 N DUP 5
SRR1766482.5136050 chr18 7984721 N chr18 7984823 N DUP 10
SRR1766480.442097 chr4 186877495 N chr4 186877686 N DUP 6
SRR1766442.14612109 chr4 186877516 N chr4 186877639 N DUP 7
SRR1766478.7078048 chr4 186877478 N chr4 186877631 N DUP 1
SRR1766442.10058503 chr4 186877598 N chr4 186877675 N DUP 7
SRR1766448.4526397 chr4 186877484 N chr4 186877673 N DEL 7
SRR1766480.1229681 chr4 186877606 N chr4 186877683 N DEL 2
SRR1766461.8065008 chr4 186877620 N chr4 186877701 N DEL 6
SRR1766444.6241753 chr4 186877437 N chr4 186877702 N DEL 5
SRR1766449.3861167 chr1 189818374 N chr1 189818441 N DEL 14
SRR1766455.6062088 chr1 189818374 N chr1 189818441 N DEL 15
SRR1766470.4180350 chr1 189818446 N chr1 189818640 N DEL 5
SRR1766458.2954119 chr1 189818463 N chr1 189818544 N DEL 6
SRR1766467.7146889 chr1 189818463 N chr1 189818544 N DEL 7
SRR1766467.2018974 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766447.90772 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766471.5742663 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766467.1640808 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766442.22141324 chr1 189818463 N chr1 189818544 N DEL 30
SRR1766478.11147337 chr1 189818463 N chr1 189818544 N DEL 32
SRR1766480.7377951 chr1 189818463 N chr1 189818544 N DEL 34
SRR1766442.23091358 chr1 189818463 N chr1 189818544 N DEL 34
SRR1766447.8843032 chr1 189818463 N chr1 189818544 N DEL 26
SRR1766457.7087631 chr1 189818463 N chr1 189818544 N DEL 19
SRR1766479.12461066 chr1 189818463 N chr1 189818544 N DEL 21
SRR1766481.905479 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766459.8411973 chr1 189818463 N chr1 189818544 N DEL 25
SRR1766474.10036292 chr1 189818463 N chr1 189818544 N DEL 28
SRR1766478.7644474 chr1 189818463 N chr1 189818544 N DEL 21
SRR1766469.7515319 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766445.2964457 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766485.5643203 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766451.8874075 chr1 189818463 N chr1 189818544 N DEL 15
SRR1766472.626444 chr1 189818465 N chr1 189818546 N DEL 13
SRR1766454.10039188 chr1 189818466 N chr1 189818547 N DEL 12
SRR1766449.6554457 chr1 189818429 N chr1 189818558 N DEL 1
SRR1766465.538163 chr1 189818429 N chr1 189818558 N DEL 1
SRR1766442.18893423 chr1 189818469 N chr1 189818550 N DEL 9
SRR1766451.6842173 chr1 189818470 N chr1 189818551 N DEL 8
SRR1766442.35552044 chr1 189818615 N chr1 189818692 N DUP 11
SRR1766447.10476117 chr1 189818615 N chr1 189818692 N DUP 13
SRR1766485.12049722 chr1 189818615 N chr1 189818692 N DUP 12
SRR1766461.5924183 chr1 21948030 N chr1 21948328 N DEL 4
SRR1766442.6565731 chr1 21948030 N chr1 21948328 N DEL 4
SRR1766485.2867948 chr1 21948038 N chr1 21948336 N DEL 1
SRR1766445.6597786 chr7 156439887 N chr7 156440150 N DEL 5
SRR1766474.10239983 chr7 156439896 N chr7 156440016 N DEL 5
SRR1766480.8204062 chr7 156439896 N chr7 156440016 N DEL 5
SRR1766486.3526512 chr7 156439918 N chr7 156440012 N DUP 8
SRR1766470.4120270 chr7 156439918 N chr7 156440012 N DUP 13
SRR1766455.9511091 chr7 156439918 N chr7 156440012 N DUP 14
SRR1766481.8055877 chr7 156439917 N chr7 156440178 N DUP 5
SRR1766484.11084322 chr7 156439918 N chr7 156440012 N DUP 16
SRR1766476.10166012 chr7 156439918 N chr7 156440012 N DUP 20
SRR1766481.12119077 chr3 48815846 N chr3 48816168 N DEL 2
SRR1766481.7938549 chr11 2560313 N chr11 2560587 N DEL 5
SRR1766455.9482432 chr8 27254786 N chr8 27254942 N DUP 5
SRR1766483.10038501 chr8 27254786 N chr8 27254942 N DUP 5
SRR1766482.8715084 chr8 27254756 N chr8 27255062 N DEL 1
SRR1766475.7520862 chr15 101763980 N chr15 101764167 N DUP 10
SRR1766485.9640921 chr15 101763983 N chr15 101764443 N DUP 5
SRR1766447.4329449 chr15 101764000 N chr15 101764525 N DUP 5
SRR1766473.9934520 chr15 101764018 N chr15 101764205 N DUP 5
SRR1766481.3494210 chr15 101764107 N chr15 101764290 N DEL 1
SRR1766463.5511179 chr15 101764114 N chr15 101764297 N DEL 5
SRR1766454.4975838 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766470.9548903 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766449.8203485 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766448.6129095 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766468.208823 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766486.3609840 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766486.8349419 chr15 101764117 N chr15 101764300 N DEL 5
SRR1766481.2264342 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766480.7998917 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766484.10597215 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766474.6860704 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766473.1611871 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766464.3563971 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766479.11169002 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766474.8199494 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766475.7389380 chr15 101764107 N chr15 101764290 N DEL 5
SRR1766485.9065566 chr15 101764133 N chr15 101764225 N DEL 5
SRR1766442.2214770 chr15 101764133 N chr15 101764225 N DEL 5
SRR1766465.602449 chr15 101764023 N chr15 101764207 N DUP 8
SRR1766442.28752490 chr15 101764137 N chr15 101764229 N DEL 4
SRR1766472.10944748 chr15 101764148 N chr15 101764238 N DUP 5
SRR1766466.2781627 chr15 101764134 N chr15 101764224 N DUP 5
SRR1766466.8453153 chr15 101764138 N chr15 101764319 N DUP 5
SRR1766460.6232167 chr15 101764138 N chr15 101764319 N DUP 5
SRR1766471.1357120 chr15 101764188 N chr15 101764278 N DUP 3
SRR1766486.8349419 chr15 101764152 N chr15 101764242 N DUP 1
SRR1766448.5979964 chr15 101763979 N chr15 101764168 N DEL 10
SRR1766485.11191357 chr15 101764138 N chr15 101764228 N DUP 3
SRR1766442.29793009 chr15 101764138 N chr15 101764228 N DUP 5
SRR1766462.9492241 chr15 101764138 N chr15 101764228 N DUP 5
SRR1766471.1857383 chr15 101764138 N chr15 101764228 N DUP 5
SRR1766452.2540848 chr15 101764225 N chr15 101764315 N DUP 5
SRR1766485.6905061 chr15 101764319 N chr15 101764411 N DEL 1
SRR1766467.4396470 chr15 101764138 N chr15 101764228 N DUP 5
SRR1766472.694450 chr15 101764224 N chr15 101764316 N DEL 5
SRR1766463.5511179 chr15 101764133 N chr15 101764225 N DEL 5
SRR1766447.3049962 chr15 101764040 N chr15 101764138 N DEL 5
SRR1766453.383796 chr15 101764040 N chr15 101764138 N DEL 5
SRR1766464.2163804 chr15 101764133 N chr15 101764225 N DEL 5
SRR1766451.4407656 chr15 101764135 N chr15 101764227 N DEL 5
SRR1766453.1733493 chr15 101764233 N chr15 101764323 N DUP 5
SRR1766455.4302704 chr15 101764319 N chr15 101764411 N DEL 10
SRR1766484.7666525 chr15 101764063 N chr15 101764341 N DUP 5
SRR1766458.1356069 chr15 101764237 N chr15 101764327 N DUP 3
SRR1766486.3609840 chr15 101764239 N chr15 101764329 N DUP 1
SRR1766460.123773 chr15 101764013 N chr15 101764114 N DEL 10
SRR1766483.4307986 chr15 101764279 N chr15 101764525 N DUP 5
SRR1766446.3617331 chr15 101764224 N chr15 101764316 N DEL 5
SRR1766453.10359876 chr15 101764224 N chr15 101764316 N DEL 5
SRR1766463.3417515 chr15 101764138 N chr15 101764319 N DUP 5
SRR1766473.2541099 chr15 101764036 N chr15 101764316 N DEL 5
SRR1766482.12207217 chr15 101764138 N chr15 101764319 N DUP 5
SRR1766446.9569808 chr15 101764038 N chr15 101764318 N DEL 5
SRR1766457.7199974 chr15 101764237 N chr15 101764329 N DEL 2
SRR1766465.10950306 chr15 101764342 N chr15 101764434 N DEL 15
SRR1766480.8022948 chr15 101764220 N chr15 101764403 N DEL 5
SRR1766467.7537170 chr15 101764319 N chr15 101764411 N DEL 10
SRR1766467.2935707 chr15 101764220 N chr15 101764403 N DEL 5
SRR1766464.2496722 chr15 101763958 N chr15 101764483 N DUP 1
SRR1766458.7596497 chr15 101763958 N chr15 101764483 N DUP 1
SRR1766464.5071485 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766448.9545282 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766442.43907360 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766448.4117458 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766479.8518422 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766479.10390903 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766478.10097603 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766449.2359167 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766486.10628431 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766450.6192012 chr15 101763958 N chr15 101764483 N DUP 5
SRR1766470.2035597 chr1 248840715 N chr1 248841040 N DEL 3
SRR1766442.2483650 chr1 248840715 N chr1 248841040 N DEL 5
SRR1766443.11101196 chr1 248840715 N chr1 248841040 N DEL 5
SRR1766442.35761985 chr1 248840715 N chr1 248841040 N DEL 5
SRR1766457.3751975 chr1 248840752 N chr1 248841239 N DEL 10
SRR1766453.1492532 chr1 248840759 N chr1 248840814 N DEL 10
SRR1766465.9754141 chr1 248840769 N chr1 248841202 N DEL 8
SRR1766450.2723894 chr1 248840795 N chr1 248841228 N DEL 5
SRR1766475.6392393 chr1 248840795 N chr1 248841228 N DEL 6
SRR1766462.10387820 chr1 248840726 N chr1 248840943 N DEL 5
SRR1766461.1976052 chr1 248840732 N chr1 248840949 N DEL 5
SRR1766442.12432060 chr1 248840732 N chr1 248840949 N DEL 5
SRR1766452.10515502 chr1 248840768 N chr1 248841039 N DEL 10
SRR1766473.8138108 chr1 248840768 N chr1 248840985 N DEL 5
SRR1766452.1060870 chr1 248840883 N chr1 248841100 N DEL 5
SRR1766461.3561336 chr1 248840883 N chr1 248841100 N DEL 5
SRR1766460.8491756 chr1 248840931 N chr1 248841040 N DEL 15
SRR1766484.9724356 chr1 248840775 N chr1 248840884 N DEL 5
SRR1766464.9035570 chr1 248840814 N chr1 248840975 N DUP 5
SRR1766452.4225571 chr1 248841011 N chr1 248841228 N DEL 5
SRR1766469.998295 chr1 248841011 N chr1 248841228 N DEL 5
SRR1766466.762248 chr1 248840951 N chr1 248841220 N DUP 5
SRR1766482.11565735 chr1 248841002 N chr1 248841165 N DEL 5
SRR1766442.33002436 chr1 248841126 N chr1 248841287 N DUP 5
SRR1766442.34935425 chr1 248840715 N chr1 248841200 N DUP 2
SRR1766465.7270031 chr1 248841102 N chr1 248841157 N DEL 20
SRR1766463.4565596 chr1 248840985 N chr1 248841202 N DEL 5
SRR1766457.3751975 chr1 248841158 N chr1 248841211 N DUP 15
SRR1766457.4628727 chr1 248841167 N chr1 248841220 N DUP 5
SRR1766482.11236279 chr1 248840901 N chr1 248841172 N DEL 1
SRR1766450.10772327 chr1 248840746 N chr1 248841179 N DEL 1
SRR1766442.34935425 chr1 248840752 N chr1 248841239 N DEL 5
SRR1766458.1620315 chr1 248840759 N chr1 248841246 N DEL 5
SRR1766450.2723894 chr1 248840763 N chr1 248841250 N DEL 4
SRR1766477.2869149 chr1 248840711 N chr1 248841252 N DEL 2
SRR1766481.1898491 chr7 56327682 N chr7 56327738 N DUP 1
SRR1766452.4869508 chr6 169955233 N chr6 169955283 N DUP 5
SRR1766469.9439705 chr6 169955233 N chr6 169955283 N DUP 5
SRR1766460.11125418 chr22 47379316 N chr22 47379377 N DEL 5
SRR1766470.10843239 chr20 46491826 N chr20 46492391 N DEL 5
SRR1766448.6656103 chr20 46491826 N chr20 46492391 N DEL 10
SRR1766467.1561176 chr20 46491974 N chr20 46492539 N DEL 1
SRR1766477.8241628 chr20 46492013 N chr20 46492578 N DEL 5
SRR1766442.26541021 chr20 46492021 N chr20 46492586 N DEL 5
SRR1766455.747913 chr20 46492079 N chr20 46492642 N DUP 5
SRR1766475.4687221 chr20 46491704 N chr20 46492269 N DEL 14
SRR1766482.5618929 chr20 46491924 N chr20 46492489 N DEL 10
SRR1766475.11413882 chr20 46491924 N chr20 46492489 N DEL 5
SRR1766481.5072789 chr20 46491999 N chr20 46492564 N DEL 5
SRR1766453.3177824 chr20 46492030 N chr20 46492595 N DEL 5
SRR1766467.6785081 chr20 46492078 N chr20 46492643 N DEL 5
SRR1766442.7216186 chr20 46492104 N chr20 46492669 N DEL 7
SRR1766444.1779596 chr9 96026767 N chr9 96027098 N DEL 14
SRR1766464.7057425 chr9 96026835 N chr9 96026914 N DEL 10
SRR1766449.1019267 chr9 96026999 N chr9 96027316 N DEL 6
SRR1766449.9526156 chr9 96026928 N chr9 96027008 N DUP 2
SRR1766467.10855619 chr9 96026858 N chr9 96027096 N DUP 5
SRR1766445.6358528 chr9 96026890 N chr9 96027110 N DUP 5
SRR1766458.5838245 chr2 210735167 N chr2 210735232 N DUP 2
SRR1766446.7607364 chr16 16650860 N chr16 16650921 N DEL 11
SRR1766442.15709929 chr3 128544871 N chr3 128544975 N DEL 5
SRR1766468.6569364 chr3 128544871 N chr3 128544975 N DEL 5
SRR1766484.6587304 chr15 50635476 N chr15 50635823 N DUP 7
SRR1766477.977347 chr15 50635468 N chr15 50635819 N DUP 6
SRR1766458.1908230 chr15 50635468 N chr15 50635823 N DUP 12
SRR1766443.1711033 chr15 50635482 N chr15 50635828 N DEL 1
SRR1766444.3033469 chr15 50635482 N chr15 50635825 N DEL 4
SRR1766484.8673329 chr15 50635482 N chr15 50635825 N DEL 4
SRR1766456.4605365 chr5 3856913 N chr5 3856964 N DEL 19
SRR1766462.1133999 chr5 3856913 N chr5 3856964 N DEL 16
SRR1766450.8934125 chr5 3856917 N chr5 3856968 N DEL 11
SRR1766472.6316736 chr5 3856920 N chr5 3856971 N DEL 8
SRR1766453.6404839 chr5 3856927 N chr5 3856978 N DEL 1
SRR1766445.9705740 chr5 3856915 N chr5 3856966 N DEL 13
SRR1766450.340076 chr5 3856914 N chr5 3856965 N DEL 14
SRR1766463.388858 chr5 3856914 N chr5 3856965 N DEL 14
SRR1766484.1667907 chr5 3856924 N chr5 3856975 N DEL 4
SRR1766478.6729064 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766442.24818813 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766444.830058 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766483.8671875 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766484.7267427 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766457.6216621 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766464.10685902 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766455.187207 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766442.31960770 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766467.1193403 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766452.1531853 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766475.9233158 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766486.4764731 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766442.583488 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766442.9698385 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766483.2992174 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766483.3425034 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766458.3861524 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766462.1353904 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766467.5116494 chr10 49965694 N chr10 49965835 N DUP 5
SRR1766482.6038576 chr10 49965696 N chr10 49965837 N DUP 5
SRR1766449.5841681 chr10 49965698 N chr10 49965839 N DUP 5
SRR1766445.3225489 chr10 49965700 N chr10 49965841 N DUP 5
SRR1766447.7586149 chr10 49965701 N chr10 49965842 N DUP 5
SRR1766455.6781495 chr10 49965701 N chr10 49965842 N DUP 5
SRR1766457.2534974 chr10 49965702 N chr10 49965843 N DUP 5
SRR1766442.34700650 chr10 49965736 N chr10 49966264 N DUP 5
SRR1766484.5640815 chr10 49965668 N chr10 49966225 N DEL 15
SRR1766470.955295 chr10 49965668 N chr10 49966225 N DEL 15
SRR1766442.32425161 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766471.9309014 chr5 10347066 N chr5 10347245 N DEL 8
SRR1766464.2361891 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766451.9536241 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766457.5140021 chr5 10347422 N chr5 10347479 N DUP 10
SRR1766473.4259472 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766479.11554488 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766479.4915557 chr5 10347121 N chr5 10347406 N DEL 14
SRR1766448.10258055 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766467.6717490 chr5 10346474 N chr5 10346553 N DEL 38
SRR1766458.727214 chr5 10347121 N chr5 10347406 N DEL 6
SRR1766455.4745641 chr5 10347459 N chr5 10347518 N DEL 10
SRR1766483.7742663 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766457.2314894 chr5 10346474 N chr5 10346553 N DEL 19
SRR1766479.1479799 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766464.3370284 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766483.2867780 chr5 10346474 N chr5 10346553 N DEL 35
SRR1766476.6734492 chr5 10346474 N chr5 10346553 N DEL 35
SRR1766464.10110253 chr5 10347121 N chr5 10347406 N DEL 5
SRR1766454.598117 chr5 10347096 N chr5 10347406 N DEL 16
SRR1766442.43566049 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766445.6967072 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766446.3883240 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766464.2146313 chr5 10346474 N chr5 10346553 N DEL 5
SRR1766453.8023538 chr5 10347623 N chr5 10347862 N DEL 5
SRR1766486.10573528 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766442.5346800 chr5 10347096 N chr5 10347406 N DEL 16
SRR1766482.799618 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766467.5434496 chr5 10347171 N chr5 10347380 N DEL 1
SRR1766486.5371104 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766473.8229187 chr5 10347064 N chr5 10347243 N DEL 8
SRR1766447.1785407 chr5 10347422 N chr5 10347479 N DUP 20
SRR1766453.2294627 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766465.5349876 chr5 10347066 N chr5 10347220 N DEL 8
SRR1766472.1277807 chr5 10347621 N chr5 10347860 N DEL 5
SRR1766459.2422768 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766442.19653289 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766442.30459796 chr5 10347043 N chr5 10347189 N DUP 8
SRR1766448.4911493 chr5 10347459 N chr5 10347518 N DEL 10
SRR1766456.4259598 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766475.3765078 chr5 10347459 N chr5 10347518 N DEL 10
SRR1766445.7189719 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766462.85102 chr5 10347121 N chr5 10347406 N DEL 14
SRR1766466.2970903 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766466.1535782 chr5 10347096 N chr5 10347406 N DEL 20
SRR1766463.7885807 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766472.603517 chr5 10347422 N chr5 10347479 N DUP 19
SRR1766455.4871127 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766479.10716328 chr5 10346422 N chr5 10346566 N DEL 2
SRR1766483.11577964 chr5 10347249 N chr5 10347403 N DUP 8
SRR1766442.30459796 chr5 10346474 N chr5 10346553 N DEL 24
SRR1766471.467521 chr5 10347117 N chr5 10347398 N DEL 14
SRR1766442.21487073 chr5 10347121 N chr5 10347406 N DEL 7
SRR1766472.3204428 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766445.1973245 chr5 10347064 N chr5 10347218 N DEL 8
SRR1766472.11734428 chr5 10347247 N chr5 10347401 N DUP 8
SRR1766449.4092371 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766447.8697643 chr5 10346618 N chr5 10346705 N DEL 5
SRR1766465.9164408 chr5 10347223 N chr5 10347402 N DUP 8
SRR1766450.5186151 chr5 10347224 N chr5 10347403 N DUP 8
SRR1766444.4825970 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766484.4694579 chr5 10346480 N chr5 10346559 N DEL 9
SRR1766453.3510036 chr5 10347462 N chr5 10347521 N DEL 10
SRR1766442.27003599 chr5 10347422 N chr5 10347479 N DUP 17
SRR1766442.38430846 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766464.6603080 chr5 10347121 N chr5 10347406 N DEL 11
SRR1766473.8755073 chr5 10347040 N chr5 10347696 N DUP 8
SRR1766476.3416377 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766447.1632621 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766461.342319 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766468.8046972 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766442.1088889 chr5 10346474 N chr5 10346553 N DEL 18
SRR1766442.17812002 chr5 10346474 N chr5 10346553 N DEL 38
SRR1766453.3959843 chr5 10346677 N chr5 10346775 N DUP 5
SRR1766460.11113871 chr5 10347171 N chr5 10347380 N DEL 3
SRR1766453.3168261 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766442.4704186 chr5 10347117 N chr5 10347398 N DEL 21
SRR1766465.11248369 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766457.5205264 chr5 10347422 N chr5 10347479 N DUP 21
SRR1766480.5179651 chr5 10347358 N chr5 10347530 N DEL 3
SRR1766477.5139514 chr5 10347355 N chr5 10347527 N DEL 6
SRR1766461.8476723 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766482.7899405 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766470.2521746 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766473.9018190 chr5 10347121 N chr5 10347406 N DEL 12
SRR1766477.974189 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766478.2778857 chr5 10347064 N chr5 10347243 N DEL 8
SRR1766464.6603080 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766465.5949856 chr5 10347353 N chr5 10347525 N DEL 8
SRR1766450.2372217 chr5 10347463 N chr5 10347522 N DEL 10
SRR1766482.7899405 chr5 10347759 N chr5 10347841 N DUP 5
SRR1766460.710752 chr5 10347246 N chr5 10347400 N DUP 8
SRR1766470.10643224 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766478.4509846 chr5 10346474 N chr5 10346553 N DEL 38
SRR1766452.7841382 chr5 10347146 N chr5 10347406 N DEL 3
SRR1766442.21349329 chr5 10347358 N chr5 10347530 N DEL 3
SRR1766461.9073438 chr5 10347066 N chr5 10347245 N DEL 8
SRR1766458.5624463 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766478.3642692 chr5 10347171 N chr5 10347380 N DEL 2
SRR1766474.5649070 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766471.7918391 chr5 10347064 N chr5 10347218 N DEL 8
SRR1766485.11054307 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766443.243909 chr5 10346474 N chr5 10346553 N DEL 22
SRR1766453.8023538 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766460.710752 chr5 10346418 N chr5 10346562 N DEL 6
SRR1766467.6090314 chr5 10347096 N chr5 10347406 N DEL 16
SRR1766483.5677680 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766473.2170372 chr5 10347171 N chr5 10347380 N DEL 2
SRR1766443.9267437 chr5 10347759 N chr5 10347841 N DUP 5
SRR1766466.178559 chr5 10347459 N chr5 10347518 N DEL 10
SRR1766458.2527066 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766451.6670309 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766482.3282579 chr5 10347043 N chr5 10347139 N DUP 8
SRR1766472.9116892 chr5 10347775 N chr5 10347859 N DEL 5
SRR1766470.5490836 chr5 10347459 N chr5 10347518 N DEL 15
SRR1766484.10025845 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766445.4596809 chr5 10347043 N chr5 10347164 N DUP 8
SRR1766482.4696391 chr5 10347043 N chr5 10347114 N DUP 8
SRR1766472.1814641 chr5 10346474 N chr5 10346553 N DEL 38
SRR1766445.4449075 chr5 10347092 N chr5 10347398 N DEL 16
SRR1766450.7122101 chr5 10347096 N chr5 10347406 N DEL 16
SRR1766470.4139289 chr5 10346474 N chr5 10346553 N DEL 23
SRR1766459.6238463 chr17 32227666 N chr17 32227797 N DUP 5
SRR1766473.7110824 chr17 32227782 N chr17 32227895 N DUP 14
SRR1766477.6279492 chr9 67775876 N chr9 67776001 N DUP 1
SRR1766477.1230708 chr9 67775876 N chr9 67776001 N DUP 1
SRR1766450.478917 chr9 67775876 N chr9 67776001 N DUP 5
SRR1766472.11606917 chr9 67775876 N chr9 67776001 N DUP 5
SRR1766446.7270238 chr9 67775876 N chr9 67776001 N DUP 5
SRR1766454.6805590 chr9 67775876 N chr9 67776001 N DUP 5
SRR1766478.546252 chr19 9948187 N chr19 9948492 N DEL 33
SRR1766449.4682985 chr19 9948161 N chr19 9948469 N DUP 1
SRR1766480.1543367 chr19 9948256 N chr19 9948561 N DEL 2
SRR1766442.10653256 chr19 9948472 N chr19 9948781 N DUP 5
SRR1766469.7414847 chr19 9948199 N chr19 9948504 N DEL 5
SRR1766457.321800 chr13 62019547 N chr13 62019606 N DEL 12
SRR1766459.9770674 chr13 62019547 N chr13 62019606 N DEL 25
SRR1766462.9835446 chr13 62019547 N chr13 62019606 N DEL 29
SRR1766482.136209 chr13 62019547 N chr13 62019606 N DEL 63
SRR1766470.214716 chr13 62019547 N chr13 62019606 N DEL 27
SRR1766477.3650423 chr13 62019617 N chr13 62019768 N DUP 4
SRR1766467.9727489 chr13 62019617 N chr13 62019768 N DUP 5
SRR1766475.11454397 chr13 62019579 N chr13 62019780 N DUP 5
SRR1766460.7246157 chr13 62019772 N chr13 62019847 N DUP 13
SRR1766481.10670481 chr13 62019789 N chr13 62019848 N DUP 30
SRR1766456.6025753 chr13 62019789 N chr13 62019848 N DUP 27
SRR1766453.6644475 chr13 62019789 N chr13 62019848 N DUP 27
SRR1766469.7787499 chr13 62019789 N chr13 62019848 N DUP 32
SRR1766462.1645298 chr13 62019593 N chr13 62019773 N DEL 7
SRR1766443.6912908 chr13 62019594 N chr13 62019774 N DEL 6
SRR1766486.4097881 chr13 62019535 N chr13 62019775 N DEL 5
SRR1766465.2160569 chr13 62019537 N chr13 62019777 N DEL 5
SRR1766482.12705189 chr13 62019790 N chr13 62019849 N DUP 11
SRR1766443.7295555 chr13 62019592 N chr13 62019825 N DEL 4
SRR1766449.10422640 chr13 62019830 N chr13 62019962 N DUP 6
SRR1766442.13221786 chr13 62019760 N chr13 62019968 N DUP 6
SRR1766457.5752772 chr14 56355292 N chr14 56355345 N DUP 12
SRR1766442.11096501 chr14 56355314 N chr14 56355425 N DUP 23
SRR1766464.7165385 chr14 56355301 N chr14 56355402 N DUP 15
SRR1766449.830077 chr14 56355301 N chr14 56355402 N DUP 14
SRR1766476.4309794 chr14 56355314 N chr14 56355425 N DUP 24
SRR1766471.6849989 chr14 56355285 N chr14 56355452 N DUP 3
SRR1766484.11336252 chr14 56355398 N chr14 56355459 N DUP 9
SRR1766442.37521161 chr14 56355301 N chr14 56355402 N DUP 15
SRR1766460.10419520 chr14 56355398 N chr14 56355459 N DUP 8
SRR1766466.86738 chr14 56355314 N chr14 56355425 N DUP 23
SRR1766476.7815557 chr14 56355337 N chr14 56355420 N DUP 14
SRR1766473.10082444 chr14 56355337 N chr14 56355420 N DUP 14
SRR1766445.417605 chr14 56355337 N chr14 56355420 N DUP 19
SRR1766452.6695738 chr14 56355377 N chr14 56355452 N DEL 15
SRR1766471.10971266 chr14 56355377 N chr14 56355452 N DEL 15
SRR1766468.5157910 chr14 56355377 N chr14 56355452 N DEL 15
SRR1766442.27903440 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766459.917116 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766459.5558079 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766442.18099783 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766454.123169 chr14 56355349 N chr14 56355452 N DEL 15
SRR1766442.352658 chr14 56355331 N chr14 56355452 N DEL 20
SRR1766443.4673862 chr14 56355331 N chr14 56355452 N DEL 20
SRR1766445.8577450 chr14 56355331 N chr14 56355452 N DEL 20
SRR1766460.9076839 chr14 56355331 N chr14 56355452 N DEL 15
SRR1766476.8144751 chr14 56355331 N chr14 56355452 N DEL 20
SRR1766471.7382822 chr14 56355331 N chr14 56355452 N DEL 19
SRR1766442.12914548 chr14 56355313 N chr14 56355452 N DEL 10
SRR1766452.1701095 chr14 56355313 N chr14 56355452 N DEL 10
SRR1766448.8583577 chr14 56355315 N chr14 56355454 N DEL 10
SRR1766451.3735200 chr14 56355315 N chr14 56355454 N DEL 10
SRR1766442.31185038 chr14 56355316 N chr14 56355455 N DEL 10
SRR1766482.2015970 chr14 56355321 N chr14 56355460 N DEL 7
SRR1766472.4282063 chr14 56355322 N chr14 56355461 N DEL 6
SRR1766474.4751411 chr14 56355322 N chr14 56355461 N DEL 6
SRR1766482.3732972 chr14 98835437 N chr14 98835550 N DUP 5
SRR1766459.6607745 chr3 106073612 N chr3 106074350 N DUP 5
SRR1766476.2687489 chr3 106073619 N chr3 106073744 N DUP 5
SRR1766445.1314203 chr3 106073628 N chr3 106073704 N DUP 5
SRR1766451.3963636 chr3 106073742 N chr3 106074531 N DEL 5
SRR1766467.3548026 chr3 106073764 N chr3 106074551 N DEL 6
SRR1766442.44602383 chr3 106073764 N chr3 106074551 N DEL 6
SRR1766461.7696843 chr3 106073780 N chr3 106073859 N DEL 1
SRR1766459.9413742 chr3 106073982 N chr3 106074332 N DEL 3
SRR1766446.9963828 chr3 106073982 N chr3 106074332 N DEL 4
SRR1766479.11971497 chr3 106073938 N chr3 106074161 N DEL 8
SRR1766468.6235911 chr3 106073607 N chr3 106073951 N DEL 5
SRR1766476.8921933 chr3 106073588 N chr3 106074103 N DUP 4
SRR1766465.4333732 chr3 106073619 N chr3 106073744 N DUP 5
SRR1766451.5126359 chr3 106073785 N chr3 106074008 N DEL 4
SRR1766451.3963636 chr3 106074011 N chr3 106074136 N DUP 5
SRR1766455.7262819 chr3 106073719 N chr3 106074033 N DEL 10
SRR1766442.1456353 chr3 106073914 N chr3 106074135 N DUP 2
SRR1766480.5272381 chr3 106073575 N chr3 106074139 N DUP 5
SRR1766475.7221324 chr3 106074060 N chr3 106074145 N DUP 3
SRR1766442.36162605 chr3 106073935 N chr3 106074156 N DUP 1
SRR1766474.10377386 chr3 106073755 N chr3 106073924 N DEL 5
SRR1766452.10478571 chr3 106073935 N chr3 106074156 N DUP 5
SRR1766442.3069708 chr3 106073938 N chr3 106074161 N DEL 10
SRR1766483.1120548 chr3 106073705 N chr3 106074145 N DEL 5
SRR1766452.326692 chr3 106073938 N chr3 106074161 N DEL 10
SRR1766479.7728884 chr3 106073938 N chr3 106074161 N DEL 9
SRR1766458.5240135 chr3 106073946 N chr3 106074169 N DEL 5
SRR1766447.4931990 chr3 106073986 N chr3 106074209 N DEL 5
SRR1766476.2687489 chr3 106073968 N chr3 106074191 N DEL 5
SRR1766448.8109841 chr3 106073600 N chr3 106074166 N DEL 3
SRR1766465.11224372 chr3 106073605 N chr3 106074171 N DEL 1
SRR1766478.3282651 chr3 106073804 N chr3 106074247 N DUP 3
SRR1766461.1228797 chr3 106073918 N chr3 106074313 N DUP 9
SRR1766469.7962070 chr3 106073690 N chr3 106074400 N DUP 5
SRR1766442.39036989 chr3 106073690 N chr3 106074400 N DUP 6
SRR1766449.6523629 chr3 106073690 N chr3 106074400 N DUP 10
SRR1766448.8153443 chr3 106073691 N chr3 106074401 N DUP 13
SRR1766468.985962 chr3 106074213 N chr3 106074388 N DUP 7
SRR1766470.9190658 chr3 106074213 N chr3 106074388 N DUP 7
SRR1766442.10781912 chr3 106073608 N chr3 106073777 N DEL 2
SRR1766464.7306329 chr3 106073619 N chr3 106073744 N DUP 5
SRR1766480.8411971 chr10 106718940 N chr10 106719007 N DEL 5
SRR1766480.6954657 chr10 106718904 N chr10 106718971 N DEL 15
SRR1766442.13005065 chr10 106718971 N chr10 106719036 N DUP 5
SRR1766476.8356049 chr10 106718971 N chr10 106719036 N DUP 5
SRR1766470.8064401 chr10 106718971 N chr10 106719036 N DUP 5
SRR1766449.74085 chr10 106718971 N chr10 106719036 N DUP 5
SRR1766474.6685559 chr10 106718971 N chr10 106719036 N DUP 5
SRR1766484.10391300 chr10 106718928 N chr10 106718995 N DEL 5
SRR1766446.10390265 chr10 106718905 N chr10 106719038 N DEL 5
SRR1766461.6998018 chr10 106719071 N chr10 106719138 N DEL 5
SRR1766466.8086662 chr10 106718905 N chr10 106719038 N DEL 5
SRR1766477.1195456 chr10 106719071 N chr10 106719138 N DEL 5
SRR1766449.8369050 chr10 106719071 N chr10 106719138 N DEL 5
SRR1766443.6792589 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766470.149485 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766476.786500 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766468.1825976 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766442.8411782 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766479.7063926 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766479.2115776 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766448.10918086 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766458.7373508 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766483.6157318 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766482.6638258 chr10 106719066 N chr10 106719133 N DEL 15
SRR1766469.6912644 chr10 106719000 N chr10 106719133 N DEL 15
SRR1766454.338703 chr10 106719000 N chr10 106719133 N DEL 15
SRR1766483.4855414 chr10 106719000 N chr10 106719133 N DEL 15
SRR1766452.6467156 chr10 106719000 N chr10 106719133 N DEL 15
SRR1766443.2265539 chr8 29667041 N chr8 29667208 N DEL 8
SRR1766483.12243578 chr8 29667041 N chr8 29667208 N DEL 8
SRR1766471.3369767 chr8 29667019 N chr8 29667116 N DUP 2
SRR1766484.7645658 chr8 29666966 N chr8 29667145 N DUP 3
SRR1766464.9895291 chr8 29666966 N chr8 29667145 N DUP 5
SRR1766483.61635 chr8 29667048 N chr8 29667117 N DEL 8
SRR1766484.4833794 chr8 29667033 N chr8 29667122 N DEL 3
SRR1766451.7593351 chr8 29667206 N chr8 29667283 N DUP 6
SRR1766470.11190758 chr8 29667216 N chr8 29667317 N DUP 13
SRR1766479.7700020 chr8 29667260 N chr8 29667315 N DUP 21
SRR1766442.6737593 chr8 29667070 N chr8 29667282 N DEL 9
SRR1766473.1063878 chr8 29666915 N chr8 29667297 N DEL 3
SRR1766461.4456442 chr8 29666962 N chr8 29667289 N DEL 11
SRR1766474.4170091 chr21 41474520 N chr21 41475903 N DEL 5
SRR1766451.5456172 chr6 158705646 N chr6 158705803 N DUP 11
SRR1766483.10479641 chr6 158705688 N chr6 158705832 N DUP 9
SRR1766458.3648309 chr6 158705688 N chr6 158705832 N DUP 9
SRR1766478.8750385 chr6 158705642 N chr6 158705801 N DEL 9
SRR1766486.3590123 chr3 5135493 N chr3 5135670 N DUP 11
SRR1766463.3020073 chr3 5135931 N chr3 5136243 N DUP 8
SRR1766462.6112610 chrX 33010119 N chrX 33010180 N DEL 18
SRR1766442.39320619 chrX 33010119 N chrX 33010180 N DEL 18
SRR1766471.1964679 chrX 33010120 N chrX 33010181 N DEL 13
SRR1766471.6413838 chrX 33010120 N chrX 33010181 N DEL 13
SRR1766455.1942686 chrX 33010095 N chrX 33010198 N DEL 10
SRR1766467.10090629 chr15 21149854 N chr15 21149933 N DUP 1
SRR1766470.7687355 chr16 75059351 N chr16 75059403 N DUP 20
SRR1766472.10295300 chr19 11153376 N chr19 11153999 N DEL 1
SRR1766443.2357380 chr19 11153376 N chr19 11153999 N DEL 8
SRR1766484.8602056 chr19 11153547 N chr19 11154171 N DUP 5
SRR1766465.7882707 chr19 11153549 N chr19 11154173 N DUP 3
SRR1766476.1632452 chr19 11153550 N chr19 11154174 N DUP 2
SRR1766457.3275109 chr19 11153551 N chr19 11154175 N DUP 1
SRR1766445.7997261 chr9 42199423 N chr9 42199552 N DEL 5
SRR1766465.3192230 chrX 123846056 N chrX 123846365 N DEL 5
SRR1766453.997981 chrX 123846064 N chrX 123846373 N DEL 10
SRR1766479.9819543 chrX 123846076 N chrX 123846383 N DUP 5
SRR1766452.7598713 chrX 123846348 N chrX 123846656 N DEL 2
SRR1766442.36498884 chr7 56367877 N chr7 56368280 N DEL 5
SRR1766477.7651209 chr7 56367950 N chr7 56368178 N DEL 5
SRR1766481.5939938 chr7 56367950 N chr7 56368096 N DEL 10
SRR1766455.5443953 chr7 56367772 N chr7 56367997 N DUP 5
SRR1766460.10648237 chr7 56367898 N chr7 56368299 N DUP 2
SRR1766459.7971264 chr7 56367943 N chr7 56368218 N DUP 5
SRR1766475.865200 chr7 56367936 N chr7 56368082 N DUP 5
SRR1766483.533353 chr7 56367860 N chr7 56368088 N DEL 11
SRR1766474.1504335 chr1 35865347 N chr1 35865651 N DEL 5
SRR1766475.4042046 chr1 35865329 N chr1 35865631 N DUP 3
SRR1766482.10232645 chr7 157057186 N chr7 157057251 N DEL 4
SRR1766455.6365799 chr7 157057113 N chr7 157057217 N DEL 5
SRR1766471.2932528 chr7 157057234 N chr7 157057377 N DUP 5
SRR1766472.10394638 chr7 157057134 N chr7 157057421 N DUP 5
SRR1766450.9562426 chr7 157057195 N chr7 157057340 N DEL 1
SRR1766442.11955018 chr7 157057373 N chr7 157057452 N DUP 5
SRR1766460.1182140 chr7 157057131 N chr7 157057420 N DEL 5
SRR1766472.5122703 chr7 157057325 N chr7 157057548 N DUP 10
SRR1766462.1570230 chr7 157057245 N chr7 157057548 N DUP 5
SRR1766463.3138776 chr7 157057310 N chr7 157057375 N DEL 5
SRR1766465.10412565 chr7 157057469 N chr7 157057548 N DUP 5
SRR1766451.2808562 chr7 157057245 N chr7 157057548 N DUP 7
SRR1766482.9014818 chr3 128954869 N chr3 128955044 N DUP 2
SRR1766469.3882093 chr3 128954864 N chr3 128955088 N DUP 5
SRR1766465.1556325 chr3 128955139 N chr3 128955495 N DUP 5
SRR1766450.3526199 chr3 128955208 N chr3 128955436 N DUP 5
SRR1766446.263932 chr3 128954879 N chr3 128955233 N DEL 5
SRR1766478.6069197 chr3 128954879 N chr3 128955233 N DEL 5
SRR1766461.11082585 chr3 128955025 N chr3 128955252 N DEL 10
SRR1766464.3991584 chr3 128955025 N chr3 128955252 N DEL 10
SRR1766462.6974829 chr3 128955030 N chr3 128955257 N DEL 5
SRR1766465.1067411 chr3 128955032 N chr3 128955259 N DEL 5
SRR1766452.3179696 chr3 128955039 N chr3 128955266 N DEL 1
SRR1766454.2532317 chr3 128955135 N chr3 128955316 N DEL 7
SRR1766484.8950616 chr3 128955044 N chr3 128955322 N DEL 3
SRR1766442.7591456 chr3 128954889 N chr3 128955342 N DEL 7
SRR1766471.4586191 chr3 128955222 N chr3 128955450 N DUP 1
SRR1766479.4083418 chr12 12944889 N chr12 12944951 N DEL 8
SRR1766457.9455848 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766442.23936417 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766463.988270 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766462.8210323 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766452.6744293 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766455.8565815 chr12 12944889 N chr12 12944951 N DEL 10
SRR1766448.10239597 chr12 12944892 N chr12 12944950 N DEL 10
SRR1766442.33013779 chr12 12944892 N chr12 12944950 N DEL 15
SRR1766479.11636452 chr12 12944896 N chr12 12944950 N DEL 12
SRR1766474.6293010 chr12 12944896 N chr12 12944950 N DEL 13
SRR1766452.6004620 chr9 96601608 N chr9 96601906 N DEL 1
SRR1766475.6040977 chr1 11145739 N chr1 11145857 N DUP 5
SRR1766478.7745262 chr10 15149213 N chr10 15149344 N DUP 5
SRR1766486.1050257 chr10 15149427 N chr10 15149682 N DEL 2
SRR1766486.5234875 chr10 15149213 N chr10 15149439 N DUP 10
SRR1766442.17362096 chr10 15149213 N chr10 15149439 N DUP 10
SRR1766475.3908330 chr10 15149487 N chr10 15149662 N DEL 5
SRR1766450.3305644 chr10 15149394 N chr10 15149506 N DUP 6
SRR1766486.8196070 chr10 15149266 N chr10 15149516 N DUP 5
SRR1766442.27007108 chr10 15149353 N chr10 15149410 N DEL 11
SRR1766478.6168211 chr10 15149418 N chr10 15149536 N DUP 9
SRR1766477.10553609 chr10 15149434 N chr10 15149549 N DUP 8
SRR1766466.3103977 chr10 15149400 N chr10 15149518 N DUP 5
SRR1766465.3435809 chr10 15149434 N chr10 15149549 N DUP 9
SRR1766462.9714871 chr10 15149414 N chr10 15149532 N DUP 7
SRR1766462.6108573 chr10 15149414 N chr10 15149532 N DUP 14
SRR1766483.3418252 chr10 15149320 N chr10 15149584 N DUP 11
SRR1766459.3240647 chr10 15149414 N chr10 15149532 N DUP 14
SRR1766484.9770339 chr10 15149414 N chr10 15149532 N DUP 18
SRR1766465.5263945 chr10 15149414 N chr10 15149532 N DUP 19
SRR1766485.3761545 chr10 15149605 N chr10 15149706 N DUP 24
SRR1766463.1853415 chr10 15149592 N chr10 15149657 N DUP 29
SRR1766480.425796 chr10 15149593 N chr10 15149658 N DUP 15
SRR1766453.3546593 chr10 15149592 N chr10 15149657 N DUP 26
SRR1766460.1628626 chr10 15149531 N chr10 15149592 N DEL 19
SRR1766447.6190164 chr10 15149464 N chr10 15149693 N DUP 17
SRR1766478.1232114 chr10 15149597 N chr10 15149698 N DUP 13
SRR1766458.7380679 chr10 15149577 N chr10 15149738 N DUP 25
SRR1766460.8561626 chr10 15149531 N chr10 15149598 N DEL 15
SRR1766450.9178643 chr10 15149531 N chr10 15149598 N DEL 16
SRR1766449.5700154 chr10 15149622 N chr10 15149690 N DUP 12
SRR1766461.6776329 chr10 15149666 N chr10 15149740 N DUP 7
SRR1766486.5771749 chr10 15149654 N chr10 15149716 N DUP 12
SRR1766445.8698855 chr10 15149345 N chr10 15149735 N DUP 14
SRR1766470.1082725 chr10 15149498 N chr10 15149628 N DEL 19
SRR1766472.3522019 chr10 15149655 N chr10 15149726 N DUP 14
SRR1766463.2112154 chr10 15149597 N chr10 15149698 N DUP 12
SRR1766446.5264582 chr10 15149481 N chr10 15149744 N DUP 9
SRR1766442.46068740 chr10 15149604 N chr10 15149708 N DUP 8
SRR1766480.3315942 chr10 15149501 N chr10 15149649 N DEL 12
SRR1766475.4714776 chr10 15149679 N chr10 15149738 N DUP 10
SRR1766486.1050257 chr10 15149601 N chr10 15149699 N DUP 17
SRR1766460.5457542 chr10 15149518 N chr10 15149597 N DEL 9
SRR1766463.5798224 chr10 15149222 N chr10 15149750 N DUP 11
SRR1766458.2349347 chr10 15149662 N chr10 15149742 N DUP 10
SRR1766481.4352701 chr10 15149230 N chr10 15149688 N DEL 3
SRR1766479.9464627 chr10 15149232 N chr10 15149690 N DEL 1
SRR1766450.3578925 chr10 15149630 N chr10 15149712 N DEL 10
SRR1766460.8561626 chr10 15149360 N chr10 15149719 N DEL 5
SRR1766463.2577476 chr10 15149619 N chr10 15149722 N DEL 5
SRR1766458.8308435 chr9 118390577 N chr9 118390778 N DUP 2
SRR1766442.11827094 chr14 104720496 N chr14 104720601 N DEL 2
SRR1766472.9746978 chr14 104720496 N chr14 104720601 N DEL 2
SRR1766442.17206080 chr14 104720558 N chr14 104720696 N DEL 5
SRR1766466.6020588 chr14 104720558 N chr14 104720696 N DEL 5
SRR1766470.7172163 chr14 104720558 N chr14 104720696 N DEL 16
SRR1766476.9015370 chr14 104720548 N chr14 104720651 N DUP 5
SRR1766450.2903937 chr14 104720548 N chr14 104720651 N DUP 5
SRR1766482.10889181 chr14 104720548 N chr14 104720651 N DUP 5
SRR1766482.9045527 chr14 104720548 N chr14 104720651 N DUP 5
SRR1766470.9390525 chr14 104720548 N chr14 104720651 N DUP 5
SRR1766454.8130397 chr14 104720548 N chr14 104720651 N DUP 5
SRR1766450.4314423 chr14 104720548 N chr14 104720651 N DUP 5
SRR1766456.3502087 chr14 104720661 N chr14 104721181 N DEL 5
SRR1766462.11216592 chr14 104720661 N chr14 104721181 N DEL 5
SRR1766442.43552980 chr14 104720532 N chr14 104720705 N DEL 6
SRR1766482.8009113 chr14 104720764 N chr14 104721006 N DEL 6
SRR1766448.6228387 chr14 104720764 N chr14 104721006 N DEL 5
SRR1766455.9730286 chr14 104720513 N chr14 104720755 N DEL 5
SRR1766443.2003789 chr14 104720764 N chr14 104721006 N DEL 7
SRR1766464.8049911 chr14 104720526 N chr14 104721009 N DEL 5
SRR1766468.4927580 chr14 104720527 N chr14 104721010 N DEL 5
SRR1766458.17230 chr14 104720509 N chr14 104720751 N DEL 7
SRR1766464.7765102 chr14 104720527 N chr14 104720941 N DEL 7
SRR1766464.3732957 chr14 104720548 N chr14 104720651 N DUP 5
SRR1766455.4255843 chr14 104720501 N chr14 104720916 N DEL 2
SRR1766458.2907655 chr14 104720522 N chr14 104720936 N DEL 7
SRR1766471.6319472 chr14 104720523 N chr14 104720937 N DEL 7
SRR1766455.4255843 chr14 104721003 N chr14 104721518 N DEL 6
SRR1766461.7718003 chr14 104720523 N chr14 104720696 N DEL 13
SRR1766457.958488 chr14 104720523 N chr14 104720903 N DEL 6
SRR1766454.8130397 chr14 104720522 N chr14 104720972 N DEL 6
SRR1766470.7353141 chr14 104720523 N chr14 104720696 N DEL 10
SRR1766446.10663172 chr14 104720523 N chr14 104721006 N DEL 5
SRR1766454.4070637 chr14 104720523 N chr14 104721006 N DEL 5
SRR1766446.8169823 chr14 104720523 N chr14 104721006 N DEL 5
SRR1766442.29458857 chr14 104720527 N chr14 104721010 N DEL 5
SRR1766450.10061137 chr14 104720533 N chr14 104721016 N DEL 5
SRR1766484.4619882 chr14 104720491 N chr14 104721208 N DUP 13
SRR1766459.10691782 chr14 104720491 N chr14 104721208 N DUP 13
SRR1766484.11737318 chr14 104720561 N chr14 104721208 N DUP 13
SRR1766448.1320047 chr14 104720601 N chr14 104721286 N DUP 10
SRR1766465.6056452 chr14 104720532 N chr14 104720630 N DUP 5
SRR1766471.6319472 chr14 104720922 N chr14 104721332 N DUP 4
SRR1766448.6103212 chr14 104720480 N chr14 104721373 N DUP 5
SRR1766465.10396959 chr14 104720575 N chr14 104721021 N DUP 1
SRR1766485.11810140 chr14 104720628 N chr14 104721450 N DUP 1
SRR1766442.41069344 chr14 104720516 N chr14 104720905 N DEL 13
SRR1766465.1675585 chr14 104720886 N chr14 104721332 N DEL 7
SRR1766478.9159002 chr14 104720564 N chr14 104721288 N DUP 5
SRR1766460.9839350 chr14 104720651 N chr14 104721475 N DEL 5
SRR1766442.24739537 chr14 104720651 N chr14 104721475 N DEL 5
SRR1766442.36347636 chr14 104720654 N chr14 104721478 N DEL 5
SRR1766453.9742371 chr14 104720675 N chr14 104721500 N DEL 2
SRR1766460.9295975 chr14 104721519 N chr14 104721587 N DUP 5
SRR1766443.3445553 chr1 2142036 N chr1 2142457 N DEL 5
SRR1766469.9620287 chr1 2142036 N chr1 2142457 N DEL 5
SRR1766482.7011433 chr1 2142095 N chr1 2142264 N DEL 5
SRR1766442.15423336 chr1 2142046 N chr1 2142299 N DEL 3
SRR1766445.2992432 chr1 2142074 N chr1 2142285 N DEL 5
SRR1766466.6178041 chr1 2142074 N chr1 2142285 N DEL 5
SRR1766449.1561701 chr1 2142074 N chr1 2142285 N DEL 5
SRR1766469.6993938 chr1 2142074 N chr1 2142285 N DEL 5
SRR1766469.1153772 chr1 2142054 N chr1 2142263 N DUP 5
SRR1766473.9986850 chr1 2142074 N chr1 2142285 N DEL 5
SRR1766475.8519840 chr1 2142074 N chr1 2142285 N DEL 5
SRR1766481.7657590 chr1 2142035 N chr1 2142288 N DEL 5
SRR1766456.4088198 chr1 2142087 N chr1 2142298 N DEL 2
SRR1766451.4416238 chr1 2142076 N chr1 2142411 N DUP 7
SRR1766453.9538600 chr1 2142069 N chr1 2142154 N DEL 5
SRR1766465.546788 chr1 2142054 N chr1 2142263 N DUP 5
SRR1766442.16107555 chr1 2142095 N chr1 2142264 N DEL 5
SRR1766449.3539188 chr1 2142022 N chr1 2142273 N DUP 5
SRR1766454.7828908 chr1 2142095 N chr1 2142264 N DEL 5
SRR1766447.5856424 chr1 2142062 N chr1 2142273 N DEL 5
SRR1766470.9194478 chr1 2142064 N chr1 2142275 N DEL 4
SRR1766459.1058799 chr1 2142088 N chr1 2142299 N DEL 5
SRR1766450.9896105 chr1 2142037 N chr1 2142290 N DEL 5
SRR1766444.6803480 chr1 2142116 N chr1 2142285 N DEL 5
SRR1766447.7716972 chr1 2142116 N chr1 2142285 N DEL 5
SRR1766471.1627380 chr1 2142116 N chr1 2142285 N DEL 5
SRR1766465.546788 chr1 2142381 N chr1 2142466 N DEL 5
SRR1766486.409004 chr1 2142074 N chr1 2142285 N DEL 5
SRR1766480.86281 chr1 2142116 N chr1 2142285 N DEL 8
SRR1766473.9986850 chr1 2142135 N chr1 2142557 N DEL 8
SRR1766477.10099352 chr1 2142035 N chr1 2142330 N DEL 1
SRR1766449.1561701 chr1 2142246 N chr1 2142457 N DEL 5
SRR1766467.8964753 chr1 2142471 N chr1 2142557 N DEL 6
SRR1766482.4266891 chr1 2142246 N chr1 2142457 N DEL 5
SRR1766455.5604169 chr1 2142173 N chr1 2142466 N DUP 6
SRR1766445.141934 chr1 2142471 N chr1 2142557 N DEL 15
SRR1766469.8249993 chr1 2142471 N chr1 2142557 N DEL 15
SRR1766467.2738637 chr1 2142414 N chr1 2142626 N DEL 8
SRR1766480.86281 chr1 2142075 N chr1 2142581 N DEL 16
SRR1766484.7670346 chr1 2142471 N chr1 2142557 N DEL 12
SRR1766453.7730850 chr1 2142471 N chr1 2142557 N DEL 14
SRR1766459.10597847 chr1 2142075 N chr1 2142581 N DEL 11
SRR1766456.6196670 chr1 2142471 N chr1 2142557 N DEL 7
SRR1766467.6325504 chr1 2142057 N chr1 2142563 N DEL 5
SRR1766475.1903748 chr1 2142099 N chr1 2142563 N DEL 9
SRR1766442.29292620 chr1 2142075 N chr1 2142581 N DEL 5
SRR1766469.7480979 chr1 2142039 N chr1 2142587 N DEL 5
SRR1766442.5473329 chr1 2142088 N chr1 2142594 N DEL 2
SRR1766455.3401840 chr1 2142089 N chr1 2142595 N DEL 1
SRR1766479.11417957 chr10 10462629 N chr10 10462784 N DUP 9
SRR1766470.5684576 chr10 10462637 N chr10 10462778 N DEL 2
SRR1766460.6359927 chr10 10462637 N chr10 10462779 N DEL 1
SRR1766467.1688184 chr10 10462637 N chr10 10462779 N DEL 1
SRR1766449.6882202 chr10 10462637 N chr10 10462777 N DEL 3
SRR1766464.8749425 chr10 10462637 N chr10 10462772 N DEL 8
SRR1766469.5569084 chr10 10462637 N chr10 10462767 N DEL 13
SRR1766470.6498967 chr10 10462637 N chr10 10462768 N DEL 12
SRR1766457.6518502 chr2 83914591 N chr2 83914660 N DEL 5
SRR1766450.5413375 chr2 83914591 N chr2 83914660 N DEL 6
SRR1766475.8180115 chr2 83914472 N chr2 83914617 N DUP 4
SRR1766484.12033461 chr2 83914554 N chr2 83914651 N DUP 8
SRR1766454.10663833 chr2 83914609 N chr2 83914757 N DUP 10
SRR1766472.11313346 chr2 83914513 N chr2 83914756 N DUP 14
SRR1766450.4542906 chr2 83914513 N chr2 83914756 N DUP 18
SRR1766469.3437505 chr2 83914553 N chr2 83914649 N DEL 8
SRR1766463.5622191 chr2 83914553 N chr2 83914649 N DEL 7
SRR1766447.10349129 chr2 83914553 N chr2 83914649 N DEL 7
SRR1766479.13786496 chr2 83914553 N chr2 83914649 N DEL 7
SRR1766473.7420994 chr2 83914554 N chr2 83914650 N DEL 7
SRR1766449.2879521 chr2 83914554 N chr2 83914650 N DEL 7
SRR1766463.10845758 chr2 83914582 N chr2 83914653 N DEL 7
SRR1766467.10901725 chr2 83914536 N chr2 83914656 N DEL 6
SRR1766466.2007458 chr2 83914591 N chr2 83914662 N DEL 2
SRR1766468.6325797 chr8 140120705 N chr8 140120870 N DEL 41
SRR1766477.11085877 chr8 140120731 N chr8 140120784 N DEL 6
SRR1766482.4114782 chr8 140120705 N chr8 140120870 N DEL 12
SRR1766473.4727613 chr8 140120804 N chr8 140120968 N DUP 5
SRR1766466.3542217 chr8 140120661 N chr8 140120970 N DUP 5
SRR1766479.11341268 chr8 140120878 N chr8 140121004 N DUP 4
SRR1766471.1081450 chr8 140120758 N chr8 140120892 N DEL 9
SRR1766465.4070334 chr8 140120706 N chr8 140121019 N DUP 5
SRR1766465.1469828 chr8 140120718 N chr8 140120964 N DEL 5
SRR1766479.5058398 chr8 140120712 N chr8 140121023 N DEL 5
SRR1766473.7101736 chr8 140120912 N chr8 140121059 N DEL 5
SRR1766465.11227638 chrX 117323959 N chrX 117324020 N DEL 7
SRR1766442.45899132 chrX 117323963 N chrX 117324024 N DEL 7
SRR1766479.4027156 chr19 37413342 N chr19 37413931 N DEL 9
SRR1766448.6778963 chr19 37413392 N chr19 37413981 N DEL 9
SRR1766481.10788732 chr19 37413828 N chr19 37414079 N DUP 5
SRR1766454.8648900 chr19 37413664 N chr19 37413917 N DEL 5
SRR1766457.3909088 chr9 83948475 N chr9 83948654 N DEL 5
SRR1766469.10169153 chr5 151650767 N chr5 151650939 N DEL 5
SRR1766447.9829239 chr16 7956972 N chr16 7957141 N DEL 3
SRR1766468.6463749 chr16 7956961 N chr16 7957132 N DEL 5
SRR1766477.2130030 chr19 36638948 N chr19 36639285 N DEL 5
SRR1766448.2455299 chr19 36638973 N chr19 36639310 N DEL 5
SRR1766454.2337188 chr4 7363561 N chr4 7363633 N DEL 5
SRR1766457.6195757 chr7 61903967 N chr7 61904479 N DUP 20
SRR1766467.7554517 chr7 61904411 N chr7 61904927 N DEL 30
SRR1766459.10524536 chr4 713396 N chr4 713574 N DEL 6
SRR1766459.805884 chr4 713574 N chr4 713627 N DEL 15
SRR1766474.8810512 chr9 134422094 N chr9 134422529 N DEL 5
SRR1766483.11669232 chr9 134422102 N chr9 134422647 N DEL 5
SRR1766485.3516091 chr9 134422270 N chr9 134422809 N DEL 8
SRR1766450.1232793 chr9 134422161 N chr9 134422290 N DUP 4
SRR1766453.7351396 chr9 134422330 N chr9 134422701 N DUP 4
SRR1766442.42495481 chr9 134422449 N chr9 134422652 N DEL 5
SRR1766465.2631222 chr9 134422474 N chr9 134422585 N DEL 6
SRR1766467.4021280 chr9 134422216 N chr9 134422409 N DEL 5
SRR1766472.5320411 chr9 134422223 N chr9 134422416 N DEL 1
SRR1766442.41340464 chr9 134422502 N chr9 134422649 N DEL 8
SRR1766483.11669232 chr9 134422466 N chr9 134422667 N DUP 3
SRR1766477.3996881 chr9 134422431 N chr9 134422760 N DEL 20
SRR1766452.2083065 chr9 134422083 N chr9 134422756 N DEL 5
SRR1766484.6145337 chr9 134422736 N chr9 134422791 N DEL 5
SRR1766481.3673602 chr9 134422087 N chr9 134422814 N DEL 4
SRR1766470.2724044 chr9 134422667 N chr9 134422830 N DEL 5
SRR1766477.10059085 chr9 134422112 N chr9 134422837 N DEL 1
SRR1766466.1861879 chr9 136307630 N chr9 136309055 N DEL 1
SRR1766486.7420566 chr9 136307772 N chr9 136308853 N DEL 6
SRR1766486.7867077 chr9 136307857 N chr9 136308336 N DEL 1
SRR1766460.2709101 chr9 136307873 N chr9 136308959 N DEL 10
SRR1766468.5250727 chr9 136307917 N chr9 136308277 N DEL 3
SRR1766442.12593267 chr9 136307993 N chr9 136309057 N DEL 5
SRR1766447.2459378 chr9 136307889 N chr9 136308418 N DUP 5
SRR1766449.8577730 chr9 136307889 N chr9 136308418 N DUP 5
SRR1766465.11138687 chr9 136307889 N chr9 136308418 N DUP 5
SRR1766459.3311665 chr9 136307753 N chr9 136307894 N DEL 8
SRR1766444.1619428 chr9 136307833 N chr9 136307896 N DEL 4
SRR1766468.2447764 chr9 136307506 N chr9 136307914 N DEL 10
SRR1766452.2701772 chr9 136307936 N chr9 136308583 N DUP 1
SRR1766458.4205770 chr9 136307625 N chr9 136307929 N DEL 5
SRR1766442.45077211 chr9 136307984 N chr9 136308074 N DUP 5
SRR1766475.1956834 chr9 136307984 N chr9 136308074 N DUP 5
SRR1766477.2740728 chr9 136308115 N chr9 136308968 N DEL 5
SRR1766453.10487929 chr9 136308044 N chr9 136308226 N DEL 14
SRR1766461.109184 chr9 136308009 N chr9 136308500 N DUP 5
SRR1766469.9529305 chr9 136307919 N chr9 136308032 N DEL 9
SRR1766484.2324684 chr9 136308028 N chr9 136308820 N DUP 5
SRR1766479.9441339 chr9 136308157 N chr9 136308616 N DEL 5
SRR1766464.5234761 chr9 136307890 N chr9 136308191 N DUP 3
SRR1766469.8541234 chr9 136308199 N chr9 136308393 N DEL 10
SRR1766453.5850425 chr9 136308089 N chr9 136308179 N DUP 2
SRR1766454.4139736 chr9 136308038 N chr9 136308219 N DUP 7
SRR1766459.264474 chr9 136307889 N chr9 136308219 N DUP 8
SRR1766484.4870893 chr9 136308038 N chr9 136308219 N DUP 7
SRR1766471.9604658 chr9 136308038 N chr9 136308219 N DUP 7
SRR1766480.7930815 chr9 136308038 N chr9 136308219 N DUP 7
SRR1766478.11013932 chr9 136308040 N chr9 136308221 N DUP 7
SRR1766484.9000563 chr9 136307980 N chr9 136308161 N DUP 12
SRR1766463.603070 chr9 136308135 N chr9 136308226 N DEL 7
SRR1766442.17445329 chr9 136307983 N chr9 136308254 N DUP 5
SRR1766448.6219012 chr9 136308135 N chr9 136308226 N DEL 7
SRR1766468.4971223 chr9 136308038 N chr9 136308219 N DUP 3
SRR1766464.1832511 chr9 136308281 N chr9 136308803 N DEL 5
SRR1766471.8432377 chr9 136308135 N chr9 136308226 N DEL 7
SRR1766463.10099757 chr9 136308044 N chr9 136308226 N DEL 17
SRR1766453.9162025 chr9 136308052 N chr9 136308234 N DEL 7
SRR1766453.5122981 chr9 136308054 N chr9 136308236 N DEL 5
SRR1766456.1203717 chr9 136308058 N chr9 136308240 N DEL 1
SRR1766480.509387 chr9 136307889 N chr9 136308361 N DUP 4
SRR1766482.12957971 chr9 136308258 N chr9 136309024 N DUP 5
SRR1766442.12593267 chr9 136307655 N chr9 136308261 N DEL 5
SRR1766448.6450734 chr9 136307490 N chr9 136308435 N DUP 10
SRR1766486.5762169 chr9 136308327 N chr9 136308544 N DUP 5
SRR1766468.7070610 chr9 136308459 N chr9 136309005 N DEL 1
SRR1766466.9760410 chr9 136308469 N chr9 136308541 N DEL 5
SRR1766448.11101830 chr9 136308277 N chr9 136308494 N DUP 5
SRR1766479.634717 chr9 136308527 N chr9 136308928 N DEL 8
SRR1766448.9661034 chr9 136307879 N chr9 136308428 N DEL 5
SRR1766456.1207086 chr9 136308524 N chr9 136308782 N DEL 26
SRR1766453.8724952 chr9 136308577 N chr9 136308729 N DEL 3
SRR1766473.9937879 chr9 136308577 N chr9 136308729 N DEL 4
SRR1766442.17445329 chr9 136308577 N chr9 136308729 N DEL 5
SRR1766463.3590186 chr9 136307485 N chr9 136308491 N DEL 1
SRR1766460.472459 chr9 136307927 N chr9 136308505 N DEL 12
SRR1766482.11133851 chr9 136308509 N chr9 136308579 N DUP 12
SRR1766486.10045348 chr9 136307938 N chr9 136308516 N DEL 4
SRR1766453.9429119 chr9 136308633 N chr9 136309162 N DEL 5
SRR1766479.9441339 chr9 136307505 N chr9 136308536 N DEL 13
SRR1766482.1942524 chr9 136307928 N chr9 136308553 N DEL 3
SRR1766453.9354321 chr9 136308547 N chr9 136309178 N DUP 15
SRR1766480.1013974 chr9 136307458 N chr9 136308577 N DEL 3
SRR1766443.4126186 chr9 136308358 N chr9 136308597 N DEL 5
SRR1766473.3228173 chr9 136308472 N chr9 136308648 N DEL 1
SRR1766460.7045752 chr9 136308026 N chr9 136308681 N DEL 9
SRR1766476.4223656 chr9 136308049 N chr9 136308695 N DEL 1
SRR1766486.8295008 chr9 136308545 N chr9 136308721 N DEL 3
SRR1766468.7070610 chr9 136308324 N chr9 136308718 N DEL 2
SRR1766470.2536131 chr9 136308307 N chr9 136308783 N DEL 10
SRR1766450.4962109 chr2 152923103 N chr2 152923271 N DUP 12
SRR1766451.7173943 chrX 71740723 N chrX 71740852 N DUP 5
SRR1766451.786606 chrX 71740804 N chrX 71741111 N DUP 4
SRR1766442.30514896 chrX 71740950 N chrX 71741021 N DEL 7
SRR1766472.1927137 chrX 71740950 N chrX 71741021 N DEL 7
SRR1766486.4217277 chrX 71740741 N chrX 71741065 N DEL 8
SRR1766452.8931481 chrX 71740761 N chrX 71741098 N DEL 11
SRR1766474.1176446 chrX 71740802 N chrX 71741152 N DEL 12
SRR1766467.8201261 chrX 71741215 N chrX 71741272 N DEL 6
SRR1766474.6727292 chrX 71741215 N chrX 71741272 N DEL 11
SRR1766464.2059664 chr19 20149842 N chr19 20149939 N DUP 2
SRR1766484.728909 chr19 20149876 N chr19 20150051 N DUP 5
SRR1766479.5645037 chr19 20149848 N chr19 20150025 N DEL 5
SRR1766473.8999509 chr19 20149915 N chr19 20150140 N DUP 1
SRR1766476.1928590 chr19 20149862 N chr19 20150039 N DEL 1
SRR1766451.3763295 chr19 20149956 N chr19 20150084 N DEL 10
SRR1766485.3725591 chr16 49210592 N chr16 49210826 N DEL 5
SRR1766445.10039870 chr1 86111253 N chr1 86111373 N DEL 4
SRR1766475.7317997 chr1 86111253 N chr1 86111373 N DEL 4
SRR1766474.10888272 chr1 86111253 N chr1 86111373 N DEL 10
SRR1766453.9487667 chr1 86111251 N chr1 86111328 N DUP 5
SRR1766446.6611307 chr1 86111215 N chr1 86111333 N DUP 5
SRR1766464.4797955 chr1 86111215 N chr1 86111333 N DUP 5
SRR1766450.8148628 chr1 86111297 N chr1 86111415 N DUP 10
SRR1766467.4074967 chr16 16350501 N chr16 16350628 N DEL 5
SRR1766465.6822460 chr6 140064306 N chr6 140064419 N DEL 2
SRR1766445.8352031 chr6 140064306 N chr6 140064417 N DEL 4
SRR1766444.4894844 chr6 140064306 N chr6 140064407 N DEL 14
SRR1766485.9700657 chr6 140064306 N chr6 140064415 N DEL 6
SRR1766444.5407570 chr9 107729163 N chr9 107729479 N DEL 9
SRR1766449.9087558 chr9 107729048 N chr9 107729364 N DEL 10
SRR1766461.9693040 chr9 107729083 N chr9 107729399 N DEL 10
SRR1766479.4315403 chr19 14002226 N chr19 14002406 N DEL 5
SRR1766479.2970189 chr19 14002241 N chr19 14002421 N DEL 5
SRR1766445.4657924 chr19 14002233 N chr19 14002583 N DEL 30
SRR1766450.6158500 chr19 14002209 N chr19 14002559 N DEL 16
SRR1766462.712330 chr19 14002341 N chr19 14002512 N DEL 3
SRR1766457.9222834 chr19 14002167 N chr19 14002517 N DEL 5
SRR1766468.5360922 chr20 22762290 N chr20 22762429 N DEL 5
SRR1766472.8993461 chr20 22762322 N chr20 22762437 N DEL 17
SRR1766447.9500600 chr20 22762292 N chr20 22762491 N DUP 7
SRR1766485.9512612 chr20 22762292 N chr20 22762491 N DUP 8
SRR1766458.4621323 chr20 22762480 N chr20 22762535 N DEL 1
SRR1766477.63389 chr20 22762323 N chr20 22762518 N DEL 5
SRR1766442.45298400 chr17 78465483 N chr17 78465638 N DUP 5
SRR1766472.586247 chr17 78465717 N chr17 78465793 N DUP 5
SRR1766471.3374555 chr17 78465889 N chr17 78465985 N DUP 1
SRR1766477.4925378 chr10 100525781 N chr10 100525866 N DUP 18
SRR1766474.10648682 chr10 100525783 N chr10 100525866 N DUP 23
SRR1766483.3724836 chr10 100525778 N chr10 100525897 N DEL 1
SRR1766448.6033794 chrY 56832640 N chrY 56832691 N DEL 13
SRR1766442.38311926 chrY 56832624 N chrY 56832703 N DUP 11
SRR1766474.7068363 chrY 56832502 N chrY 56832678 N DUP 1
SRR1766486.6418731 chrY 56832505 N chrY 56832676 N DUP 2
SRR1766444.6432607 chrY 56832482 N chrY 56832663 N DUP 5
SRR1766482.9979460 chrY 56832516 N chrY 56832689 N DEL 5
SRR1766484.11243453 chrY 56832668 N chrY 56832866 N DEL 1
SRR1766455.3415925 chrY 56832521 N chrY 56832689 N DEL 9
SRR1766442.26244332 chrY 56832501 N chrY 56832672 N DUP 4
SRR1766479.10093370 chrY 56832521 N chrY 56832689 N DEL 12
SRR1766469.8651742 chrY 56832541 N chrY 56832637 N DUP 5
SRR1766442.31466519 chrY 56832624 N chrY 56832703 N DUP 13
SRR1766475.8007632 chrY 56832533 N chrY 56832646 N DEL 15
SRR1766454.1477437 chrY 56832632 N chrY 56832686 N DUP 5
SRR1766479.8201704 chrY 56832627 N chrY 56832828 N DUP 1
SRR1766466.2012533 chrY 56832479 N chrY 56832667 N DEL 10
SRR1766463.5068019 chrY 56832638 N chrY 56832694 N DEL 10
SRR1766475.2164559 chrY 56832624 N chrY 56832703 N DUP 11
SRR1766466.7735684 chrY 56832505 N chrY 56832676 N DUP 3
SRR1766485.3371475 chrY 56832536 N chrY 56832704 N DEL 2
SRR1766471.11010484 chrY 56832501 N chrY 56832672 N DUP 5
SRR1766442.4626513 chrY 56832479 N chrY 56832697 N DEL 2
SRR1766452.9900474 chrY 56832518 N chrY 56832696 N DEL 3
SRR1766458.8372337 chrY 56832501 N chrY 56832672 N DUP 10
SRR1766442.11752887 chrY 56832521 N chrY 56832694 N DEL 5
SRR1766442.27326158 chrY 56832625 N chrY 56832808 N DEL 1
SRR1766478.5573406 chrY 56832518 N chrY 56832691 N DEL 5
SRR1766475.1481515 chrY 56832521 N chrY 56832694 N DEL 5
SRR1766462.9955769 chrY 56832526 N chrY 56832694 N DEL 15
SRR1766451.4929332 chrY 56832537 N chrY 56832723 N DUP 4
SRR1766486.8525340 chrY 56832502 N chrY 56832658 N DUP 18
SRR1766485.9780615 chrY 56832502 N chrY 56832678 N DUP 5
SRR1766486.72152 chrY 56832526 N chrY 56832637 N DUP 4
SRR1766485.2749192 chrY 56832480 N chrY 56832693 N DEL 5
SRR1766463.6734647 chrY 56832526 N chrY 56832674 N DEL 15
SRR1766483.8270574 chrY 56832638 N chrY 56832699 N DEL 5
SRR1766477.9933165 chrY 56832641 N chrY 56832702 N DEL 5
SRR1766478.3281477 chrY 56832639 N chrY 56832700 N DEL 4
SRR1766465.6276068 chrY 56832516 N chrY 56832689 N DEL 5
SRR1766465.129010 chrY 56832628 N chrY 56832806 N DEL 8
SRR1766454.7585016 chrY 56832502 N chrY 56832678 N DUP 5
SRR1766484.2910610 chrY 56832536 N chrY 56832694 N DEL 8
SRR1766445.10308449 chrY 56832502 N chrY 56832688 N DUP 18
SRR1766448.9488299 chrY 56832625 N chrY 56832694 N DUP 5
SRR1766459.7148932 chrY 56832521 N chrY 56832694 N DEL 5
SRR1766468.2839629 chrY 56832521 N chrY 56832689 N DEL 9
SRR1766457.9295719 chrY 56832521 N chrY 56832689 N DEL 6
SRR1766483.9136165 chrY 56832521 N chrY 56832689 N DEL 10
SRR1766477.10570622 chrY 56832615 N chrY 56832679 N DUP 5
SRR1766470.5725053 chrY 56832502 N chrY 56832678 N DUP 5
SRR1766473.6377599 chrY 56832692 N chrY 56832828 N DUP 3
SRR1766452.7235622 chrY 56832515 N chrY 56832648 N DEL 8
SRR1766460.6140139 chrY 56832502 N chrY 56832678 N DUP 9
SRR1766457.7921007 chrY 56832536 N chrY 56832704 N DEL 1
SRR1766471.3819600 chrY 56832638 N chrY 56832699 N DEL 5
SRR1766451.7460928 chrY 56832639 N chrY 56832700 N DEL 4
SRR1766473.9665699 chrY 56832502 N chrY 56832678 N DUP 4
SRR1766443.3522593 chrY 56832541 N chrY 56832637 N DUP 5
SRR1766459.3971472 chrY 56832516 N chrY 56832689 N DEL 5
SRR1766470.2415744 chrY 56832505 N chrY 56832676 N DUP 4
SRR1766442.15898942 chrY 56832527 N chrY 56832820 N DUP 3
SRR1766448.9731267 chrY 56832639 N chrY 56832700 N DEL 4
SRR1766448.221779 chrY 56832541 N chrY 56832637 N DUP 5
SRR1766442.17120129 chrY 56832503 N chrY 56832649 N DUP 6
SRR1766443.4851682 chrY 56832516 N chrY 56832694 N DEL 5
SRR1766479.10303115 chrY 56832521 N chrY 56832689 N DEL 15
SRR1766484.11567279 chrY 56832536 N chrY 56832694 N DEL 10
SRR1766457.1794972 chrY 56832502 N chrY 56832678 N DUP 4
SRR1766467.11107821 chrY 56832512 N chrY 56832663 N DUP 3
SRR1766478.3691734 chrY 56832638 N chrY 56832694 N DEL 10
SRR1766478.3374520 chrY 56832517 N chrY 56832690 N DEL 5
SRR1766466.10126700 chrY 56832640 N chrY 56832701 N DEL 3
SRR1766452.8104357 chrY 56832527 N chrY 56832820 N DUP 3
SRR1766465.7381685 chrY 56832638 N chrY 56832699 N DEL 5
SRR1766442.15505116 chrY 56832625 N chrY 56832694 N DUP 5
SRR1766453.5125318 chrY 56832639 N chrY 56832700 N DEL 4
SRR1766456.4773548 chrY 56832541 N chrY 56832637 N DUP 5
SRR1766486.566765 chrY 56832521 N chrY 56832689 N DEL 8
SRR1766477.10034290 chrY 56832521 N chrY 56832689 N DEL 9
SRR1766484.4156069 chrY 56832633 N chrY 56832866 N DEL 6
SRR1766442.45774751 chrY 56832497 N chrY 56832645 N DEL 10
SRR1766486.1471825 chrY 56832642 N chrY 56832693 N DEL 11
SRR1766466.7808909 chr4 117720751 N chr4 117720812 N DEL 10
SRR1766442.24019877 chr4 117720752 N chr4 117720813 N DEL 9
SRR1766454.3218652 chr4 117720753 N chr4 117720814 N DEL 9
SRR1766454.6326349 chr4 117720753 N chr4 117720814 N DEL 9
SRR1766482.12311138 chr4 117720763 N chr4 117720824 N DEL 2
SRR1766464.1294522 chr20 7435684 N chr20 7435764 N DEL 4
SRR1766469.7618563 chr20 7435684 N chr20 7435764 N DEL 4
SRR1766461.7091329 chr20 7435684 N chr20 7435764 N DEL 5
SRR1766485.6757061 chr20 7435684 N chr20 7435764 N DEL 8
SRR1766448.7879238 chr20 7435649 N chr20 7435727 N DUP 9
SRR1766479.2587893 chr20 7435649 N chr20 7435727 N DUP 10
SRR1766483.4645820 chr20 7435646 N chr20 7435724 N DUP 10
SRR1766452.9837535 chr20 7435649 N chr20 7435727 N DUP 10
SRR1766457.9327095 chr20 7435649 N chr20 7435727 N DUP 10
SRR1766460.1446938 chr20 7435649 N chr20 7435727 N DUP 10
SRR1766451.9451264 chr20 7435646 N chr20 7435724 N DUP 9
SRR1766470.1923036 chr20 7435646 N chr20 7435724 N DUP 11
SRR1766484.4910515 chr20 7435646 N chr20 7435724 N DUP 11
SRR1766483.10479412 chr20 7435649 N chr20 7435727 N DUP 14
SRR1766476.980463 chr20 7435646 N chr20 7435724 N DUP 15
SRR1766473.5591225 chr20 7435649 N chr20 7435727 N DUP 15
SRR1766478.6252182 chr20 7435647 N chr20 7435809 N DUP 7
SRR1766450.3199741 chr20 7435564 N chr20 7435649 N DEL 11
SRR1766454.10202566 chr20 7435687 N chr20 7435800 N DUP 21
SRR1766461.585810 chr20 7435687 N chr20 7435800 N DUP 21
SRR1766475.5692948 chr20 7435687 N chr20 7435800 N DUP 21
SRR1766453.5504645 chr20 7435687 N chr20 7435800 N DUP 21
SRR1766443.311436 chr20 7435654 N chr20 7435773 N DUP 5
SRR1766451.6086716 chr20 7435716 N chr20 7435799 N DUP 11
SRR1766464.10206603 chr20 7435716 N chr20 7435799 N DUP 14
SRR1766470.4212007 chr20 7435716 N chr20 7435799 N DUP 13
SRR1766443.10559064 chr20 7435666 N chr20 7435787 N DUP 9
SRR1766456.5998792 chr20 7435716 N chr20 7435799 N DUP 14
SRR1766443.4427402 chr20 7435716 N chr20 7435799 N DUP 16
SRR1766467.9584497 chr20 7435666 N chr20 7435787 N DUP 11
SRR1766442.7553470 chr20 7435565 N chr20 7435691 N DEL 11
SRR1766472.4935429 chr20 7435564 N chr20 7435690 N DEL 12
SRR1766460.344135 chr6 31773851 N chr6 31774159 N DEL 6
SRR1766456.4351115 chr18 2503138 N chr18 2503241 N DUP 13
SRR1766465.2727385 chr18 2503137 N chr18 2503240 N DUP 14
SRR1766462.936562 chr18 2503140 N chr18 2503243 N DUP 11
SRR1766471.11903613 chr18 2503139 N chr18 2503242 N DUP 12
SRR1766452.7797528 chr8 30767739 N chr8 30767872 N DUP 2
SRR1766452.7797528 chr8 30767881 N chr8 30768056 N DEL 4
SRR1766454.6023189 chr8 142127818 N chr8 142127929 N DUP 1
SRR1766458.1792935 chr3 129818550 N chr3 129818726 N DEL 9
SRR1766479.8949503 chr3 129818550 N chr3 129818726 N DEL 10
SRR1766460.8110663 chr3 129818550 N chr3 129818726 N DEL 10
SRR1766455.1902287 chr3 129818550 N chr3 129818726 N DEL 14
SRR1766448.5035490 chr3 129818551 N chr3 129818702 N DEL 3
SRR1766468.2583838 chr3 129818552 N chr3 129818703 N DEL 4
SRR1766459.10215504 chr3 129818554 N chr3 129818705 N DEL 6
SRR1766448.10218172 chr3 129818561 N chr3 129818712 N DEL 4
SRR1766474.1866702 chr3 129818563 N chr3 129818714 N DEL 2
SRR1766458.7446049 chr3 129818557 N chr3 129818733 N DEL 8
SRR1766471.8016846 chr7 21377602 N chr7 21377773 N DUP 1
SRR1766442.43691869 chr7 21377648 N chr7 21377706 N DEL 5
SRR1766479.6287562 chr10 3786001 N chr10 3786076 N DEL 5
SRR1766483.5105136 chr10 3786002 N chr10 3786077 N DEL 5
SRR1766476.8503507 chr5 15411073 N chr5 15411139 N DEL 6
SRR1766454.7017368 chr10 74695622 N chr10 74695754 N DUP 1
SRR1766459.1296593 chr10 74695623 N chr10 74695769 N DUP 4
SRR1766474.4737281 chr10 97528330 N chr10 97528825 N DUP 5
SRR1766457.694704 chr10 97528346 N chr10 97528941 N DUP 5
SRR1766461.8396779 chr10 97528346 N chr10 97528941 N DUP 5
SRR1766460.6816562 chr10 97528427 N chr10 97529024 N DEL 7
SRR1766442.42396860 chr10 97528270 N chr10 97528445 N DUP 1
SRR1766442.21803889 chr10 97528270 N chr10 97528445 N DUP 2
SRR1766462.903279 chr10 97528270 N chr10 97528445 N DUP 2
SRR1766449.7857778 chr10 97528346 N chr10 97528569 N DUP 5
SRR1766453.2999338 chr10 97528263 N chr10 97528438 N DUP 9
SRR1766451.7535987 chr10 97528346 N chr10 97528569 N DUP 5
SRR1766485.7318057 chr10 97528346 N chr10 97528569 N DUP 5
SRR1766459.8595727 chr10 97528280 N chr10 97528454 N DUP 5
SRR1766459.9280978 chr10 97528280 N chr10 97528454 N DUP 5
SRR1766447.9472493 chr10 97528280 N chr10 97528454 N DUP 5
SRR1766455.9063861 chr10 97528410 N chr10 97528633 N DUP 5
SRR1766482.6437712 chr10 97528266 N chr10 97528489 N DUP 4
SRR1766461.6413901 chr10 97528266 N chr10 97528489 N DUP 5
SRR1766486.7919190 chr10 97528266 N chr10 97528489 N DUP 5
SRR1766459.7798327 chr10 97528266 N chr10 97528713 N DUP 10
SRR1766464.6723733 chr10 97528266 N chr10 97528489 N DUP 5
SRR1766442.7710854 chr10 97528266 N chr10 97528489 N DUP 5
SRR1766448.7387847 chr10 97528266 N chr10 97528489 N DUP 5
SRR1766474.9418331 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766486.11765817 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766463.3387578 chr10 97528460 N chr10 97528828 N DUP 5
SRR1766478.10634670 chr10 97528269 N chr10 97528542 N DUP 12
SRR1766447.6853971 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766481.11789013 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766451.933543 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766464.3514000 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766485.4316907 chr10 97528285 N chr10 97528462 N DEL 12
SRR1766459.11373543 chr10 97528462 N chr10 97529058 N DUP 5
SRR1766443.5256016 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766450.9369262 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766442.29192102 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766480.8724002 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766482.8103838 chr10 97528318 N chr10 97528494 N DEL 10
SRR1766449.10959511 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766482.3121676 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766442.38007697 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766478.3385295 chr10 97528742 N chr10 97528891 N DEL 10
SRR1766457.694704 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766442.7522057 chr10 97528502 N chr10 97528875 N DEL 5
SRR1766460.10167645 chr10 97528283 N chr10 97528508 N DEL 1
SRR1766485.5542960 chr10 97528301 N chr10 97528526 N DEL 5
SRR1766447.3297753 chr10 97528301 N chr10 97528526 N DEL 5
SRR1766465.9256580 chr10 97528301 N chr10 97528526 N DEL 5
SRR1766442.30163700 chr10 97528312 N chr10 97528537 N DEL 4
SRR1766466.5433112 chr10 97528314 N chr10 97528539 N DEL 2
SRR1766476.2602257 chr10 97528280 N chr10 97528554 N DEL 5
SRR1766466.7640524 chr10 97528669 N chr10 97529042 N DEL 3
SRR1766475.7116546 chr10 97528283 N chr10 97528681 N DUP 5
SRR1766442.31550173 chr10 97528280 N chr10 97528678 N DUP 5
SRR1766476.5385921 chr10 97528410 N chr10 97528633 N DUP 2
SRR1766481.7122630 chr10 97528713 N chr10 97528811 N DEL 1
SRR1766463.10183971 chr10 97528410 N chr10 97528633 N DUP 5
SRR1766472.10435807 chr10 97528266 N chr10 97528713 N DUP 7
SRR1766471.10122187 chr10 97528266 N chr10 97528713 N DUP 10
SRR1766459.7798327 chr10 97528266 N chr10 97528713 N DUP 10
SRR1766447.6587341 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766455.1609261 chr10 97528501 N chr10 97528726 N DEL 5
SRR1766466.4707542 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766442.21617368 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766446.5274089 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766453.7178381 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766459.544123 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766472.662253 chr10 97528461 N chr10 97528781 N DUP 5
SRR1766486.10015861 chr10 97528461 N chr10 97528781 N DUP 6
SRR1766452.2676140 chr10 97528522 N chr10 97528747 N DEL 10
SRR1766442.35961471 chr10 97528298 N chr10 97528747 N DEL 10
SRR1766443.3835791 chr10 97528781 N chr10 97528832 N DEL 7
SRR1766454.2360020 chr10 97528776 N chr10 97528827 N DEL 11
SRR1766461.2334760 chr10 97528263 N chr10 97528857 N DUP 1
SRR1766442.4698095 chr10 97528558 N chr10 97528930 N DUP 6
SRR1766454.3364077 chr10 97528327 N chr10 97528826 N DEL 7
SRR1766462.6602921 chr10 97528327 N chr10 97528826 N DEL 7
SRR1766465.3078363 chr10 97528327 N chr10 97528826 N DEL 7
SRR1766479.7559003 chr10 97528489 N chr10 97528861 N DEL 7
SRR1766485.1261982 chr10 97528717 N chr10 97528963 N DUP 5
SRR1766473.4108898 chr10 97528489 N chr10 97528861 N DEL 10
SRR1766482.7666020 chr10 97528554 N chr10 97528875 N DUP 5
SRR1766443.6706448 chr10 97528326 N chr10 97528874 N DEL 6
SRR1766479.9423446 chr10 97528326 N chr10 97528874 N DEL 6
SRR1766481.3648221 chr10 97528283 N chr10 97528880 N DEL 5
SRR1766464.7703393 chr10 97528292 N chr10 97528889 N DEL 1
SRR1766463.7342927 chr10 97528292 N chr10 97528889 N DEL 1
SRR1766462.6602921 chr10 97528346 N chr10 97528941 N DUP 5
SRR1766465.6038375 chr10 97528308 N chr10 97528533 N DEL 5
SRR1766452.3044930 chr10 97528346 N chr10 97528941 N DUP 5
SRR1766452.2630857 chr10 97528346 N chr10 97528941 N DUP 5
SRR1766482.3121676 chr10 97528828 N chr10 97528929 N DEL 5
SRR1766475.982098 chr10 97528298 N chr10 97528944 N DEL 5
SRR1766450.2325619 chr10 97528330 N chr10 97529050 N DUP 11
SRR1766463.7890113 chr10 97528429 N chr10 97529026 N DEL 5
SRR1766451.6065250 chr10 97528270 N chr10 97529088 N DUP 1
SRR1766483.4507615 chr10 97528831 N chr10 97529059 N DEL 5
SRR1766472.4878735 chr10 97528405 N chr10 97529250 N DUP 10
SRR1766483.9019743 chr18 46546536 N chr18 46546667 N DEL 3
SRR1766470.10294740 chr3 184414636 N chr3 184414785 N DEL 12
SRR1766479.13137944 chr3 184414761 N chr3 184414915 N DEL 7
SRR1766449.5866435 chr3 184414761 N chr3 184414915 N DEL 10
SRR1766482.11599982 chr3 184414763 N chr3 184414888 N DEL 25
SRR1766483.6629982 chr3 184414763 N chr3 184414888 N DEL 43
SRR1766442.1638286 chr3 184414930 N chr3 184414994 N DEL 1
SRR1766453.10053538 chr3 184414955 N chr3 184415048 N DEL 5
SRR1766472.4608855 chr3 184414961 N chr3 184415050 N DEL 13
SRR1766453.9313997 chr3 184414629 N chr3 184415071 N DEL 2
SRR1766468.1279516 chr19 42370669 N chr19 42370780 N DEL 1
SRR1766482.9523995 chr1 9549482 N chr1 9549658 N DEL 5
SRR1766461.7685584 chr12 40773785 N chr12 40773846 N DEL 5
SRR1766450.8091176 chr12 40773785 N chr12 40773846 N DEL 8
SRR1766442.7352387 chr12 40773785 N chr12 40773846 N DEL 10
SRR1766472.7203057 chr12 40773785 N chr12 40773846 N DEL 14
SRR1766443.2546600 chr12 40773791 N chr12 40773852 N DEL 9
SRR1766444.5456784 chr12 40773794 N chr12 40773855 N DEL 6
SRR1766462.8851844 chr12 40773794 N chr12 40773855 N DEL 6
SRR1766477.4198063 chr12 40773795 N chr12 40773856 N DEL 5
SRR1766482.195527 chr12 40773796 N chr12 40773857 N DEL 4
SRR1766467.1267319 chr12 40773794 N chr12 40773855 N DEL 6
SRR1766467.2441763 chr12 40773794 N chr12 40773855 N DEL 6
SRR1766467.9983187 chr12 40773791 N chr12 40773852 N DEL 9
SRR1766473.2772632 chr12 40773787 N chr12 40773848 N DEL 13
SRR1766452.5319159 chrX 532911 N chrX 533084 N DUP 10
SRR1766479.3812222 chrX 532911 N chrX 533084 N DUP 10
SRR1766459.6091257 chrX 532358 N chrX 532698 N DUP 25
SRR1766461.6522231 chrX 532736 N chrX 532905 N DEL 20
SRR1766477.8092036 chrX 532736 N chrX 532905 N DEL 20
SRR1766442.31760687 chrX 532358 N chrX 532698 N DUP 25
SRR1766459.10428374 chrX 532395 N chrX 532905 N DEL 5
SRR1766459.8470207 chrX 532911 N chrX 533084 N DUP 10
SRR1766461.7756351 chrX 532911 N chrX 533084 N DUP 10
SRR1766461.7307005 chrX 532911 N chrX 533084 N DUP 10
SRR1766470.10824691 chrX 532736 N chrX 532905 N DEL 20
SRR1766471.8122851 chrX 532395 N chrX 532905 N DEL 5
SRR1766457.9194010 chrX 532736 N chrX 532905 N DEL 20
SRR1766472.9522075 chrX 532910 N chrX 533083 N DUP 10
SRR1766442.4712355 chrX 532736 N chrX 532905 N DEL 20
SRR1766448.7771131 chrX 532736 N chrX 532905 N DEL 20
SRR1766476.5803771 chrX 532395 N chrX 532905 N DEL 5
SRR1766480.2328076 chrX 532395 N chrX 532905 N DEL 5
SRR1766455.2629016 chrX 532736 N chrX 532905 N DEL 18
SRR1766446.1965177 chrX 532736 N chrX 532905 N DEL 17
SRR1766460.9147976 chrX 532492 N chrX 532846 N DEL 21
SRR1766458.1053295 chrX 532498 N chrX 532846 N DEL 13
SRR1766459.408763 chrX 532492 N chrX 532846 N DEL 25
SRR1766455.8427191 chrX 532616 N chrX 532938 N DEL 5
SRR1766442.37256079 chrX 532616 N chrX 532938 N DEL 5
SRR1766478.856559 chrX 532616 N chrX 532938 N DEL 5
SRR1766478.7152973 chrX 532616 N chrX 532938 N DEL 5
SRR1766474.1664745 chrX 532616 N chrX 532938 N DEL 5
SRR1766464.5201002 chrX 532334 N chrX 532489 N DUP 38
SRR1766455.161523 chrX 532358 N chrX 532698 N DUP 5
SRR1766451.2428632 chrX 532406 N chrX 532746 N DUP 1
SRR1766448.211756 chrX 532358 N chrX 532698 N DUP 9
SRR1766450.6752566 chrX 532358 N chrX 532698 N DUP 12
SRR1766484.10044483 chrX 532358 N chrX 532698 N DUP 12
SRR1766483.6348287 chrX 532358 N chrX 532698 N DUP 14
SRR1766477.4200360 chrX 532358 N chrX 532698 N DUP 25
SRR1766447.6321340 chrX 532358 N chrX 532698 N DUP 25
SRR1766470.6796442 chrX 532358 N chrX 532698 N DUP 25
SRR1766442.45090361 chrX 532358 N chrX 532698 N DUP 25
SRR1766448.8150322 chrX 532358 N chrX 532698 N DUP 25
SRR1766450.3143119 chrX 532358 N chrX 532698 N DUP 25
SRR1766474.4455774 chrX 532358 N chrX 532698 N DUP 25
SRR1766479.12130205 chrX 532358 N chrX 532698 N DUP 30
SRR1766484.10425771 chrX 532358 N chrX 532698 N DUP 30
SRR1766483.2085544 chrX 532358 N chrX 532698 N DUP 31
SRR1766485.8417833 chrX 532358 N chrX 532698 N DUP 31
SRR1766443.9657364 chrX 532358 N chrX 532698 N DUP 32
SRR1766442.34448767 chrX 532358 N chrX 532698 N DUP 32
SRR1766459.7002795 chrX 532814 N chrX 532984 N DUP 21
SRR1766478.9997886 chrX 532846 N chrX 533001 N DUP 27
SRR1766471.11981734 chrX 532846 N chrX 533001 N DUP 27
SRR1766472.6611511 chrX 532846 N chrX 533001 N DUP 27
SRR1766476.9652760 chrX 532814 N chrX 532984 N DUP 21
SRR1766483.9362901 chrX 532814 N chrX 532984 N DUP 21
SRR1766457.624091 chrX 532846 N chrX 533001 N DUP 27
SRR1766486.9501071 chrX 532814 N chrX 532984 N DUP 21
SRR1766468.7416564 chrX 532846 N chrX 533001 N DUP 24
SRR1766469.2266229 chrX 532846 N chrX 533001 N DUP 24
SRR1766442.17972795 chrX 532814 N chrX 532987 N DUP 21
SRR1766470.10694971 chrX 532814 N chrX 532984 N DUP 11
SRR1766475.3914026 chrX 532334 N chrX 532836 N DUP 16
SRR1766471.7625282 chrX 532334 N chrX 532836 N DUP 16
SRR1766468.3061584 chrX 532489 N chrX 532825 N DEL 4
SRR1766451.5814113 chrX 532334 N chrX 532836 N DUP 11
SRR1766455.1843895 chrX 532334 N chrX 532495 N DUP 10
SRR1766466.741586 chrX 532402 N chrX 533084 N DUP 15
SRR1766479.12130205 chrX 532334 N chrX 532489 N DUP 10
SRR1766452.9736373 chrX 532358 N chrX 532698 N DUP 28
SRR1766482.3287684 chrX 532688 N chrX 532857 N DEL 10
SRR1766442.42037449 chrX 532402 N chrX 533084 N DUP 15
SRR1766451.2837471 chrX 532338 N chrX 532487 N DUP 10
SRR1766462.325216 chrX 532770 N chrX 532937 N DUP 10
SRR1766463.2937286 chrX 532963 N chrX 533138 N DEL 2
SRR1766481.5743445 chrX 532913 N chrX 533086 N DUP 5
SRR1766479.7259905 chrX 532910 N chrX 533083 N DUP 15
SRR1766477.911756 chrX 532508 N chrX 532853 N DEL 5
SRR1766447.7195572 chrX 532963 N chrX 533138 N DEL 5
SRR1766485.7632539 chrX 532736 N chrX 532905 N DEL 23
SRR1766485.8417833 chrX 532880 N chrX 533053 N DUP 15
SRR1766448.8150322 chrX 532911 N chrX 533084 N DUP 11
SRR1766479.7224712 chrX 532348 N chrX 532858 N DEL 3
SRR1766476.5417712 chrX 532348 N chrX 532858 N DEL 3
SRR1766483.8662027 chrX 532911 N chrX 533084 N DUP 10
SRR1766455.8427191 chrX 532405 N chrX 532915 N DEL 5
SRR1766465.10786183 chrX 532736 N chrX 532905 N DEL 20
SRR1766447.4543671 chrX 532911 N chrX 533084 N DUP 10
SRR1766470.10694971 chrX 532964 N chrX 533139 N DEL 5
SRR1766477.3122202 chrX 532963 N chrX 533138 N DEL 5
SRR1766449.5255823 chrX 532736 N chrX 532905 N DEL 20
SRR1766481.6379179 chrX 532905 N chrX 533078 N DUP 15
SRR1766449.6873246 chrX 532963 N chrX 533138 N DEL 5
SRR1766478.8490390 chrX 532963 N chrX 533138 N DEL 5
SRR1766462.4987836 chrX 532360 N chrX 532868 N DUP 5
SRR1766451.9448856 chrX 532405 N chrX 532915 N DEL 5
SRR1766463.4414053 chrX 532485 N chrX 532981 N DUP 1
SRR1766459.6091257 chrX 532371 N chrX 532535 N DUP 5
SRR1766483.2085544 chrX 532905 N chrX 533078 N DUP 10
SRR1766442.4712355 chrX 532535 N chrX 532880 N DEL 5
SRR1766442.45090361 chrX 532911 N chrX 533084 N DUP 15
SRR1766486.1970114 chrX 532911 N chrX 533084 N DUP 15
SRR1766463.5423529 chrX 532910 N chrX 533083 N DUP 15
SRR1766445.5901442 chrX 532396 N chrX 532906 N DEL 3
SRR1766482.5839177 chrX 532476 N chrX 532981 N DUP 1
SRR1766470.10824691 chrX 532476 N chrX 532981 N DUP 6
SRR1766442.37256079 chrX 532478 N chrX 532814 N DEL 4
SRR1766473.6477425 chrX 532334 N chrX 533004 N DUP 8
SRR1766459.5797587 chrX 532911 N chrX 533084 N DUP 10
SRR1766448.847277 chrX 532473 N chrX 532987 N DUP 4
SRR1766452.2924394 chrX 532911 N chrX 533084 N DUP 10
SRR1766463.2794026 chrX 532477 N chrX 532990 N DEL 5
SRR1766449.8737437 chrX 532477 N chrX 532816 N DEL 11
SRR1766455.7942497 chrX 532477 N chrX 532816 N DEL 11
SRR1766459.5079220 chrX 532477 N chrX 532816 N DEL 13
SRR1766467.3456470 chrX 532477 N chrX 532990 N DEL 8
SRR1766471.11981734 chrX 532478 N chrX 532814 N DEL 9
SRR1766484.10425771 chrX 532477 N chrX 532816 N DEL 18
SRR1766442.45639657 chrX 532911 N chrX 533084 N DUP 10
SRR1766460.2188702 chrX 532477 N chrX 532816 N DEL 18
SRR1766461.6522231 chrX 532911 N chrX 533084 N DUP 10
SRR1766470.6796442 chrX 532477 N chrX 532816 N DEL 18
SRR1766445.5797316 chrX 532477 N chrX 532990 N DEL 8
SRR1766464.10919875 chrX 532454 N chrX 532796 N DEL 9
SRR1766481.451998 chrX 532408 N chrX 532918 N DEL 2
SRR1766477.11445418 chrX 532846 N chrX 533001 N DUP 33
SRR1766481.7843412 chrX 532846 N chrX 533001 N DUP 33
SRR1766448.4524579 chrX 532814 N chrX 532987 N DUP 15
SRR1766457.2827369 chrX 532814 N chrX 532984 N DUP 23
SRR1766481.10632956 chrX 532846 N chrX 533001 N DUP 32
SRR1766454.3179782 chrX 532814 N chrX 532987 N DUP 15
SRR1766477.11106464 chrX 532814 N chrX 532987 N DUP 25
SRR1766462.4664999 chrX 532814 N chrX 532987 N DUP 25
SRR1766443.5911404 chrX 532814 N chrX 532987 N DUP 25
SRR1766447.4543671 chrX 532334 N chrX 533004 N DUP 20
SRR1766451.4329360 chrX 532334 N chrX 533004 N DUP 20
SRR1766442.41208733 chrX 532813 N chrX 532988 N DEL 11
SRR1766476.7169450 chrX 532813 N chrX 532985 N DEL 8
SRR1766475.9741166 chrX 532814 N chrX 532986 N DEL 8
SRR1766442.44552150 chrX 532816 N chrX 532988 N DEL 8
SRR1766481.8043450 chrX 532816 N chrX 532988 N DEL 8
SRR1766448.8015409 chrX 532822 N chrX 532994 N DEL 6
SRR1766478.10407683 chrX 532822 N chrX 532994 N DEL 6
SRR1766466.4858301 chrX 532823 N chrX 532995 N DEL 5
SRR1766466.741586 chrX 532827 N chrX 532999 N DEL 1
SRR1766482.5839177 chrX 532512 N chrX 533031 N DEL 5
SRR1766455.1920327 chrX 532698 N chrX 533041 N DEL 5
SRR1766453.6694744 chrX 532359 N chrX 533043 N DEL 8
SRR1766451.2428632 chrX 532814 N chrX 533157 N DEL 5
SRR1766467.11936841 chr7 4125032 N chr7 4125529 N DEL 5
SRR1766477.5930342 chr7 4125047 N chr7 4125493 N DEL 7
SRR1766471.4497294 chr7 4125056 N chr7 4125301 N DEL 14
SRR1766486.10138534 chr7 4125175 N chr7 4125538 N DEL 10
SRR1766478.3592999 chr7 4125081 N chr7 4125182 N DUP 5
SRR1766476.11171341 chr7 4125034 N chr7 4125265 N DUP 10
SRR1766484.573583 chr7 4125023 N chr7 4125157 N DEL 10
SRR1766477.10519006 chr7 4125174 N chr7 4125271 N DUP 5
SRR1766452.3954220 chr7 4125196 N chr7 4125407 N DUP 5
SRR1766483.11842484 chr7 4125054 N chr7 4125317 N DUP 1
SRR1766444.6082632 chr7 4125231 N chr7 4125686 N DUP 4
SRR1766457.1353461 chr7 4125054 N chr7 4125263 N DEL 6
SRR1766465.7784291 chr7 4125325 N chr7 4125398 N DUP 1
SRR1766470.2172997 chr7 4125061 N chr7 4125318 N DEL 5
SRR1766479.8338793 chr7 4125071 N chr7 4125367 N DEL 5
SRR1766457.4842981 chr7 4125082 N chr7 4125374 N DEL 5
SRR1766478.8662302 chr7 4125084 N chr7 4125376 N DEL 5
SRR1766469.8353976 chr7 4125057 N chr7 4125381 N DEL 6
SRR1766485.6945862 chr7 4125059 N chr7 4125493 N DEL 15
SRR1766482.518402 chr7 4125095 N chr7 4125501 N DEL 4
SRR1766442.7998604 chr7 4125058 N chr7 4125504 N DEL 4
SRR1766460.2223474 chr7 4125055 N chr7 4125497 N DEL 11
SRR1766463.444526 chr7 4125237 N chr7 4125565 N DEL 2
SRR1766481.9157094 chr7 4125069 N chr7 4125573 N DEL 5
SRR1766445.8578877 chr7 4125274 N chr7 4125606 N DEL 1
SRR1766470.7032325 chr7 4125051 N chr7 4125607 N DEL 3
SRR1766476.1873146 chr7 4125057 N chr7 4125653 N DEL 1
SRR1766486.6071078 chr11 39227958 N chr11 39228049 N DEL 2
SRR1766453.10211856 chr11 39227973 N chr11 39228088 N DEL 16
SRR1766469.10040682 chr11 39227973 N chr11 39228088 N DEL 17
SRR1766442.34386644 chr11 39228018 N chr11 39228077 N DUP 4
SRR1766467.4683945 chr11 39228020 N chr11 39228079 N DUP 2
SRR1766460.3845140 chr11 39227967 N chr11 39228042 N DEL 9
SRR1766468.5064553 chr11 39227967 N chr11 39228042 N DEL 9
SRR1766442.17931865 chr11 39227967 N chr11 39228042 N DEL 9
SRR1766453.10062123 chr11 39227967 N chr11 39228042 N DEL 9
SRR1766461.5969618 chr11 39227968 N chr11 39228043 N DEL 9
SRR1766442.14911280 chr11 39227969 N chr11 39228044 N DEL 9
SRR1766468.5333061 chr11 39227969 N chr11 39228044 N DEL 9
SRR1766450.1924135 chr11 39227970 N chr11 39228045 N DEL 9
SRR1766479.13238288 chr11 39227973 N chr11 39228048 N DEL 9
SRR1766469.2324673 chr11 39227976 N chr11 39228051 N DEL 6
SRR1766478.7916475 chr11 39227974 N chr11 39228049 N DEL 8
SRR1766470.4291055 chr3 197602823 N chr3 197602900 N DEL 5
SRR1766486.8261215 chr3 197602798 N chr3 197602874 N DUP 5
SRR1766465.9581788 chr3 197602679 N chr3 197602910 N DUP 5
SRR1766472.3283146 chr3 197602791 N chr3 197602908 N DEL 6
SRR1766467.8664836 chr3 83741640 N chr3 83741732 N DUP 2
SRR1766466.7695446 chr22 10851006 N chr22 10851403 N DEL 11
SRR1766470.7182439 chr22 10851067 N chr22 10851264 N DUP 5
SRR1766479.1788208 chr22 10851268 N chr22 10851468 N DEL 5
SRR1766470.5824672 chr22 10851268 N chr22 10851468 N DEL 5
SRR1766445.5127916 chr22 10851081 N chr22 10851280 N DEL 5
SRR1766453.10867409 chr22 10851284 N chr22 10851482 N DUP 4
SRR1766466.1283208 chr22 10850908 N chr22 10851503 N DUP 1
SRR1766457.8596287 chr22 10851006 N chr22 10851403 N DEL 11
SRR1766454.5562365 chr5 95927538 N chr5 95927687 N DEL 9
SRR1766462.9388745 chr5 95927538 N chr5 95927687 N DEL 9
SRR1766464.10795041 chr5 95927538 N chr5 95927687 N DEL 9
SRR1766448.8537627 chr5 95927538 N chr5 95927687 N DEL 11
SRR1766482.5734359 chr5 95927538 N chr5 95927687 N DEL 12
SRR1766453.4684209 chr5 95927538 N chr5 95927687 N DEL 13
SRR1766473.2657398 chr5 95927538 N chr5 95927687 N DEL 14
SRR1766448.1948502 chr5 95927538 N chr5 95927687 N DEL 18
SRR1766456.4332329 chr5 95927538 N chr5 95927687 N DEL 18
SRR1766484.7202850 chr5 95927538 N chr5 95927687 N DEL 18
SRR1766442.19374397 chr5 95927575 N chr5 95927626 N DEL 8
SRR1766453.9194829 chr5 95927538 N chr5 95927687 N DEL 18
SRR1766464.10687207 chr5 95927575 N chr5 95927626 N DEL 10
SRR1766474.1518101 chr5 95927534 N chr5 95927585 N DUP 3
SRR1766453.1566577 chr5 95927534 N chr5 95927585 N DUP 3
SRR1766450.3401078 chr5 95927602 N chr5 95927673 N DUP 14
SRR1766485.6700458 chr5 95927602 N chr5 95927673 N DUP 14
SRR1766450.907134 chr5 95927575 N chr5 95927626 N DEL 13
SRR1766442.2632727 chr5 95927575 N chr5 95927626 N DEL 9
SRR1766479.10926599 chr5 95927575 N chr5 95927626 N DEL 13
SRR1766447.4395770 chr5 95927575 N chr5 95927626 N DEL 9
SRR1766455.5298750 chr5 95927523 N chr5 95927628 N DEL 9
SRR1766442.22206083 chr5 95927525 N chr5 95927608 N DEL 7
SRR1766462.4474523 chr5 95927526 N chr5 95927609 N DEL 7
SRR1766453.4150939 chr5 95927526 N chr5 95927609 N DEL 7
SRR1766463.1469534 chr5 95927563 N chr5 95927616 N DEL 1
SRR1766451.1875257 chr5 95927575 N chr5 95927626 N DEL 9
SRR1766442.25678286 chr5 95927575 N chr5 95927626 N DEL 9
SRR1766485.3520738 chr5 95927528 N chr5 95927633 N DEL 8
SRR1766452.3337225 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766479.7592797 chr5 95927550 N chr5 95927601 N DUP 7
SRR1766446.494000 chr5 95927650 N chr5 95927777 N DUP 7
SRR1766450.10676330 chr5 95927650 N chr5 95927777 N DUP 7
SRR1766475.4472248 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766473.2140803 chr5 95927550 N chr5 95927601 N DUP 7
SRR1766448.3094478 chr5 95927550 N chr5 95927627 N DUP 4
SRR1766472.390523 chr5 95927538 N chr5 95927687 N DEL 17
SRR1766462.1362974 chr5 95927538 N chr5 95927687 N DEL 16
SRR1766442.20756671 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766479.12868825 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766450.8802746 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766459.8336509 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766480.8285736 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766447.8596740 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766462.9388745 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766449.3861440 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766464.10795041 chr5 95927625 N chr5 95927804 N DEL 7
SRR1766475.10572458 chr5 95927599 N chr5 95927804 N DEL 7
SRR1766485.2472895 chr5 95927599 N chr5 95927804 N DEL 7
SRR1766448.1948502 chr5 95927599 N chr5 95927804 N DEL 7
SRR1766449.8778324 chr5 95927599 N chr5 95927804 N DEL 7
SRR1766480.2514503 chr5 95927599 N chr5 95927804 N DEL 7
SRR1766474.9791763 chr5 95927599 N chr5 95927804 N DEL 7
SRR1766448.8537627 chr5 95927723 N chr5 95927856 N DEL 14
SRR1766442.17561281 chr5 95927723 N chr5 95927856 N DEL 14
SRR1766442.42413776 chr5 95927723 N chr5 95927856 N DEL 14
SRR1766453.9194829 chr5 95927723 N chr5 95927856 N DEL 14
SRR1766474.3141017 chr5 95927599 N chr5 95927856 N DEL 14
SRR1766447.2933504 chr5 95927599 N chr5 95927856 N DEL 13
SRR1766449.4709640 chr5 95927599 N chr5 95927856 N DEL 10
SRR1766460.5377270 chr5 95927599 N chr5 95927856 N DEL 7
SRR1766448.10558401 chr5 95927599 N chr5 95927856 N DEL 7
SRR1766447.192606 chr5 95927599 N chr5 95927856 N DEL 7
SRR1766474.6903853 chr5 95927599 N chr5 95927856 N DEL 7
SRR1766442.45687085 chr5 95927599 N chr5 95927856 N DEL 7
SRR1766485.1385375 chr5 95927599 N chr5 95927886 N DEL 10
SRR1766442.39842660 chr5 95927599 N chr5 95927886 N DEL 13
SRR1766482.8962914 chr5 95927599 N chr5 95927886 N DEL 15
SRR1766457.1080109 chr5 95927854 N chr5 95927941 N DUP 15
SRR1766451.6600763 chr5 95927573 N chr5 95927886 N DEL 10
SRR1766445.3112775 chr5 95927573 N chr5 95927886 N DEL 7
SRR1766462.4474523 chr5 95927573 N chr5 95927886 N DEL 7
SRR1766442.29748881 chr5 95927575 N chr5 95927888 N DEL 7
SRR1766466.2542705 chr5 95927575 N chr5 95927888 N DEL 7
SRR1766477.2458410 chr5 95927576 N chr5 95927889 N DEL 7
SRR1766442.5064651 chr13 27998900 N chr13 27999013 N DEL 1
SRR1766474.8435483 chr13 27998900 N chr13 27999013 N DEL 1
SRR1766477.4423267 chr13 27998916 N chr13 27998997 N DUP 4
SRR1766481.2901421 chr13 27998916 N chr13 27998997 N DUP 4
SRR1766480.2377444 chr13 27998890 N chr13 27999040 N DUP 6
SRR1766442.35315888 chr13 27998968 N chr13 27999019 N DUP 24
SRR1766475.4958283 chr13 27998968 N chr13 27999019 N DUP 25
SRR1766484.9177243 chr13 27998968 N chr13 27999019 N DUP 27
SRR1766449.7027146 chr13 27998968 N chr13 27999019 N DUP 28
SRR1766442.10168482 chr13 27998912 N chr13 27999042 N DUP 14
SRR1766472.11307815 chr13 27998968 N chr13 27999019 N DUP 30
SRR1766463.6908159 chr13 27998968 N chr13 27999019 N DUP 30
SRR1766483.6258830 chr13 27998983 N chr13 27999041 N DEL 21
SRR1766442.29273071 chr13 27998968 N chr13 27999019 N DUP 22
SRR1766452.1060388 chr13 27998964 N chr13 27999037 N DUP 19
SRR1766447.5182355 chr13 27998962 N chr13 27999066 N DUP 28
SRR1766477.5162579 chr13 27998968 N chr13 27999019 N DUP 26
SRR1766448.3961823 chr13 27998968 N chr13 27999019 N DUP 27
SRR1766481.1593684 chr13 27998968 N chr13 27999019 N DUP 30
SRR1766466.3304096 chr13 27998909 N chr13 27998968 N DEL 7
SRR1766464.3101435 chr13 27999088 N chr13 27999286 N DEL 11
SRR1766476.1476588 chr13 27998960 N chr13 27999064 N DUP 15
SRR1766486.2975113 chr13 27998960 N chr13 27999064 N DUP 18
SRR1766473.3760361 chr13 27998911 N chr13 27999024 N DEL 4
SRR1766486.6846917 chr13 27998987 N chr13 27999047 N DEL 2
SRR1766473.217054 chr13 27999047 N chr13 27999112 N DUP 14
SRR1766455.5249921 chr13 27999047 N chr13 27999112 N DUP 14
SRR1766449.1535673 chr13 27999107 N chr13 27999188 N DEL 6
SRR1766445.7825528 chr13 27998984 N chr13 27999042 N DEL 14
SRR1766453.780664 chr13 27998960 N chr13 27999064 N DUP 19
SRR1766463.10567222 chr13 27999013 N chr13 27999149 N DUP 26
SRR1766465.3351649 chr13 27999042 N chr13 27999107 N DUP 18
SRR1766476.9413642 chr13 27998982 N chr13 27999042 N DEL 7
SRR1766478.8560053 chr13 27998961 N chr13 27999171 N DUP 7
SRR1766453.2406926 chr13 27998967 N chr13 27999171 N DUP 17
SRR1766454.4206526 chr13 27998983 N chr13 27999041 N DEL 16
SRR1766485.427727 chr13 27998960 N chr13 27999174 N DUP 15
SRR1766462.2537060 chr13 27998964 N chr13 27999258 N DUP 19
SRR1766473.3699132 chr13 27999047 N chr13 27999112 N DUP 22
SRR1766452.7910045 chr13 27998967 N chr13 27999171 N DUP 23
SRR1766453.3680967 chr13 27998950 N chr13 27999150 N DUP 27
SRR1766486.6316215 chr13 27998961 N chr13 27999127 N DUP 18
SRR1766445.1502972 chr13 27999109 N chr13 27999172 N DEL 16
SRR1766475.9643434 chr13 27999109 N chr13 27999172 N DEL 15
SRR1766476.10462932 chr13 27999196 N chr13 27999260 N DUP 42
SRR1766482.8602446 chr13 27999093 N chr13 27999246 N DEL 15
SRR1766482.9737075 chr13 27999112 N chr13 27999286 N DEL 13
SRR1766448.6395271 chr13 27999093 N chr13 27999246 N DEL 16
SRR1766454.9377414 chr13 27998911 N chr13 27999235 N DEL 9
SRR1766472.9208603 chr13 27999093 N chr13 27999246 N DEL 16
SRR1766454.143376 chr13 27999305 N chr13 27999364 N DUP 8
SRR1766469.3160727 chr13 27999305 N chr13 27999364 N DUP 8
SRR1766485.5335596 chr13 27998911 N chr13 27999235 N DEL 9
SRR1766442.33258567 chr13 27999305 N chr13 27999364 N DUP 13
SRR1766470.6193709 chr13 27999305 N chr13 27999364 N DUP 27
SRR1766468.3392298 chr13 27999305 N chr13 27999364 N DUP 15
SRR1766448.10015345 chr13 27999125 N chr13 27999307 N DEL 5
SRR1766449.7959744 chr13 27999291 N chr13 27999368 N DEL 20
SRR1766448.2538942 chr13 27999298 N chr13 27999375 N DEL 8
SRR1766465.3351649 chr13 27999292 N chr13 27999369 N DEL 14
SRR1766485.2124696 chr13 27999291 N chr13 27999398 N DEL 5
SRR1766445.4562627 chr13 27999291 N chr13 27999398 N DEL 5
SRR1766450.4672932 chr13 27999292 N chr13 27999399 N DEL 5
SRR1766442.29233473 chr13 27999292 N chr13 27999399 N DEL 5
SRR1766470.9841752 chr8 141107273 N chr8 141107956 N DEL 5
SRR1766456.486476 chr8 141107319 N chr8 141107786 N DEL 5
SRR1766449.2341929 chr8 141107329 N chr8 141108064 N DEL 10
SRR1766480.4582855 chr8 141107330 N chr8 141107605 N DEL 4
SRR1766479.3837233 chr8 141107332 N chr8 141108067 N DEL 7
SRR1766475.1530968 chr8 141107330 N chr8 141107605 N DEL 5
SRR1766443.2124347 chr8 141107340 N chr8 141107615 N DEL 5
SRR1766466.3563887 chr8 141107366 N chr8 141107613 N DEL 10
SRR1766442.6644827 chr8 141107278 N chr8 141107387 N DUP 5
SRR1766475.2671557 chr8 141107386 N chr8 141107633 N DEL 5
SRR1766467.8858381 chr8 141107338 N chr8 141107777 N DEL 6
SRR1766475.5792338 chr8 141107429 N chr8 141108108 N DEL 7
SRR1766461.1907734 chr8 141107427 N chr8 141107890 N DEL 5
SRR1766467.6929163 chr8 141107496 N chr8 141107663 N DEL 6
SRR1766474.3954979 chr8 141107486 N chr8 141107541 N DEL 8
SRR1766442.22819411 chr8 141107280 N chr8 141107447 N DEL 3
SRR1766479.4036519 chr8 141107540 N chr8 141107949 N DEL 19
SRR1766443.1832361 chr8 141107405 N chr8 141107566 N DUP 2
SRR1766455.3537393 chr8 141107469 N chr8 141107794 N DUP 5
SRR1766479.9989100 chr8 141107566 N chr8 141107623 N DEL 1
SRR1766464.10959847 chr8 141107566 N chr8 141107623 N DEL 4
SRR1766479.503744 chr8 141107528 N chr8 141107801 N DUP 10
SRR1766443.2124347 chr8 141107451 N chr8 141107532 N DEL 8
SRR1766476.10924834 chr8 141107655 N chr8 141108116 N DEL 8
SRR1766462.4683611 chr8 141107467 N chr8 141107602 N DEL 10
SRR1766485.300084 chr8 141107639 N chr8 141107774 N DUP 17
SRR1766446.1661137 chr8 141107613 N chr8 141108074 N DUP 5
SRR1766480.1068179 chr8 141107450 N chr8 141107613 N DEL 5
SRR1766480.3151908 chr8 141107639 N chr8 141107828 N DUP 15
SRR1766456.1171620 chr8 141107639 N chr8 141107720 N DUP 8
SRR1766484.2206904 chr8 141107277 N chr8 141107634 N DEL 2
SRR1766445.3470910 chr8 141107553 N chr8 141107636 N DEL 2
SRR1766460.9761426 chr8 141107669 N chr8 141107776 N DUP 5
SRR1766461.1907734 chr8 141107723 N chr8 141107778 N DEL 5
SRR1766443.9061337 chr8 141107443 N chr8 141107690 N DEL 5
SRR1766442.38256591 chr8 141107683 N chr8 141107738 N DEL 5
SRR1766466.4814945 chr8 141107639 N chr8 141107774 N DUP 3
SRR1766453.9259003 chr8 141107639 N chr8 141107774 N DUP 17
SRR1766477.4812811 chr8 141107639 N chr8 141107774 N DUP 23
SRR1766451.8751495 chr8 141107435 N chr8 141107842 N DUP 4
SRR1766442.22819411 chr8 141107688 N chr8 141107743 N DEL 5
SRR1766475.5882689 chr8 141107745 N chr8 141107824 N DUP 6
SRR1766482.8536402 chr8 141107637 N chr8 141107776 N DEL 5
SRR1766475.10162709 chr8 141107550 N chr8 141107743 N DEL 5
SRR1766462.8497548 chr8 141107751 N chr8 141108074 N DUP 5
SRR1766463.2999767 chr8 141107637 N chr8 141107774 N DEL 10
SRR1766465.4474064 chr8 141107440 N chr8 141107955 N DUP 5
SRR1766474.4286031 chr8 141107604 N chr8 141107959 N DEL 5
SRR1766452.2832708 chr8 141107749 N chr8 141108046 N DEL 5
SRR1766474.3954979 chr8 141107749 N chr8 141108046 N DEL 5
SRR1766444.2055085 chr8 141107458 N chr8 141108055 N DEL 5
SRR1766467.8108957 chr8 141107426 N chr8 141108077 N DEL 5
SRR1766471.12193054 chr8 141107459 N chr8 141108110 N DEL 5
SRR1766465.2183344 chr14 94803992 N chr14 94804114 N DUP 12
SRR1766448.5616626 chr12 128205768 N chr12 128205899 N DUP 4
SRR1766472.3866853 chr12 128205761 N chr12 128205892 N DUP 5
SRR1766466.8204700 chr12 128205868 N chr12 128205975 N DUP 5
SRR1766449.10352324 chr12 128205803 N chr12 128205972 N DEL 5
SRR1766475.8341306 chr12 128205929 N chr12 128206001 N DEL 1
SRR1766454.1789467 chr12 128205899 N chr12 128206045 N DEL 5
SRR1766443.11202283 chr2 41747326 N chr2 41747782 N DEL 12
SRR1766467.3668075 chr2 41747361 N chr2 41747716 N DEL 6
SRR1766473.7426786 chr2 41747326 N chr2 41747782 N DEL 17
SRR1766457.3619805 chr2 41747377 N chr2 41747602 N DUP 8
SRR1766475.9833552 chr2 41747401 N chr2 41747610 N DUP 26
SRR1766443.6881291 chr2 41747407 N chr2 41747811 N DUP 9
SRR1766442.30575574 chr2 41747247 N chr2 41747376 N DEL 1
SRR1766442.38353285 chr2 41747240 N chr2 41747543 N DUP 5
SRR1766465.9079019 chr2 41747529 N chr2 41747708 N DEL 10
SRR1766476.2541200 chr2 41747243 N chr2 41747499 N DEL 5
SRR1766444.7066972 chr2 41747242 N chr2 41747547 N DEL 5
SRR1766471.1078284 chr2 41747607 N chr2 41747834 N DUP 8
SRR1766465.5318652 chr2 41747587 N chr2 41747816 N DUP 7
SRR1766467.4834416 chr2 41747387 N chr2 41747742 N DEL 4
SRR1766468.1525396 chr2 41747265 N chr2 41747977 N DEL 1
SRR1766443.11202283 chr2 41747651 N chr2 41747881 N DEL 5
SRR1766478.1213841 chr2 41747633 N chr2 41747990 N DEL 5
SRR1766443.3115765 chr2 41747852 N chr2 41748257 N DEL 1
SRR1766468.1525396 chr2 41747930 N chr2 41748257 N DEL 10
SRR1766480.3775410 chr10 478464 N chr10 478533 N DEL 9
SRR1766453.8571653 chr7 158404837 N chr7 158404986 N DEL 5
SRR1766473.6673531 chr7 158405128 N chr7 158405229 N DUP 3
SRR1766480.5092687 chr7 158404920 N chr7 158405141 N DEL 2
SRR1766480.2047595 chr7 158404960 N chr7 158405194 N DEL 5
SRR1766447.6175468 chr9 136849046 N chr9 136849144 N DEL 5
SRR1766463.9424319 chr5 79341638 N chr5 79341803 N DUP 5
SRR1766446.3448120 chr17 79555640 N chr17 79555759 N DUP 5
SRR1766453.5686119 chr17 79555643 N chr17 79555708 N DUP 10
SRR1766444.1074239 chr17 79555690 N chr17 79555779 N DUP 8
SRR1766468.1056974 chr17 79555761 N chr17 79555844 N DUP 10
SRR1766483.10739498 chr17 79555628 N chr17 79555761 N DEL 15
SRR1766462.5364184 chr17 79555761 N chr17 79556027 N DUP 9
SRR1766454.8108139 chr17 79555764 N chr17 79555847 N DUP 6
SRR1766473.10793314 chr17 79555762 N chr17 79555845 N DUP 5
SRR1766467.5260141 chr17 79555664 N chr17 79555761 N DEL 8
SRR1766464.10862645 chr17 79555668 N chr17 79555765 N DEL 5
SRR1766447.9384166 chr17 79555658 N chr17 79555773 N DEL 3
SRR1766454.8108139 chr17 79555630 N chr17 79555763 N DEL 8
SRR1766483.6638679 chr17 79555670 N chr17 79555803 N DEL 1
SRR1766442.26958715 chr17 79555669 N chr17 79555805 N DEL 2
SRR1766442.40057164 chr17 79555688 N chr17 79555836 N DEL 15
SRR1766471.6174033 chr17 79555627 N chr17 79555980 N DUP 3
SRR1766484.6121431 chr17 79555627 N chr17 79555980 N DUP 4
SRR1766459.1549019 chr17 79555669 N chr17 79555859 N DEL 5
SRR1766482.7277531 chr17 79555627 N chr17 79555980 N DUP 8
SRR1766442.23473056 chr17 79555848 N chr17 79555939 N DEL 11
SRR1766469.3835578 chr8 143711797 N chr8 143711906 N DEL 3
SRR1766443.5700751 chr11 9339959 N chr11 9340014 N DEL 2
SRR1766457.2029768 chr11 9339959 N chr11 9340014 N DEL 5
SRR1766457.8181538 chr11 9339959 N chr11 9340014 N DEL 5
SRR1766453.10712269 chr11 9339959 N chr11 9340014 N DEL 5
SRR1766461.4684254 chr11 9340001 N chr11 9340054 N DUP 5
SRR1766448.1141443 chr11 9340001 N chr11 9340054 N DUP 5
SRR1766463.10769524 chr11 9340003 N chr11 9340056 N DUP 5
SRR1766483.3846030 chr11 9340001 N chr11 9340054 N DUP 5
SRR1766447.1661809 chr11 9340001 N chr11 9340054 N DUP 5
SRR1766485.128906 chr11 9340001 N chr11 9340054 N DUP 5
SRR1766442.16186636 chr11 9340001 N chr11 9340054 N DUP 5
SRR1766486.18231 chr11 9340001 N chr11 9340054 N DUP 5
SRR1766458.8310233 chr11 9340005 N chr11 9340058 N DUP 5
SRR1766479.6792745 chr11 9340013 N chr11 9340066 N DUP 3
SRR1766482.945828 chr4 46977386 N chr4 46977480 N DEL 2
SRR1766473.1377218 chr22 44813415 N chr22 44813503 N DUP 5
SRR1766465.1771996 chr22 44813507 N chr22 44813579 N DEL 2
SRR1766455.3753854 chr22 44813507 N chr22 44813579 N DEL 4
SRR1766478.6765001 chr22 44813507 N chr22 44813579 N DEL 18
SRR1766466.518549 chr22 44813507 N chr22 44813579 N DEL 18
SRR1766442.2530365 chr22 44813507 N chr22 44813579 N DEL 18
SRR1766443.1886040 chr22 44813507 N chr22 44813579 N DEL 18
SRR1766453.4508940 chr22 44813408 N chr22 44813579 N DEL 16
SRR1766451.2645951 chr22 44813408 N chr22 44813579 N DEL 15
SRR1766463.6244956 chr22 44813514 N chr22 44813586 N DEL 8
SRR1766482.3296350 chr13 38036071 N chr13 38036346 N DUP 4
SRR1766471.9280067 chr16 22161740 N chr16 22161902 N DUP 1
SRR1766456.1721926 chr6 5035776 N chr6 5035912 N DEL 7
SRR1766461.58592 chr7 135096710 N chr7 135096898 N DEL 5
SRR1766481.10873199 chr7 135096709 N chr7 135096905 N DEL 2
SRR1766450.6818925 chr5 105934152 N chr5 105934279 N DUP 4
SRR1766462.2657546 chr5 105934178 N chr5 105934227 N DUP 1
SRR1766474.3387641 chr5 105934197 N chr5 105934254 N DEL 14
SRR1766479.1327134 chr5 105934197 N chr5 105934254 N DEL 14
SRR1766451.784357 chr5 105934197 N chr5 105934254 N DEL 13
SRR1766480.6446357 chr5 105934189 N chr5 105934254 N DEL 9
SRR1766455.533850 chr5 105934189 N chr5 105934254 N DEL 7
SRR1766442.8858546 chr5 105934189 N chr5 105934254 N DEL 7
SRR1766484.5750022 chr5 105934185 N chr5 105934254 N DEL 7
SRR1766442.10791018 chr5 105934181 N chr5 105934254 N DEL 7
SRR1766471.8097316 chr5 105934181 N chr5 105934254 N DEL 7
SRR1766468.1650417 chr5 105934177 N chr5 105934254 N DEL 7
SRR1766464.10917141 chr5 105934173 N chr5 105934254 N DEL 7
SRR1766456.5851116 chr5 105934173 N chr5 105934254 N DEL 7
SRR1766485.7888787 chr5 105934173 N chr5 105934254 N DEL 7
SRR1766468.1883784 chr5 105934169 N chr5 105934254 N DEL 7
SRR1766451.8174136 chr5 105934201 N chr5 105934254 N DEL 14
SRR1766460.6981384 chr5 105934212 N chr5 105934296 N DEL 6
SRR1766454.3530422 chr5 105934208 N chr5 105934296 N DEL 6
SRR1766464.10471731 chr5 105934196 N chr5 105934296 N DEL 6
SRR1766460.8063660 chr5 105934196 N chr5 105934296 N DEL 6
SRR1766445.4595235 chr5 105934192 N chr5 105934296 N DEL 6
SRR1766461.3075758 chr5 105934188 N chr5 105934296 N DEL 6
SRR1766461.7497638 chr5 105934184 N chr5 105934296 N DEL 6
SRR1766462.7177482 chr5 105934180 N chr5 105934296 N DEL 6
SRR1766446.7068426 chr5 105934153 N chr5 105934306 N DEL 1
SRR1766472.6919951 chr5 105934153 N chr5 105934306 N DEL 1
SRR1766455.9704275 chr5 105934155 N chr5 105934308 N DEL 3
SRR1766447.2796041 chr22 16311039 N chr22 16311090 N DUP 5
SRR1766471.10894678 chr22 16311144 N chr22 16311220 N DEL 10
SRR1766450.9270371 chr22 16311144 N chr22 16311220 N DEL 12
SRR1766452.719356 chr22 16311103 N chr22 16311154 N DUP 6
SRR1766443.6420772 chr22 16311144 N chr22 16311220 N DEL 5
SRR1766464.2099505 chr22 16311144 N chr22 16311220 N DEL 5
SRR1766447.6053161 chr22 16311103 N chr22 16311154 N DUP 4
SRR1766483.5637666 chr22 16311144 N chr22 16311220 N DEL 5
SRR1766466.1891627 chr22 16311144 N chr22 16311220 N DEL 5
SRR1766442.13274391 chr22 16311116 N chr22 16311216 N DUP 13
SRR1766442.38890689 chr22 16311028 N chr22 16311130 N DEL 10
SRR1766469.3650084 chr22 16311137 N chr22 16311237 N DUP 4
SRR1766468.4745036 chr19 2796463 N chr19 2796645 N DEL 4
SRR1766482.10859598 chr3 59012508 N chr3 59012647 N DEL 1
SRR1766462.2059369 chr5 76812173 N chr5 76812561 N DUP 1
SRR1766482.4511387 chr5 76812173 N chr5 76812561 N DUP 5
SRR1766456.557089 chr5 76812328 N chr5 76812562 N DEL 12
SRR1766471.10978943 chr5 76812197 N chr5 76812587 N DEL 5
SRR1766454.781516 chr5 76812200 N chr5 76812590 N DEL 2
SRR1766455.5593417 chr5 76812201 N chr5 76812591 N DEL 1
SRR1766451.2681979 chr5 76812641 N chr5 76812691 N DUP 4
SRR1766467.1209413 chr20 57090921 N chr20 57090991 N DEL 5
SRR1766453.3855985 chr20 57091054 N chr20 57091133 N DEL 5
SRR1766482.1075519 chr14 103896736 N chr14 103896870 N DEL 5
SRR1766480.7537691 chr14 103896736 N chr14 103896870 N DEL 12
SRR1766455.7545021 chr14 103896736 N chr14 103896870 N DEL 14
SRR1766456.3212529 chr14 103896736 N chr14 103896870 N DEL 14
SRR1766463.9267279 chr14 103896736 N chr14 103896870 N DEL 14
SRR1766460.651924 chr14 103896736 N chr14 103896870 N DEL 32
SRR1766462.8889482 chr14 103896737 N chr14 103896902 N DUP 27
SRR1766475.5539064 chr14 103896746 N chr14 103896911 N DUP 9
SRR1766442.18313176 chr14 103896746 N chr14 103896911 N DUP 9
SRR1766443.4492413 chr14 103896746 N chr14 103896911 N DUP 9
SRR1766464.3217137 chr14 103896748 N chr14 103896880 N DUP 4
SRR1766464.2306483 chr14 103896744 N chr14 103896909 N DUP 8
SRR1766475.8483473 chr14 103896777 N chr14 103896877 N DUP 10
SRR1766449.8307387 chr14 103896728 N chr14 103896793 N DEL 5
SRR1766477.11111545 chr17 32027468 N chr17 32027703 N DEL 12
SRR1766464.7045650 chr17 32027469 N chr17 32027546 N DEL 33
SRR1766442.35916864 chr17 32027530 N chr17 32027665 N DEL 3
SRR1766449.10273736 chr17 32027499 N chr17 32027692 N DUP 16
SRR1766465.8638326 chr17 32027521 N chr17 32027640 N DEL 5
SRR1766465.5382969 chr17 32027519 N chr17 32027654 N DEL 2
SRR1766479.11758575 chr17 32027516 N chr17 32027665 N DEL 10
SRR1766458.5469163 chr1 27086658 N chr1 27086808 N DUP 2
SRR1766485.5433374 chr1 27086658 N chr1 27086808 N DUP 2
SRR1766483.8941785 chr1 27086672 N chr1 27087071 N DUP 4
SRR1766450.8432816 chr1 27086689 N chr1 27086919 N DUP 4
SRR1766458.5217232 chr1 27086744 N chr1 27087193 N DUP 11
SRR1766455.1047524 chr1 27086877 N chr1 27087108 N DEL 2
SRR1766446.5051086 chr1 27086975 N chr1 27087122 N DEL 10
SRR1766480.6404983 chr1 27086808 N chr1 27086978 N DEL 6
SRR1766442.9779386 chr10 127016801 N chr10 127017074 N DEL 2
SRR1766444.4473200 chr10 127016806 N chr10 127016897 N DEL 6
SRR1766467.6479431 chr10 127016910 N chr10 127017019 N DUP 5
SRR1766481.2658246 chr10 127017056 N chr10 127017195 N DEL 13
SRR1766457.402049 chr10 127016934 N chr10 127017126 N DUP 7
SRR1766476.9554196 chr10 127016787 N chr10 127017192 N DUP 2
SRR1766458.7463648 chr10 127017024 N chr10 127017217 N DUP 10
SRR1766451.10080637 chr10 127017088 N chr10 127017199 N DEL 1
SRR1766448.3976412 chr10 127016971 N chr10 127017202 N DEL 5
SRR1766476.4687958 chr10 127016796 N chr10 127017333 N DUP 4
SRR1766444.4416943 chr10 127017065 N chr10 127017237 N DEL 1
SRR1766452.402351 chr10 127017289 N chr10 127017386 N DUP 7
SRR1766451.5955766 chr10 127017129 N chr10 127017424 N DUP 9
SRR1766480.4291630 chr10 127017132 N chr10 127017347 N DEL 27
SRR1766480.4291630 chr10 127017135 N chr10 127017350 N DEL 12
SRR1766454.3056840 chr10 127016938 N chr10 127017486 N DUP 9
SRR1766458.4727321 chr19 29128480 N chr19 29128598 N DUP 5
SRR1766485.2363443 chr19 29128717 N chr19 29128995 N DUP 4
SRR1766454.8868857 chr19 29128612 N chr19 29129084 N DUP 5
SRR1766471.9651396 chr19 29129186 N chr19 29129664 N DEL 5
SRR1766442.5450879 chr19 29129268 N chr19 29129743 N DEL 5
SRR1766453.5058560 chr19 29129283 N chr19 29129949 N DEL 5
SRR1766450.5059803 chr19 29129088 N chr19 29129209 N DEL 5
SRR1766480.4849262 chr19 29129281 N chr19 29129754 N DUP 5
SRR1766442.14534437 chr19 29128730 N chr19 29129802 N DUP 2
SRR1766479.3698653 chr13 21186896 N chr13 21187090 N DEL 5
SRR1766479.2419548 chr13 21186866 N chr13 21187098 N DUP 5
SRR1766465.5244032 chr13 21187006 N chr13 21187161 N DUP 10
SRR1766451.4877539 chr13 21186956 N chr13 21187111 N DUP 5
SRR1766464.6347688 chr13 21186961 N chr13 21187116 N DUP 13
SRR1766465.931454 chrX 532964 N chrX 533139 N DEL 1
SRR1766463.2937286 chrX 532963 N chrX 533138 N DEL 2
SRR1766481.5743445 chrX 532910 N chrX 533083 N DUP 15
SRR1766471.2101902 chrX 532942 N chrX 533117 N DEL 3
SRR1766479.7259905 chrX 532910 N chrX 533083 N DUP 15
SRR1766477.911756 chrX 532853 N chrX 533026 N DUP 5
SRR1766447.7195572 chrX 532963 N chrX 533138 N DEL 5
SRR1766485.7632539 chrX 532905 N chrX 533078 N DUP 20
SRR1766485.8417833 chrX 532880 N chrX 533053 N DUP 15
SRR1766448.8150322 chrX 532911 N chrX 533084 N DUP 14
SRR1766483.8662027 chrX 532911 N chrX 533084 N DUP 12
SRR1766455.8427191 chrX 532910 N chrX 533083 N DUP 10
SRR1766465.10786183 chrX 532905 N chrX 533078 N DUP 15
SRR1766447.4543671 chrX 532911 N chrX 533084 N DUP 10
SRR1766470.10694971 chrX 532964 N chrX 533139 N DEL 5
SRR1766477.3122202 chrX 532963 N chrX 533138 N DEL 5
SRR1766449.5255823 chrX 532905 N chrX 533078 N DUP 15
SRR1766481.6379179 chrX 532905 N chrX 533078 N DUP 15
SRR1766446.9583030 chrX 532832 N chrX 532981 N DUP 5
SRR1766449.6873246 chrX 532963 N chrX 533138 N DEL 5
SRR1766459.6091257 chrX 532880 N chrX 533053 N DUP 5
SRR1766483.2085544 chrX 532905 N chrX 533078 N DUP 10
SRR1766442.4712355 chrX 532880 N chrX 533053 N DUP 5
SRR1766442.45090361 chrX 532911 N chrX 533084 N DUP 15
SRR1766486.1970114 chrX 532911 N chrX 533084 N DUP 15
SRR1766463.5423529 chrX 532910 N chrX 533083 N DUP 15
SRR1766459.5797587 chrX 532911 N chrX 533084 N DUP 10
SRR1766452.2924394 chrX 532911 N chrX 533084 N DUP 10
SRR1766449.8737437 chrX 532832 N chrX 533002 N DUP 11
SRR1766455.7942497 chrX 532832 N chrX 533002 N DUP 11
SRR1766459.5079220 chrX 532832 N chrX 533002 N DUP 13
SRR1766471.11981734 chrX 532832 N chrX 533005 N DUP 9
SRR1766484.10425771 chrX 532832 N chrX 533002 N DUP 18
SRR1766442.45639657 chrX 532911 N chrX 533084 N DUP 10
SRR1766460.2188702 chrX 532832 N chrX 533002 N DUP 18
SRR1766461.6522231 chrX 532911 N chrX 533084 N DUP 10
SRR1766470.6796442 chrX 532911 N chrX 533084 N DUP 10
SRR1766464.10919875 chrX 532913 N chrX 533086 N DUP 7
SRR1766477.11445418 chrX 532846 N chrX 533001 N DUP 33
SRR1766481.7843412 chrX 532846 N chrX 533001 N DUP 33
SRR1766448.4524579 chrX 532832 N chrX 533005 N DUP 15
SRR1766457.2827369 chrX 532832 N chrX 533002 N DUP 23
SRR1766481.10632956 chrX 532846 N chrX 533001 N DUP 32
SRR1766454.3179782 chrX 532832 N chrX 533005 N DUP 15
SRR1766477.11106464 chrX 532832 N chrX 533005 N DUP 25
SRR1766462.4664999 chrX 532832 N chrX 533005 N DUP 25
SRR1766443.5911404 chrX 532832 N chrX 533005 N DUP 25
SRR1766447.4543671 chrX 532911 N chrX 533084 N DUP 8
SRR1766451.4329360 chrX 532911 N chrX 533084 N DUP 8
SRR1766470.10057164 chr2 605326 N chr2 605399 N DUP 1
SRR1766475.10489133 chr2 605329 N chr2 605558 N DUP 10
SRR1766469.3246983 chr2 605280 N chr2 605333 N DEL 5
SRR1766465.9930226 chr2 605283 N chr2 605336 N DEL 5
SRR1766478.1592908 chr2 605283 N chr2 605336 N DEL 5
SRR1766474.10381981 chr2 605285 N chr2 605338 N DEL 3
SRR1766478.837368 chr2 605430 N chr2 605480 N DUP 5
SRR1766448.920701 chr2 605430 N chr2 605480 N DUP 5
SRR1766462.10637781 chr2 605271 N chr2 605480 N DEL 5
SRR1766449.10429990 chr3 160593979 N chr3 160594077 N DUP 3
SRR1766459.833798 chr3 160593979 N chr3 160594077 N DUP 5
SRR1766456.6339988 chr3 160593979 N chr3 160594077 N DUP 5
SRR1766459.6363408 chr3 160593979 N chr3 160594077 N DUP 5
SRR1766476.3010283 chr3 160593979 N chr3 160594077 N DUP 5
SRR1766474.7275166 chr3 160593979 N chr3 160594077 N DUP 5
SRR1766466.3646592 chr3 160593979 N chr3 160594077 N DUP 5
SRR1766476.6345955 chrX 140724592 N chrX 140724650 N DUP 17
SRR1766451.2489842 chrX 140724592 N chrX 140724656 N DUP 15
SRR1766465.1961337 chrX 140724651 N chrX 140724715 N DUP 5
SRR1766483.4138432 chr3 96621696 N chr3 96621774 N DEL 9
SRR1766464.711321 chr15 66130824 N chr15 66130895 N DUP 2
SRR1766455.962946 chr15 66130825 N chr15 66130896 N DUP 1
SRR1766456.2899665 chr10 132335404 N chr10 132335501 N DEL 5
SRR1766454.3443467 chr10 132335439 N chr10 132335536 N DEL 10
SRR1766462.1476549 chr10 132335460 N chr10 132335657 N DEL 26
SRR1766470.3114172 chr10 132335452 N chr10 132335547 N DUP 3
SRR1766449.6932787 chr10 132335461 N chr10 132335556 N DUP 5
SRR1766475.2115389 chr10 132335405 N chr10 132335596 N DUP 10
SRR1766471.3368258 chr10 132335405 N chr10 132335696 N DUP 5
SRR1766442.45456188 chr10 132335405 N chr10 132335696 N DUP 5
SRR1766450.607182 chr10 132335582 N chr10 132335782 N DEL 20
SRR1766445.3074113 chr1 193588247 N chr1 193588304 N DEL 1
SRR1766458.1795229 chr1 193588247 N chr1 193588304 N DEL 5
SRR1766445.1395671 chr1 193588247 N chr1 193588304 N DEL 6
SRR1766443.3564480 chr1 193588279 N chr1 193588366 N DUP 20
SRR1766453.1152432 chr1 193588279 N chr1 193588366 N DUP 25
SRR1766470.610446 chr1 193588279 N chr1 193588366 N DUP 20
SRR1766460.8957935 chr7 148365872 N chr7 148365999 N DUP 6
SRR1766485.10450576 chr7 148365899 N chr7 148366052 N DUP 4
SRR1766456.5030743 chr7 148365899 N chr7 148366052 N DUP 4
SRR1766444.7366380 chr7 148365899 N chr7 148366052 N DUP 5
SRR1766442.31600632 chr6 31068210 N chr6 31068287 N DEL 5
SRR1766447.9716661 chr6 31068343 N chr6 31068407 N DEL 14
SRR1766474.7883228 chr6 31068350 N chr6 31068414 N DEL 8
SRR1766452.10522602 chr6 31068379 N chr6 31068442 N DEL 5
SRR1766478.371039 chr4 103834851 N chr4 103835167 N DEL 3
SRR1766444.2088856 chr5 154652435 N chr5 154652756 N DEL 17
SRR1766444.3071076 chr5 154652441 N chr5 154652762 N DEL 9
SRR1766465.9233155 chr6 112528600 N chr6 112528834 N DEL 10
SRR1766486.1736144 chr6 112528624 N chr6 112528855 N DEL 3
SRR1766442.5732660 chr22 31355209 N chr22 31355513 N DEL 1
SRR1766483.11730131 chr1 68898314 N chr1 68898456 N DEL 7
SRR1766462.8294406 chr1 68898315 N chr1 68898457 N DEL 7
SRR1766453.9648669 chr1 68898316 N chr1 68898458 N DEL 7
SRR1766444.1016580 chr19 32954938 N chr19 32955259 N DEL 24
SRR1766457.2611892 chr19 32954935 N chr19 32955256 N DEL 5
SRR1766482.9998207 chr16 46382023 N chr16 46382152 N DUP 5
SRR1766469.731876 chr16 46382024 N chr16 46382153 N DUP 5
SRR1766463.5700014 chr16 46382025 N chr16 46382154 N DUP 5
SRR1766465.9882331 chr16 46382025 N chr16 46382154 N DUP 5
SRR1766475.935907 chr16 46382002 N chr16 46382196 N DUP 11
SRR1766450.5351797 chr16 46382002 N chr16 46382222 N DUP 11
SRR1766445.10481479 chr16 46382002 N chr16 46382222 N DUP 12
SRR1766469.7048807 chr16 46382002 N chr16 46382222 N DUP 13
SRR1766463.2338987 chr16 46382130 N chr16 46382207 N DUP 14
SRR1766480.2133975 chr16 46382002 N chr16 46382232 N DUP 3
SRR1766485.11056827 chr16 46382002 N chr16 46382232 N DUP 4
SRR1766448.6396761 chr16 46382002 N chr16 46382232 N DUP 4
SRR1766473.8515477 chr16 46382113 N chr16 46382291 N DUP 7
SRR1766472.5988805 chr16 46382002 N chr16 46382232 N DUP 5
SRR1766471.2773015 chr8 1368328 N chr8 1368544 N DEL 5
SRR1766472.620186 chr22 32564693 N chr22 32564789 N DEL 1
SRR1766469.568040 chr22 32564730 N chr22 32564967 N DEL 3
SRR1766473.3886724 chr22 32564775 N chr22 32565132 N DEL 3
SRR1766477.1060338 chr22 32564720 N chr22 32564815 N DUP 5
SRR1766448.4433470 chr22 32564820 N chr22 32565321 N DEL 5
SRR1766462.6431756 chr22 32564820 N chr22 32565321 N DEL 5
SRR1766460.2705199 chr22 32564795 N chr22 32565128 N DEL 14
SRR1766482.7946696 chr22 32564795 N chr22 32565104 N DEL 15
SRR1766486.7994384 chr22 32564820 N chr22 32565321 N DEL 5
SRR1766459.11473252 chr22 32564855 N chr22 32565020 N DEL 5
SRR1766452.7683969 chr22 32565007 N chr22 32565128 N DEL 22
SRR1766483.1025822 chr22 32564725 N chr22 32565032 N DUP 10
SRR1766451.9147954 chr22 32565043 N chr22 32565140 N DEL 18
SRR1766448.9008747 chr22 32564843 N chr22 32565054 N DUP 10
SRR1766447.9579897 chr22 32565061 N chr22 32565134 N DEL 4
SRR1766459.323124 chr22 32565060 N chr22 32565179 N DUP 5
SRR1766442.22811814 chr22 32565026 N chr22 32565193 N DUP 15
SRR1766475.5344120 chr22 32564858 N chr22 32564999 N DEL 5
SRR1766448.660446 chr22 32564692 N chr22 32565000 N DEL 5
SRR1766468.5860496 chr22 32564743 N chr22 32565004 N DEL 1
SRR1766473.10817027 chr22 32565161 N chr22 32565306 N DEL 4
SRR1766459.11473252 chr22 32564880 N chr22 32565045 N DEL 5
SRR1766479.6453026 chr22 32565154 N chr22 32565299 N DEL 8
SRR1766447.6659521 chr22 32565178 N chr22 32565299 N DEL 10
SRR1766443.3463904 chr22 32565178 N chr22 32565299 N DEL 10
SRR1766463.3201162 chr22 32564840 N chr22 32565195 N DUP 10
SRR1766447.9579897 chr22 32564854 N chr22 32565211 N DEL 5
SRR1766469.568040 chr22 32565188 N chr22 32565261 N DEL 5
SRR1766462.6431756 chr22 32565188 N chr22 32565261 N DEL 10
SRR1766465.5754144 chr22 32564823 N chr22 32565228 N DEL 5
SRR1766477.1060338 chr22 32564829 N chr22 32565234 N DEL 15
SRR1766452.7683969 chr22 32564880 N chr22 32565261 N DEL 8
SRR1766468.1247888 chr22 32564880 N chr22 32565261 N DEL 5
SRR1766473.3886724 chr22 32564880 N chr22 32565261 N DEL 5
SRR1766443.9126532 chr22 32565175 N chr22 32565296 N DEL 5
SRR1766442.34022770 chr22 32564747 N chr22 32565296 N DEL 5
SRR1766442.20815922 chr22 32564750 N chr22 32565299 N DEL 10
SRR1766473.8466007 chr22 32564958 N chr22 32565319 N DEL 5
SRR1766479.4114818 chr22 32564958 N chr22 32565319 N DEL 5
SRR1766478.1996432 chr22 32565179 N chr22 32565324 N DEL 3
SRR1766482.1704254 chr22 32564746 N chr22 32565319 N DEL 5
SRR1766442.35126576 chr22 32565019 N chr22 32565332 N DEL 10
SRR1766446.4746328 chr15 95761094 N chr15 95761148 N DUP 5
SRR1766477.11109204 chr5 120331265 N chr5 120331571 N DEL 10
SRR1766447.5881935 chr5 120331263 N chr5 120331571 N DEL 17
SRR1766448.8231890 chr5 120331265 N chr5 120331571 N DEL 13
SRR1766466.8467543 chr5 120331265 N chr5 120331571 N DEL 14
SRR1766446.1600829 chr5 120331266 N chr5 120331571 N DEL 15
SRR1766468.3080200 chr5 120331267 N chr5 120331571 N DEL 15
SRR1766485.9066541 chr22 31018597 N chr22 31018760 N DEL 3
SRR1766466.8113798 chr22 31018597 N chr22 31018760 N DEL 5
SRR1766483.7684297 chr22 31018598 N chr22 31018647 N DUP 10
SRR1766471.2434897 chr22 31018617 N chr22 31018830 N DUP 8
SRR1766478.10808845 chr22 31018615 N chr22 31018770 N DUP 10
SRR1766474.8443907 chr22 31018616 N chr22 31018829 N DUP 9
SRR1766459.7504193 chr22 31018660 N chr22 31018735 N DEL 6
SRR1766449.8725714 chr22 31018771 N chr22 31018830 N DEL 7
SRR1766443.7852719 chr22 31018660 N chr22 31018831 N DEL 5
SRR1766443.2655468 chr8 144513892 N chr8 144513946 N DEL 5
SRR1766450.6266288 chr8 144513900 N chr8 144513984 N DEL 10
SRR1766466.632635 chr8 144513900 N chr8 144513984 N DEL 11
SRR1766471.2806676 chr8 144513878 N chr8 144513960 N DUP 10
SRR1766470.9687831 chr8 144513945 N chr8 144514004 N DUP 24
SRR1766475.1370340 chr8 144513942 N chr8 144514031 N DUP 9
SRR1766466.9869156 chr8 144513883 N chr8 144513997 N DEL 9
SRR1766479.12350631 chr4 20084257 N chr4 20084401 N DUP 5
SRR1766479.897308 chr4 20084257 N chr4 20084401 N DUP 5
SRR1766444.2011287 chr4 20084508 N chr4 20084587 N DEL 2
SRR1766442.28463641 chr4 20084508 N chr4 20084587 N DEL 5
SRR1766446.5357297 chr4 20084508 N chr4 20084587 N DEL 7
SRR1766465.8939860 chr4 20084508 N chr4 20084587 N DEL 7
SRR1766453.942433 chr4 20084508 N chr4 20084587 N DEL 7
SRR1766446.9664949 chr4 20084508 N chr4 20084587 N DEL 7
SRR1766485.6732823 chr4 20084508 N chr4 20084587 N DEL 9
SRR1766455.3617250 chr4 20084508 N chr4 20084587 N DEL 10
SRR1766483.11307263 chr4 20084522 N chr4 20084601 N DEL 1
SRR1766454.4390265 chr4 20084521 N chr4 20084600 N DEL 2
SRR1766447.990765 chr4 20084529 N chr4 20084606 N DEL 9
SRR1766481.1040560 chr4 20084529 N chr4 20084606 N DEL 9
SRR1766475.11357017 chr4 20084529 N chr4 20084606 N DEL 9
SRR1766465.212443 chr4 20084537 N chr4 20084614 N DEL 7
SRR1766486.8742558 chr4 20084563 N chr4 20084640 N DEL 5
SRR1766477.6910360 chr4 20084563 N chr4 20084640 N DEL 5
SRR1766478.8515853 chr4 20084563 N chr4 20084640 N DEL 5
SRR1766461.9308606 chr4 20084525 N chr4 20084641 N DEL 5
SRR1766447.5103744 chr4 20084290 N chr4 20084664 N DEL 5
SRR1766442.26788231 chr4 20084291 N chr4 20084665 N DEL 5
SRR1766475.9307999 chr4 20084394 N chr4 20084666 N DEL 5
SRR1766483.3626812 chr16 30492415 N chr16 30492723 N DEL 2
SRR1766448.4405401 chr16 30492452 N chr16 30492759 N DEL 2
SRR1766473.8911220 chr16 30492454 N chr16 30492761 N DEL 5
SRR1766443.9818036 chr16 30492485 N chr16 30492792 N DEL 5
SRR1766442.16562425 chr20 29231810 N chr20 29232154 N DEL 6
SRR1766465.6274804 chr20 29232237 N chr20 29232577 N DUP 4
SRR1766465.7761975 chr20 29231754 N chr20 29232439 N DEL 15
SRR1766475.4809720 chr20 29231843 N chr20 29232526 N DUP 2
SRR1766469.8350954 chr3 129069510 N chr3 129069653 N DUP 2
SRR1766442.36751983 chr21 46691914 N chr21 46692194 N DEL 5
SRR1766447.4460022 chr21 46691879 N chr21 46692345 N DEL 15
SRR1766453.1649804 chr21 46691940 N chr21 46692683 N DEL 5
SRR1766475.4159702 chr21 46691914 N chr21 46692194 N DEL 5
SRR1766466.10818050 chr21 46691879 N chr21 46692345 N DEL 5
SRR1766472.1887632 chr21 46691939 N chr21 46692312 N DEL 5
SRR1766475.3495715 chr21 46691940 N chr21 46692313 N DEL 1
SRR1766452.10067194 chr21 46691914 N chr21 46692194 N DEL 5
SRR1766442.28599789 chr21 46691939 N chr21 46692589 N DEL 5
SRR1766481.4880136 chr21 46691914 N chr21 46692194 N DEL 5
SRR1766475.4756982 chr21 46691914 N chr21 46692194 N DEL 5
SRR1766452.5364863 chr21 46691862 N chr21 46692069 N DUP 11
SRR1766467.11783074 chr21 46691940 N chr21 46692313 N DEL 5
SRR1766467.570523 chr21 46691924 N chr21 46692297 N DEL 5
SRR1766462.6401292 chr21 46691923 N chr21 46692664 N DUP 5
SRR1766444.723462 chr21 46691924 N chr21 46692204 N DEL 6
SRR1766445.8958413 chr21 46691924 N chr21 46692204 N DEL 8
SRR1766478.2331386 chr21 46692016 N chr21 46692573 N DEL 5
SRR1766454.6505443 chr21 46692016 N chr21 46692573 N DEL 5
SRR1766461.157720 chr21 46692021 N chr21 46692115 N DEL 5
SRR1766442.39925528 chr21 46692021 N chr21 46692115 N DEL 5
SRR1766477.2349635 chr21 46691947 N chr21 46692039 N DUP 5
SRR1766442.18938873 chr21 46691947 N chr21 46692039 N DUP 5
SRR1766442.42054103 chr21 46691947 N chr21 46692039 N DUP 5
SRR1766463.9531752 chr21 46692033 N chr21 46692311 N DUP 5
SRR1766458.8737904 chr21 46692021 N chr21 46692115 N DEL 5
SRR1766442.42729999 chr21 46692033 N chr21 46692311 N DUP 5
SRR1766443.3943619 chr21 46691974 N chr21 46692345 N DUP 5
SRR1766451.6282302 chr21 46691947 N chr21 46692039 N DUP 5
SRR1766442.8486511 chr21 46691947 N chr21 46692039 N DUP 5
SRR1766482.5170815 chr21 46691947 N chr21 46692039 N DUP 5
SRR1766462.5033484 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766442.27976247 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766449.5717455 chr21 46691947 N chr21 46692039 N DUP 8
SRR1766465.2581381 chr21 46691973 N chr21 46692065 N DUP 4
SRR1766442.47148570 chr21 46691947 N chr21 46692039 N DUP 11
SRR1766451.7194082 chr21 46692114 N chr21 46692301 N DEL 5
SRR1766473.2960419 chr21 46692061 N chr21 46692343 N DEL 7
SRR1766442.3746511 chr21 46691947 N chr21 46692132 N DUP 5
SRR1766464.2573548 chr21 46692044 N chr21 46692506 N DUP 5
SRR1766448.2550757 chr21 46692125 N chr21 46692589 N DEL 10
SRR1766485.5883544 chr21 46692114 N chr21 46692301 N DEL 5
SRR1766454.3167232 chr21 46691995 N chr21 46692090 N DEL 15
SRR1766482.8541410 chr21 46691947 N chr21 46692132 N DUP 5
SRR1766442.22852177 chr21 46692125 N chr21 46692589 N DEL 10
SRR1766464.5766953 chr21 46692159 N chr21 46692530 N DEL 5
SRR1766478.3153880 chr21 46692132 N chr21 46692319 N DEL 5
SRR1766464.9451647 chr21 46691894 N chr21 46692081 N DEL 1
SRR1766458.5689457 chr21 46692159 N chr21 46692530 N DEL 13
SRR1766460.7883951 chr21 46692115 N chr21 46692207 N DUP 10
SRR1766486.2401640 chr21 46692021 N chr21 46692115 N DEL 5
SRR1766474.10768803 chr21 46692132 N chr21 46692319 N DEL 5
SRR1766481.2320907 chr21 46692021 N chr21 46692115 N DEL 5
SRR1766481.6236072 chr21 46692021 N chr21 46692115 N DEL 5
SRR1766483.1149532 chr21 46692159 N chr21 46692623 N DEL 10
SRR1766450.4572773 chr21 46692129 N chr21 46692314 N DUP 1
SRR1766479.10789831 chr21 46692218 N chr21 46692589 N DEL 5
SRR1766444.3635163 chr21 46691973 N chr21 46692160 N DEL 5
SRR1766454.7716912 chr21 46692193 N chr21 46692287 N DEL 5
SRR1766471.11965796 chr21 46691960 N chr21 46692147 N DEL 1
SRR1766452.3403749 chr21 46691973 N chr21 46692160 N DEL 5
SRR1766451.904271 chr21 46692193 N chr21 46692287 N DEL 5
SRR1766452.5034067 chr21 46692163 N chr21 46692255 N DUP 1
SRR1766442.20254511 chr21 46692414 N chr21 46692506 N DEL 8
SRR1766486.4534790 chr21 46692228 N chr21 46692506 N DEL 4
SRR1766454.3140822 chr21 46692219 N chr21 46692590 N DEL 10
SRR1766454.1534689 chr21 46691940 N chr21 46692404 N DUP 10
SRR1766449.1990844 chr21 46691892 N chr21 46692172 N DEL 2
SRR1766476.5643943 chr21 46692228 N chr21 46692506 N DEL 9
SRR1766465.10589477 chr21 46692295 N chr21 46692573 N DEL 5
SRR1766442.26888038 chr21 46692228 N chr21 46692506 N DEL 10
SRR1766478.10342993 chr21 46691914 N chr21 46692194 N DEL 5
SRR1766451.2021055 chr21 46692228 N chr21 46692506 N DEL 10
SRR1766453.9792203 chr21 46691924 N chr21 46692204 N DEL 10
SRR1766453.1618882 chr21 46691944 N chr21 46692036 N DUP 5
SRR1766482.6705002 chr21 46692219 N chr21 46692590 N DEL 15
SRR1766478.2309426 chr21 46691923 N chr21 46692203 N DEL 5
SRR1766450.990571 chr21 46692228 N chr21 46692506 N DEL 10
SRR1766463.1160325 chr21 46692219 N chr21 46692313 N DEL 5
SRR1766460.4193916 chr21 46691944 N chr21 46692224 N DEL 5
SRR1766482.704237 chr21 46691949 N chr21 46692506 N DEL 5
SRR1766445.7257402 chr21 46692222 N chr21 46692684 N DUP 12
SRR1766474.9280975 chr21 46692039 N chr21 46692226 N DEL 15
SRR1766478.467534 chr21 46692311 N chr21 46692589 N DEL 5
SRR1766473.318038 chr21 46692311 N chr21 46692589 N DEL 5
SRR1766452.6947660 chr21 46692311 N chr21 46692589 N DEL 5
SRR1766484.9650494 chr21 46692256 N chr21 46692348 N DUP 5
SRR1766478.4111649 chr21 46692133 N chr21 46692318 N DUP 2
SRR1766454.5778624 chr21 46692065 N chr21 46692252 N DEL 5
SRR1766461.2389548 chr21 46692133 N chr21 46692318 N DUP 5
SRR1766471.4277039 chr21 46692159 N chr21 46692253 N DEL 5
SRR1766455.6462125 chr21 46691947 N chr21 46692132 N DUP 10
SRR1766481.1223679 chr21 46692133 N chr21 46692318 N DUP 5
SRR1766442.20678799 chr21 46692345 N chr21 46692530 N DEL 2
SRR1766478.2322463 chr21 46692133 N chr21 46692318 N DUP 5
SRR1766472.3554045 chr21 46692133 N chr21 46692318 N DUP 5
SRR1766442.6529872 chr21 46692321 N chr21 46692506 N DEL 10
SRR1766444.3635163 chr21 46692133 N chr21 46692318 N DUP 5
SRR1766483.1653048 chr21 46692013 N chr21 46692384 N DUP 1
SRR1766467.9976925 chr21 46692013 N chr21 46692384 N DUP 4
SRR1766482.3990530 chr21 46692345 N chr21 46692530 N DEL 10
SRR1766445.8958413 chr21 46692033 N chr21 46692220 N DEL 10
SRR1766459.1494706 chr21 46692387 N chr21 46692665 N DEL 5
SRR1766442.4205767 chr21 46692478 N chr21 46692665 N DEL 11
SRR1766476.1413096 chr21 46692198 N chr21 46692292 N DEL 5
SRR1766446.8526451 chr21 46692254 N chr21 46692344 N DUP 7
SRR1766450.3549229 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766476.7331748 chr21 46692388 N chr21 46692573 N DEL 5
SRR1766477.5796702 chr21 46692392 N chr21 46692577 N DEL 5
SRR1766476.8716028 chr21 46692345 N chr21 46692530 N DEL 11
SRR1766470.3399220 chr21 46692032 N chr21 46692312 N DEL 5
SRR1766453.1949814 chr21 46692039 N chr21 46692319 N DEL 5
SRR1766443.7091697 chr21 46692157 N chr21 46692433 N DUP 5
SRR1766473.5530273 chr21 46692344 N chr21 46692438 N DEL 5
SRR1766442.42054103 chr21 46692350 N chr21 46692442 N DEL 4
SRR1766446.5968838 chr21 46691947 N chr21 46692502 N DUP 5
SRR1766462.4393885 chr21 46692014 N chr21 46692476 N DUP 5
SRR1766466.10355654 chr21 46692505 N chr21 46692599 N DEL 4
SRR1766461.8926206 chr21 46691977 N chr21 46692441 N DEL 9
SRR1766459.1775662 chr21 46692164 N chr21 46692442 N DEL 7
SRR1766481.7412759 chr21 46692169 N chr21 46692447 N DEL 2
SRR1766481.539788 chr21 46691982 N chr21 46692446 N DEL 6
SRR1766470.7895946 chr21 46691982 N chr21 46692446 N DEL 6
SRR1766465.302334 chr21 46691986 N chr21 46692450 N DEL 2
SRR1766446.10311746 chr21 46692025 N chr21 46692489 N DEL 11
SRR1766481.668459 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766442.19772023 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766442.39925528 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766457.2652553 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766476.10135851 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766481.10875142 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766485.6998333 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766478.2331386 chr21 46691914 N chr21 46692471 N DEL 5
SRR1766442.3612491 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766481.231902 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766445.9763279 chr21 46692025 N chr21 46692489 N DEL 10
SRR1766453.1618882 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766455.7853259 chr21 46692211 N chr21 46692489 N DEL 5
SRR1766464.2499478 chr21 46692025 N chr21 46692489 N DEL 9
SRR1766465.5044106 chr21 46692025 N chr21 46692489 N DEL 5
SRR1766457.1577120 chr21 46692025 N chr21 46692489 N DEL 5
SRR1766444.6266353 chr21 46692025 N chr21 46692489 N DEL 5
SRR1766458.7058430 chr21 46692318 N chr21 46692503 N DEL 15
SRR1766456.5327254 chr21 46692028 N chr21 46692492 N DEL 5
SRR1766472.11358348 chr21 46692032 N chr21 46692496 N DEL 5
SRR1766457.7823847 chr21 46692032 N chr21 46692496 N DEL 5
SRR1766467.7358080 chr21 46692572 N chr21 46692666 N DEL 3
SRR1766451.198811 chr21 46692036 N chr21 46692500 N DEL 4
SRR1766466.9201840 chr21 46692038 N chr21 46692502 N DEL 2
SRR1766451.6282302 chr21 46692046 N chr21 46692510 N DEL 5
SRR1766461.2051635 chr21 46692048 N chr21 46692512 N DEL 5
SRR1766446.7447435 chr21 46692050 N chr21 46692514 N DEL 5
SRR1766474.9280975 chr21 46692053 N chr21 46692517 N DEL 4
SRR1766479.6234112 chr21 46692053 N chr21 46692517 N DEL 4
SRR1766448.2550757 chr21 46691961 N chr21 46692518 N DEL 3
SRR1766462.673356 chr21 46691962 N chr21 46692519 N DEL 2
SRR1766446.5267120 chr21 46692388 N chr21 46692573 N DEL 11
SRR1766473.3935525 chr21 46692579 N chr21 46692671 N DUP 12
SRR1766455.9580449 chr21 46692016 N chr21 46692573 N DEL 5
SRR1766463.5783961 chr21 46692572 N chr21 46692664 N DUP 6
SRR1766465.5359671 chr21 46691960 N chr21 46692517 N DEL 4
SRR1766471.7927364 chr21 46691960 N chr21 46692517 N DEL 4
SRR1766452.7854478 chr21 46692572 N chr21 46692664 N DUP 5
SRR1766446.7097061 chr21 46692016 N chr21 46692573 N DEL 5
SRR1766473.5291074 chr21 46692016 N chr21 46692573 N DEL 5
SRR1766481.6236072 chr21 46692016 N chr21 46692573 N DEL 5
SRR1766479.2824430 chr21 46692016 N chr21 46692573 N DEL 5
SRR1766478.630594 chr21 46692312 N chr21 46692588 N DUP 5
SRR1766446.6766721 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766464.9797292 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766478.10872389 chr21 46692572 N chr21 46692664 N DUP 5
SRR1766449.8392860 chr21 46692503 N chr21 46692595 N DUP 12
SRR1766460.10115496 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766459.4255384 chr21 46692016 N chr21 46692573 N DEL 5
SRR1766466.10355654 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766478.8232437 chr21 46692388 N chr21 46692573 N DEL 8
SRR1766481.7896101 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766458.5689457 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766454.3140822 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766478.4157743 chr21 46692572 N chr21 46692664 N DUP 5
SRR1766461.5546154 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766452.2603472 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766470.4827682 chr21 46692579 N chr21 46692671 N DUP 10
SRR1766454.4475499 chr21 46692193 N chr21 46692564 N DEL 5
SRR1766451.1404094 chr21 46691923 N chr21 46692573 N DEL 5
SRR1766476.7331748 chr21 46691923 N chr21 46692573 N DEL 5
SRR1766449.9752047 chr21 46692572 N chr21 46692664 N DUP 5
SRR1766464.6243082 chr21 46692311 N chr21 46692589 N DEL 10
SRR1766479.12925842 chr21 46691923 N chr21 46692573 N DEL 5
SRR1766454.4686249 chr21 46691923 N chr21 46692573 N DEL 5
SRR1766471.1047566 chr21 46691941 N chr21 46692589 N DUP 10
SRR1766473.3242413 chr21 46691923 N chr21 46692573 N DEL 5
SRR1766444.6733882 chr21 46691923 N chr21 46692573 N DEL 5
SRR1766447.10489924 chr21 46692579 N chr21 46692671 N DUP 2
SRR1766478.630594 chr21 46692579 N chr21 46692671 N DUP 2
SRR1766479.10496384 chr21 46692579 N chr21 46692671 N DUP 2
SRR1766460.8476075 chr21 46692572 N chr21 46692664 N DUP 5
SRR1766466.10315026 chr21 46692044 N chr21 46692508 N DEL 3
SRR1766483.6751339 chr21 46692572 N chr21 46692664 N DUP 8
SRR1766442.36378806 chr21 46692579 N chr21 46692671 N DUP 4
SRR1766479.5975899 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766454.4838714 chr21 46692027 N chr21 46692584 N DEL 5
SRR1766442.24064084 chr21 46692028 N chr21 46692585 N DEL 5
SRR1766447.10847520 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766442.43173751 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766450.6968047 chr21 46692202 N chr21 46692573 N DEL 7
SRR1766472.3557867 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766445.8277325 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766483.6459969 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766483.11000449 chr21 46692311 N chr21 46692589 N DEL 8
SRR1766482.3892203 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766459.4329808 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766445.7257402 chr21 46692579 N chr21 46692671 N DUP 5
SRR1766467.9976925 chr21 46692030 N chr21 46692587 N DEL 1
SRR1766481.2320907 chr21 46692311 N chr21 46692589 N DEL 6
SRR1766481.10206302 chr21 46692506 N chr21 46692598 N DUP 5
SRR1766467.6428920 chr21 46692579 N chr21 46692671 N DUP 6
SRR1766442.45738844 chr21 46692579 N chr21 46692671 N DUP 11
SRR1766442.8213125 chr21 46692579 N chr21 46692671 N DUP 15
SRR1766454.10116196 chr21 46692146 N chr21 46692610 N DEL 8
SRR1766480.6907702 chr21 46692053 N chr21 46692610 N DEL 3
SRR1766486.2954728 chr21 46692053 N chr21 46692610 N DEL 2
SRR1766447.6488578 chr21 46692052 N chr21 46692609 N DEL 2
SRR1766486.4534790 chr21 46692159 N chr21 46692623 N DEL 5
SRR1766448.4546985 chr21 46692015 N chr21 46692665 N DEL 5
SRR1766466.4447283 chr21 46692197 N chr21 46692661 N DEL 5
SRR1766444.5139845 chr9 125623367 N chr9 125623678 N DUP 5
SRR1766477.431558 chr9 125623549 N chr9 125623664 N DUP 1
SRR1766471.7077942 chr9 125623558 N chr9 125623633 N DUP 3
SRR1766465.8775750 chr9 125623453 N chr9 125623805 N DUP 2
SRR1766442.32485493 chr2 159874943 N chr2 159875000 N DEL 7
SRR1766457.3132729 chr2 159874943 N chr2 159875000 N DEL 7
SRR1766463.9442736 chr2 159874943 N chr2 159875000 N DEL 7
SRR1766456.2761193 chr2 159874943 N chr2 159875000 N DEL 7
SRR1766467.421770 chr2 159874943 N chr2 159875000 N DEL 7
SRR1766462.7202058 chr2 159874943 N chr2 159875000 N DEL 7
SRR1766485.3731305 chr2 159874926 N chr2 159875010 N DEL 5
SRR1766474.8423523 chr2 159874930 N chr2 159875014 N DEL 1
SRR1766466.1799476 chr2 159874934 N chr2 159875068 N DEL 5
SRR1766445.10390828 chr7 107680010 N chr7 107680071 N DEL 3
SRR1766467.1699318 chr7 107680010 N chr7 107680071 N DEL 4
SRR1766448.11080743 chr7 107680025 N chr7 107680087 N DUP 9
SRR1766460.11257622 chr7 107679963 N chr7 107680055 N DEL 11
SRR1766466.5498767 chr6 16616704 N chr6 16616761 N DEL 11
SRR1766470.5382874 chr13 113734047 N chr13 113734113 N DEL 7
SRR1766485.11596683 chr16 28442261 N chr16 28442472 N DEL 14
SRR1766475.7129747 chr2 4449607 N chr2 4449787 N DUP 14
SRR1766481.825180 chr3 79850093 N chr3 79850143 N DUP 2
SRR1766467.10393611 chr14 70477693 N chr14 70477774 N DUP 11
SRR1766453.7766679 chr14 70477693 N chr14 70477774 N DUP 5
SRR1766477.11410261 chr14 70477609 N chr14 70477806 N DEL 2
SRR1766463.5291959 chr4 163537154 N chr4 163537216 N DEL 5
SRR1766482.3348683 chr1 15494709 N chr1 15495008 N DEL 1
SRR1766442.23424258 chrY 10763749 N chrY 10763863 N DUP 5
SRR1766442.22049114 chr20 61173321 N chr20 61173422 N DEL 5
SRR1766463.6801109 chr20 61173334 N chr20 61173415 N DEL 10
SRR1766470.5927921 chr20 61173354 N chr20 61173415 N DEL 5
SRR1766455.7617254 chr20 61173354 N chr20 61173415 N DEL 11
SRR1766451.2071800 chr20 61173395 N chr20 61173574 N DEL 5
SRR1766483.9131959 chr20 61173389 N chr20 61173450 N DEL 5
SRR1766461.10203077 chr20 61173354 N chr20 61173415 N DEL 5
SRR1766468.4218410 chr20 61173396 N chr20 61173575 N DEL 20
SRR1766473.2005969 chr20 61173480 N chr20 61173659 N DEL 5
SRR1766450.6120215 chr20 61173345 N chr20 61173523 N DEL 5
SRR1766450.2697726 chr20 61173336 N chr20 61173595 N DEL 3
SRR1766476.8507470 chr20 61173438 N chr20 61173834 N DEL 3
SRR1766450.9665060 chr20 61173424 N chr20 61173860 N DEL 5
SRR1766458.3818111 chr8 67831163 N chr8 67831216 N DEL 7
SRR1766457.6255076 chr8 67831217 N chr8 67831268 N DEL 17
SRR1766442.47100960 chr8 67831206 N chr8 67831280 N DEL 4
SRR1766448.970184 chr8 67831206 N chr8 67831280 N DEL 3
SRR1766481.10486062 chr2 108765460 N chr2 108765989 N DEL 24
SRR1766482.12785928 chr2 108765372 N chr2 108765560 N DUP 10
SRR1766477.8843202 chr2 108765656 N chr2 108766008 N DEL 5
SRR1766458.6437249 chr2 108765517 N chr2 108765872 N DEL 5
SRR1766468.3654191 chr2 108765585 N chr2 108765940 N DEL 15
SRR1766445.2550083 chr4 9981210 N chr4 9981460 N DEL 20
SRR1766446.8711744 chr4 9981273 N chr4 9981489 N DEL 13
SRR1766447.8246958 chr4 9981302 N chr4 9981485 N DEL 5
SRR1766472.3725687 chr4 9981304 N chr4 9981481 N DEL 7
SRR1766461.6242935 chr4 9981313 N chr4 9981502 N DEL 5
SRR1766443.9746749 chr4 9981325 N chr4 9981481 N DEL 4
SRR1766451.1242499 chr4 9981407 N chr4 9981494 N DEL 5
SRR1766476.10307082 chr4 9981324 N chr4 9981419 N DUP 6
SRR1766481.2654541 chr4 9981324 N chr4 9981419 N DUP 9
SRR1766463.689315 chr4 9981324 N chr4 9981419 N DUP 12
SRR1766442.35794695 chr4 9981324 N chr4 9981419 N DUP 15
SRR1766442.40441387 chr4 9981324 N chr4 9981419 N DUP 10
SRR1766481.8003392 chr4 9981348 N chr4 9981458 N DUP 8
SRR1766447.11182975 chr4 9981366 N chr4 9981514 N DUP 5
SRR1766482.6149530 chr4 9981355 N chr4 9981500 N DUP 7
SRR1766461.718464 chr4 9981366 N chr4 9981455 N DUP 5
SRR1766463.7436736 chr4 9981355 N chr4 9981441 N DUP 10
SRR1766465.10929225 chr4 9981386 N chr4 9981501 N DUP 8
SRR1766484.5025744 chr4 9981386 N chr4 9981501 N DUP 8
SRR1766479.13025578 chr4 9981386 N chr4 9981501 N DUP 8
SRR1766455.6329570 chr2 234899245 N chr2 234899296 N DEL 7
SRR1766454.1305986 chr2 234899245 N chr2 234899296 N DEL 8
SRR1766474.1433164 chr2 234899245 N chr2 234899296 N DEL 12
SRR1766475.6598973 chr2 234899245 N chr2 234899296 N DEL 13
SRR1766451.9590040 chr9 65201754 N chr9 65201876 N DEL 3
SRR1766459.11359228 chr7 71592649 N chr7 71592726 N DUP 6
SRR1766442.4487998 chr7 71592663 N chr7 71592727 N DEL 1
SRR1766445.10074319 chr7 71592661 N chr7 71592725 N DEL 3
SRR1766448.8533779 chr7 71592660 N chr7 71592724 N DEL 4
SRR1766463.71635 chr7 71592660 N chr7 71592724 N DEL 4
SRR1766460.4989477 chr7 71592662 N chr7 71592716 N DEL 12
SRR1766474.8212249 chr7 71592662 N chr7 71592721 N DEL 7
SRR1766465.6964994 chr18 54806602 N chr18 54806716 N DUP 5
SRR1766486.5653256 chr20 37572380 N chr20 37572432 N DEL 7
SRR1766442.29211788 chr20 37572379 N chr20 37572435 N DEL 7
SRR1766447.10317714 chr20 37572379 N chr20 37572540 N DEL 9
SRR1766484.9220929 chr20 37572377 N chr20 37572546 N DEL 7
SRR1766485.4522751 chr20 37572377 N chr20 37572546 N DEL 7
SRR1766459.9617478 chr20 37572372 N chr20 37572558 N DEL 4
SRR1766448.4869614 chr20 37572382 N chr20 37572566 N DEL 7
SRR1766451.8313100 chr20 37572386 N chr20 37572566 N DEL 4
SRR1766482.1154359 chr20 37572380 N chr20 37572568 N DEL 7
SRR1766482.1517502 chr20 37572379 N chr20 37572567 N DEL 7
SRR1766451.6940329 chr20 37572379 N chr20 37572571 N DEL 7
SRR1766470.3871151 chr3 126008535 N chr3 126008616 N DUP 3
SRR1766444.130694 chr3 126008563 N chr3 126008665 N DEL 23
SRR1766483.8361032 chr18 71428589 N chr18 71428738 N DEL 5
SRR1766462.37377 chr5 125632894 N chr5 125633008 N DUP 21
SRR1766445.1525882 chr5 125632894 N chr5 125633007 N DUP 20
SRR1766467.1085788 chr2 239017529 N chr2 239018448 N DEL 4
SRR1766478.5604409 chr2 239017597 N chr2 239017992 N DEL 9
SRR1766450.6179352 chr2 239017444 N chr2 239018267 N DEL 10
SRR1766483.5890898 chr2 239017691 N chr2 239018494 N DEL 7
SRR1766452.3129435 chr2 239017691 N chr2 239017942 N DEL 5
SRR1766464.6106891 chr2 239017750 N chr2 239018267 N DEL 10
SRR1766476.7027381 chr2 239017793 N chr2 239018364 N DEL 5
SRR1766468.913407 chr2 239017397 N chr2 239017752 N DEL 6
SRR1766465.3719918 chr2 239017885 N chr2 239018358 N DEL 5
SRR1766448.8637884 chr2 239017383 N chr2 239017884 N DUP 5
SRR1766467.9175636 chr2 239017418 N chr2 239017919 N DUP 3
SRR1766442.21311475 chr2 239017850 N chr2 239017951 N DUP 5
SRR1766475.7767158 chr2 239017398 N chr2 239017901 N DEL 2
SRR1766471.3041204 chr2 239017445 N chr2 239017948 N DEL 5
SRR1766479.13180651 chr2 239017381 N chr2 239018046 N DUP 6
SRR1766444.6678286 chr2 239017965 N chr2 239018508 N DUP 12
SRR1766478.5604409 chr2 239017403 N chr2 239017962 N DEL 1
SRR1766483.4941127 chr2 239017383 N chr2 239018102 N DUP 5
SRR1766484.546083 chr2 239017380 N chr2 239018103 N DUP 8
SRR1766445.1366370 chr2 239017430 N chr2 239018149 N DUP 7
SRR1766480.6616642 chr2 239017994 N chr2 239018157 N DUP 6
SRR1766453.1642506 chr2 239017994 N chr2 239018157 N DUP 6
SRR1766444.758361 chr2 239017617 N chr2 239018182 N DUP 5
SRR1766476.1595318 chr2 239017412 N chr2 239018077 N DEL 5
SRR1766467.1228826 chr2 239018003 N chr2 239018118 N DEL 5
SRR1766474.4871269 chr2 239017470 N chr2 239018239 N DUP 5
SRR1766461.10118290 chr2 239017722 N chr2 239018235 N DUP 2
SRR1766458.8387934 chr2 239017414 N chr2 239018185 N DEL 5
SRR1766462.7505371 chr2 239018313 N chr2 239018364 N DEL 5
SRR1766463.6243033 chr2 239018166 N chr2 239018269 N DEL 2
SRR1766482.4766478 chr2 239017443 N chr2 239018266 N DEL 5
SRR1766479.1954541 chr2 239017835 N chr2 239018258 N DEL 1
SRR1766470.1261992 chr2 239018195 N chr2 239018298 N DEL 10
SRR1766444.2839974 chr2 239017418 N chr2 239018389 N DUP 5
SRR1766467.7002710 chr2 239017689 N chr2 239018358 N DEL 5
SRR1766460.10796559 chr2 239017437 N chr2 239018360 N DEL 5
SRR1766459.10322999 chr2 239017442 N chr2 239018365 N DEL 5
SRR1766476.8783596 chr2 239017439 N chr2 239018362 N DEL 5
SRR1766445.6011786 chr2 239018009 N chr2 239018386 N DEL 7
SRR1766450.6971947 chr18 12873899 N chr18 12874053 N DEL 5
SRR1766481.4886833 chr18 12874110 N chr18 12874268 N DEL 4
SRR1766462.521502 chr9 37918523 N chr9 37918584 N DEL 17
SRR1766480.6460053 chr9 37918523 N chr9 37918584 N DEL 17
SRR1766486.4586852 chr9 37918523 N chr9 37918584 N DEL 26
SRR1766484.288518 chr9 37918523 N chr9 37918584 N DEL 26
SRR1766448.4003445 chr5 23894222 N chr5 23894739 N DEL 1
SRR1766466.7090593 chr5 23894795 N chr5 23895140 N DEL 3
SRR1766484.1566948 chr19 39153429 N chr19 39153611 N DUP 10
SRR1766468.3243441 chr19 39153429 N chr19 39153611 N DUP 15
SRR1766450.181568 chr19 39153437 N chr19 39153619 N DUP 5
SRR1766472.614869 chr19 39153429 N chr19 39153611 N DUP 15
SRR1766475.5294056 chr19 39153429 N chr19 39153611 N DUP 20
SRR1766442.35551343 chr19 39153429 N chr19 39153611 N DUP 34
SRR1766452.5236743 chr19 39153429 N chr19 39153611 N DUP 36
SRR1766472.11328600 chr19 39153429 N chr19 39153611 N DUP 46
SRR1766468.2261208 chr12 86502818 N chr12 86502946 N DEL 25
SRR1766462.241223 chr12 86502860 N chr12 86502938 N DUP 5
SRR1766454.1822591 chr12 86502963 N chr12 86503678 N DEL 11
SRR1766446.8169602 chr12 86502963 N chr12 86503678 N DEL 9
SRR1766459.9954864 chr12 86502963 N chr12 86503678 N DEL 9
SRR1766467.4198919 chr12 86502963 N chr12 86503678 N DEL 9
SRR1766451.747059 chr12 86502963 N chr12 86503678 N DEL 16
SRR1766452.10672015 chr12 86502936 N chr12 86503678 N DEL 16
SRR1766479.8499000 chr12 86502936 N chr12 86503678 N DEL 16
SRR1766483.12476605 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766458.1954919 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766475.8305492 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766470.2589770 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766476.3414480 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766486.5654796 chr12 86503015 N chr12 86503757 N DEL 16
SRR1766459.5270646 chr12 86503042 N chr12 86503095 N DEL 7
SRR1766467.4198919 chr12 86502796 N chr12 86502993 N DEL 4
SRR1766473.8354185 chr12 86503067 N chr12 86503784 N DEL 7
SRR1766447.5951024 chr12 86503015 N chr12 86503757 N DEL 9
SRR1766458.5674146 chr12 86503015 N chr12 86503757 N DEL 9
SRR1766451.5670355 chr12 86503015 N chr12 86503757 N DEL 9
SRR1766442.28799040 chr12 86502799 N chr12 86503764 N DEL 8
SRR1766482.11208037 chr12 86502869 N chr12 86503765 N DEL 7
SRR1766483.6704966 chr12 86503067 N chr12 86503430 N DEL 6
SRR1766442.36802092 chr12 86503179 N chr12 86503798 N DUP 7
SRR1766450.1765989 chr12 86503218 N chr12 86503477 N DUP 7
SRR1766443.2252384 chr12 86503218 N chr12 86503477 N DUP 10
SRR1766473.6911452 chr12 86503218 N chr12 86503781 N DUP 9
SRR1766481.6768283 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766452.4805788 chr12 86503218 N chr12 86503623 N DUP 12
SRR1766447.4420733 chr12 86503218 N chr12 86503623 N DUP 12
SRR1766459.8578456 chr12 86503218 N chr12 86503477 N DUP 7
SRR1766450.1765989 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766448.4502342 chr12 86503218 N chr12 86503623 N DUP 11
SRR1766483.7132869 chr12 86503218 N chr12 86503623 N DUP 11
SRR1766480.7626066 chr12 86503218 N chr12 86503623 N DUP 10
SRR1766472.10981418 chr12 86503218 N chr12 86503477 N DUP 7
SRR1766473.8354185 chr12 86503218 N chr12 86503623 N DUP 9
SRR1766478.3619440 chr12 86503218 N chr12 86503623 N DUP 8
SRR1766468.2453815 chr12 86503218 N chr12 86503477 N DUP 7
SRR1766467.8295699 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766476.3671024 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766442.31246583 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766472.11196187 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766479.8949922 chr12 86503218 N chr12 86503477 N DUP 7
SRR1766486.7741371 chr12 86503218 N chr12 86503477 N DUP 7
SRR1766478.10032979 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766472.347763 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766482.8823903 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766483.9951095 chr12 86503119 N chr12 86503218 N DEL 7
SRR1766465.4167578 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766442.37357185 chr12 86503013 N chr12 86503218 N DEL 7
SRR1766470.3716674 chr12 86503013 N chr12 86503218 N DEL 7
SRR1766461.4316363 chr12 86503013 N chr12 86503218 N DEL 7
SRR1766446.6686697 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766486.8227023 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766457.396067 chr12 86503040 N chr12 86503218 N DEL 7
SRR1766460.4683302 chr12 86502997 N chr12 86503077 N DUP 3
SRR1766474.1438118 chr12 86503013 N chr12 86503218 N DEL 7
SRR1766448.4914540 chr12 86503014 N chr12 86503219 N DEL 7
SRR1766478.2505300 chr12 86503016 N chr12 86503221 N DEL 7
SRR1766446.493056 chr12 86503040 N chr12 86503218 N DEL 7
SRR1766481.5841633 chr12 86503040 N chr12 86503218 N DEL 7
SRR1766485.8861738 chr12 86503040 N chr12 86503218 N DEL 9
SRR1766444.6279104 chr12 86503028 N chr12 86503229 N DEL 2
SRR1766478.11617144 chr12 86503121 N chr12 86503624 N DEL 3
SRR1766450.9708057 chr12 86503115 N chr12 86503239 N DEL 2
SRR1766484.10211309 chr12 86503121 N chr12 86503243 N DEL 5
SRR1766479.10755295 chr12 86503121 N chr12 86503243 N DEL 6
SRR1766482.11208037 chr12 86503121 N chr12 86503243 N DEL 9
SRR1766452.6321681 chr12 86503121 N chr12 86503243 N DEL 9
SRR1766458.4940290 chr12 86503121 N chr12 86503243 N DEL 9
SRR1766479.1221450 chr12 86503121 N chr12 86503243 N DEL 9
SRR1766482.2192603 chr12 86503121 N chr12 86503243 N DEL 9
SRR1766485.421895 chr12 86503121 N chr12 86503243 N DEL 9
SRR1766476.7877247 chr12 86503121 N chr12 86503243 N DEL 9
SRR1766485.421895 chr12 86503121 N chr12 86503349 N DEL 2
SRR1766442.7022776 chr12 86503042 N chr12 86503349 N DEL 3
SRR1766483.2408027 chr12 86503026 N chr12 86503254 N DEL 4
SRR1766485.8521350 chr12 86503015 N chr12 86503349 N DEL 7
SRR1766444.5931563 chr12 86503218 N chr12 86503781 N DUP 9
SRR1766463.921458 chr12 86503171 N chr12 86503786 N DUP 9
SRR1766482.238544 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766454.7950493 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766467.6692147 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766442.27219978 chr12 86503015 N chr12 86503349 N DEL 7
SRR1766445.3146777 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766484.262550 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766457.1230279 chr12 86502840 N chr12 86503351 N DEL 7
SRR1766466.3995621 chr12 86502840 N chr12 86503351 N DEL 7
SRR1766468.2261208 chr12 86502840 N chr12 86503351 N DEL 7
SRR1766484.685932 chr12 86503067 N chr12 86503218 N DEL 7
SRR1766486.344163 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766478.10032979 chr12 86502797 N chr12 86503354 N DEL 7
SRR1766459.5270646 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766444.635520 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766442.46745300 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766449.7259289 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766447.6081674 chr12 86503067 N chr12 86503218 N DEL 7
SRR1766453.9763572 chr12 86503067 N chr12 86503218 N DEL 7
SRR1766446.493056 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766459.9954864 chr12 86503040 N chr12 86503218 N DEL 7
SRR1766478.11617144 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766486.9118110 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766481.5841633 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766447.4420733 chr12 86503067 N chr12 86503218 N DEL 7
SRR1766466.6703242 chr12 86503040 N chr12 86503218 N DEL 7
SRR1766467.8295699 chr12 86503067 N chr12 86503218 N DEL 7
SRR1766466.8416415 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766470.8861870 chr12 86503583 N chr12 86503796 N DEL 14
SRR1766442.31246583 chr12 86503009 N chr12 86503349 N DEL 9
SRR1766482.238544 chr12 86503583 N chr12 86503796 N DEL 12
SRR1766446.3770000 chr12 86503583 N chr12 86503796 N DEL 12
SRR1766461.7049418 chr12 86503015 N chr12 86503349 N DEL 7
SRR1766464.2335191 chr12 86502842 N chr12 86503353 N DEL 7
SRR1766464.689097 chr12 86503218 N chr12 86503623 N DUP 14
SRR1766450.8208644 chr12 86503015 N chr12 86503757 N DEL 13
SRR1766470.8861870 chr12 86503067 N chr12 86503784 N DEL 7
SRR1766474.293744 chr12 86503069 N chr12 86503836 N DEL 7
SRR1766479.1221450 chr12 86503067 N chr12 86503784 N DEL 7
SRR1766483.6704966 chr12 86503067 N chr12 86503784 N DEL 7
SRR1766471.10647577 chr12 86503040 N chr12 86503784 N DEL 9
SRR1766451.7805933 chr12 86503040 N chr12 86503784 N DEL 9
SRR1766486.5654796 chr12 86503042 N chr12 86503095 N DEL 7
SRR1766465.4167578 chr12 86503040 N chr12 86503784 N DEL 9
SRR1766448.8535540 chr12 86503067 N chr12 86503430 N DEL 7
SRR1766460.9088046 chr12 86503040 N chr12 86503784 N DEL 11
SRR1766443.4173443 chr12 86503067 N chr12 86503430 N DEL 7
SRR1766442.25669914 chr12 86503040 N chr12 86503430 N DEL 7
SRR1766458.5674146 chr12 86503040 N chr12 86503430 N DEL 7
SRR1766442.9009358 chr12 86503015 N chr12 86503095 N DEL 1
SRR1766476.1227802 chr12 86503452 N chr12 86503753 N DUP 11
SRR1766483.10274482 chr12 86503121 N chr12 86503478 N DEL 5
SRR1766485.8726289 chr12 86503121 N chr12 86503478 N DEL 5
SRR1766462.1627407 chr12 86503121 N chr12 86503478 N DEL 9
SRR1766458.1954919 chr12 86503088 N chr12 86503516 N DUP 9
SRR1766454.7315669 chr12 86503146 N chr12 86503480 N DEL 14
SRR1766445.10648095 chr12 86503015 N chr12 86503478 N DEL 16
SRR1766463.3142576 chr12 86503015 N chr12 86503478 N DEL 10
SRR1766442.6255515 chr12 86503015 N chr12 86503478 N DEL 9
SRR1766472.347763 chr12 86503015 N chr12 86503478 N DEL 9
SRR1766457.5215980 chr12 86503015 N chr12 86503478 N DEL 9
SRR1766485.5136630 chr12 86503015 N chr12 86503478 N DEL 9
SRR1766486.1012353 chr12 86502870 N chr12 86503487 N DEL 6
SRR1766473.4693034 chr12 86503026 N chr12 86503489 N DEL 4
SRR1766475.7871132 chr12 86503026 N chr12 86503489 N DEL 4
SRR1766444.6279104 chr12 86503030 N chr12 86503491 N DEL 2
SRR1766451.6688853 chr12 86502793 N chr12 86503504 N DEL 5
SRR1766486.7741371 chr12 86503028 N chr12 86503512 N DEL 5
SRR1766482.11393718 chr12 86503413 N chr12 86503583 N DUP 7
SRR1766480.8743910 chr12 86503413 N chr12 86503583 N DUP 9
SRR1766469.1182654 chr12 86503413 N chr12 86503583 N DUP 9
SRR1766447.10962633 chr12 86503413 N chr12 86503583 N DUP 9
SRR1766472.11196187 chr12 86503583 N chr12 86503796 N DEL 11
SRR1766448.5492515 chr12 86503583 N chr12 86503796 N DEL 13
SRR1766450.5038210 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766469.3903658 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766479.5023210 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766452.5596729 chr12 86503218 N chr12 86503623 N DUP 16
SRR1766447.1817290 chr12 86502797 N chr12 86503225 N DEL 7
SRR1766464.7231028 chr12 86502797 N chr12 86503225 N DEL 7
SRR1766474.1438118 chr12 86503015 N chr12 86503243 N DEL 7
SRR1766476.7877247 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766467.7770464 chr12 86503015 N chr12 86503243 N DEL 7
SRR1766471.8860052 chr12 86503015 N chr12 86503243 N DEL 7
SRR1766459.9443104 chr12 86503015 N chr12 86503243 N DEL 7
SRR1766456.867414 chr12 86503015 N chr12 86503243 N DEL 7
SRR1766452.5769201 chr12 86503015 N chr12 86503243 N DEL 7
SRR1766442.9009358 chr12 86502840 N chr12 86502991 N DEL 7
SRR1766449.7593825 chr12 86503042 N chr12 86503243 N DEL 9
SRR1766486.10254790 chr12 86503015 N chr12 86503757 N DEL 9
SRR1766457.1208404 chr12 86503016 N chr12 86503758 N DEL 9
SRR1766461.9798580 chr12 86503027 N chr12 86503769 N DEL 3
SRR1766454.7950493 chr12 86503040 N chr12 86503784 N DEL 8
SRR1766445.3268784 chr12 86503040 N chr12 86503784 N DEL 12
SRR1766476.7549176 chr12 86503044 N chr12 86503811 N DEL 5
SRR1766474.4794869 chr12 86503027 N chr12 86503769 N DEL 3
SRR1766448.9201487 chr12 86503040 N chr12 86503784 N DEL 7
SRR1766453.2439139 chr12 86503013 N chr12 86503784 N DEL 7
SRR1766486.4077096 chr12 86503013 N chr12 86503784 N DEL 7
SRR1766483.6302124 chr12 86503013 N chr12 86503784 N DEL 7
SRR1766471.8919009 chr12 86503014 N chr12 86503785 N DEL 7
SRR1766452.4805788 chr12 86503014 N chr12 86503785 N DEL 7
SRR1766486.1012353 chr12 86503014 N chr12 86503785 N DEL 7
SRR1766474.11369929 chr12 86503015 N chr12 86503786 N DEL 7
SRR1766473.1010296 chr12 86502841 N chr12 86503789 N DEL 7
SRR1766485.6605288 chr12 86503218 N chr12 86503781 N DUP 9
SRR1766478.587340 chr12 86503040 N chr12 86503786 N DEL 7
SRR1766465.10237541 chr12 86503040 N chr12 86503786 N DEL 7
SRR1766450.1823113 chr12 86503119 N chr12 86503403 N DEL 8
SRR1766471.2656444 chr12 86503040 N chr12 86503786 N DEL 6
SRR1766442.6255515 chr12 86503119 N chr12 86503403 N DEL 8
SRR1766457.2510486 chr12 86503218 N chr12 86503623 N DUP 14
SRR1766482.10220538 chr12 86503013 N chr12 86503786 N DEL 6
SRR1766485.5007137 chr12 86503119 N chr12 86503403 N DEL 8
SRR1766466.552884 chr12 86503119 N chr12 86503403 N DEL 8
SRR1766463.5580732 chr12 86503070 N chr12 86503477 N DUP 8
SRR1766474.4900596 chr12 86502841 N chr12 86503791 N DEL 6
SRR1766481.4531237 chr12 86502797 N chr12 86503793 N DEL 6
SRR1766447.10962633 chr12 86503173 N chr12 86503937 N DEL 17
SRR1766448.4914540 chr12 86503173 N chr12 86503937 N DEL 17
SRR1766475.8163142 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766442.36290555 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766475.5221749 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766479.8525665 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766480.7626066 chr12 86503679 N chr12 86503937 N DEL 18
SRR1766450.5038210 chr12 86502870 N chr12 86503899 N DEL 4
SRR1766458.6030704 chr12 86503000 N chr12 86503937 N DEL 19
SRR1766453.1978957 chr12 86502842 N chr12 86503937 N DEL 17
SRR1766473.6012036 chr12 86502842 N chr12 86503937 N DEL 17
SRR1766442.32326032 chr12 86502799 N chr12 86503940 N DEL 12
SRR1766474.10867554 chr12 86503002 N chr12 86503939 N DEL 13
SRR1766442.46745300 chr12 86503029 N chr12 86503947 N DEL 5
SRR1766465.5883884 chr12 86502799 N chr12 86503940 N DEL 12
SRR1766466.6703242 chr12 86503029 N chr12 86503945 N DEL 7
SRR1766444.7137215 chr5 1422500 N chr5 1423283 N DEL 5
SRR1766442.151381 chr5 1422500 N chr5 1422763 N DEL 5
SRR1766466.2603788 chr5 1422500 N chr5 1422763 N DEL 5
SRR1766454.5392723 chr5 1422500 N chr5 1422763 N DEL 5
SRR1766443.1518904 chr5 1422508 N chr5 1422621 N DEL 14
SRR1766451.6565019 chr5 1422521 N chr5 1422598 N DEL 10
SRR1766457.9437292 chr5 1422521 N chr5 1422598 N DEL 5
SRR1766467.4156380 chr5 1422521 N chr5 1422598 N DEL 5
SRR1766447.4323510 chr5 1422521 N chr5 1422598 N DEL 5
SRR1766467.4733064 chr5 1422521 N chr5 1422598 N DEL 5
SRR1766453.4421351 chr5 1422521 N chr5 1422598 N DEL 10
SRR1766460.10481947 chr5 1422521 N chr5 1422598 N DEL 15
SRR1766442.31006958 chr5 1422521 N chr5 1422598 N DEL 20
SRR1766446.7632159 chr5 1422521 N chr5 1422598 N DEL 10
SRR1766462.7793342 chr5 1422521 N chr5 1422598 N DEL 10
SRR1766467.4156380 chr5 1422929 N chr5 1423232 N DEL 14
SRR1766442.29156634 chr5 1422580 N chr5 1422913 N DUP 8
SRR1766464.3065887 chr5 1422606 N chr5 1422755 N DUP 7
SRR1766479.8661184 chr5 1422595 N chr5 1422674 N DEL 9
SRR1766456.3987549 chr5 1422962 N chr5 1423037 N DEL 15
SRR1766470.2632024 chr5 1422726 N chr5 1423283 N DEL 7
SRR1766452.8274267 chr5 1422659 N chr5 1423366 N DEL 15
SRR1766446.8387355 chr5 1422721 N chr5 1422904 N DEL 15
SRR1766475.8622079 chr5 1422726 N chr5 1423021 N DEL 7
SRR1766475.933545 chr5 1422726 N chr5 1422909 N DEL 8
SRR1766450.1367771 chr5 1422601 N chr5 1422750 N DUP 7
SRR1766444.6197426 chr5 1422604 N chr5 1422753 N DUP 7
SRR1766459.11405611 chr5 1422743 N chr5 1422926 N DEL 10
SRR1766483.9581925 chr5 1422645 N chr5 1422904 N DEL 14
SRR1766455.6400678 chr5 1422574 N chr5 1423281 N DUP 1
SRR1766459.531360 chr5 1422613 N chr5 1423282 N DUP 8
SRR1766451.6565019 chr5 1422598 N chr5 1422893 N DUP 17
SRR1766455.4750083 chr5 1422770 N chr5 1423365 N DEL 4
SRR1766461.6318056 chr5 1422704 N chr5 1423187 N DEL 10
SRR1766474.1471987 chr5 1422659 N chr5 1423068 N DEL 5
SRR1766448.1305371 chr5 1422693 N chr5 1423288 N DEL 5
SRR1766450.4864914 chr5 1422617 N chr5 1423288 N DEL 5
SRR1766450.2401568 chr5 1422710 N chr5 1423115 N DUP 13
SRR1766464.10125897 chr5 1422633 N chr5 1422712 N DEL 7
SRR1766455.6400678 chr5 1422562 N chr5 1422675 N DUP 9
SRR1766454.5392723 chr5 1422712 N chr5 1422929 N DUP 8
SRR1766445.4143533 chr5 1422643 N chr5 1422754 N DUP 3
SRR1766450.1367771 chr5 1422571 N chr5 1422648 N DEL 5
SRR1766447.10224711 chr5 1422510 N chr5 1422807 N DUP 5
SRR1766475.10436697 chr5 1422783 N chr5 1422858 N DEL 5
SRR1766442.151381 chr5 1422704 N chr5 1422851 N DEL 9
SRR1766468.1017296 chr5 1422659 N chr5 1423366 N DEL 11
SRR1766485.5893723 chr5 1422562 N chr5 1422933 N DUP 5
SRR1766467.7203391 chr5 1422686 N chr5 1422907 N DEL 18
SRR1766442.17409400 chr5 1422735 N chr5 1422918 N DEL 9
SRR1766464.9260686 chr5 1422678 N chr5 1422751 N DUP 7
SRR1766486.11290022 chr5 1422919 N chr5 1423030 N DUP 5
SRR1766452.3373823 chr5 1423394 N chr5 1423531 N DUP 22
SRR1766444.2682053 chr5 1423121 N chr5 1423394 N DEL 26
SRR1766486.6287211 chr5 1422562 N chr5 1423157 N DUP 5
SRR1766458.5605945 chr5 1422602 N chr5 1423087 N DEL 3
SRR1766470.913081 chr5 1422682 N chr5 1423163 N DUP 3
SRR1766461.559133 chr5 1422993 N chr5 1423180 N DEL 18
SRR1766463.7541807 chr5 1422640 N chr5 1423199 N DEL 23
SRR1766442.23686459 chr5 1422583 N chr5 1423180 N DEL 6
SRR1766477.2435146 chr5 1422586 N chr5 1423183 N DEL 3
SRR1766448.5245341 chr5 1422628 N chr5 1423225 N DEL 25
SRR1766480.6248292 chr5 1422949 N chr5 1423250 N DEL 16
SRR1766479.2081966 chr5 1422545 N chr5 1423218 N DEL 5
SRR1766469.1984519 chr5 1422778 N chr5 1423225 N DEL 9
SRR1766458.4364186 chr5 1422887 N chr5 1423262 N DEL 10
SRR1766448.4973613 chr5 1422598 N chr5 1423345 N DEL 10
SRR1766455.8397902 chr5 1422971 N chr5 1423356 N DEL 20
SRR1766481.8306630 chr5 1422881 N chr5 1423330 N DEL 10
SRR1766457.5667459 chr5 1422960 N chr5 1423345 N DEL 13
SRR1766452.3551185 chr5 1423356 N chr5 1423419 N DUP 26
SRR1766473.8570077 chr5 1422960 N chr5 1423421 N DEL 17
SRR1766442.38880851 chr5 1422960 N chr5 1423421 N DEL 15
SRR1766442.37700247 chr5 1422771 N chr5 1423478 N DEL 5
SRR1766443.5896391 chr5 1422587 N chr5 1423482 N DEL 2
SRR1766480.4762618 chr5 1423056 N chr5 1423505 N DEL 5
SRR1766484.3203624 chr5 1423056 N chr5 1423505 N DEL 5
SRR1766485.2364021 chr7 79625289 N chr7 79625731 N DEL 19
SRR1766460.5126526 chr7 79625289 N chr7 79625731 N DEL 15
SRR1766480.2526661 chr7 79625289 N chr7 79625731 N DEL 13
SRR1766463.3156830 chr7 79625387 N chr7 79625527 N DUP 3
SRR1766473.11175073 chr7 79625387 N chr7 79625546 N DUP 13
SRR1766442.12609679 chr7 79625272 N chr7 79625565 N DUP 13
SRR1766480.1090496 chr7 79625186 N chr7 79625493 N DEL 4
SRR1766463.6259944 chr7 79625272 N chr7 79625565 N DUP 1
SRR1766482.7370956 chr7 79625272 N chr7 79625565 N DUP 1
SRR1766483.4786567 chr7 79625564 N chr7 79625619 N DUP 2
SRR1766476.3754791 chr7 79625437 N chr7 79625575 N DEL 13
SRR1766443.6920293 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766457.7808506 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766474.7472757 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766463.5958978 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766474.259067 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766448.9678324 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766477.11399962 chr7 79625303 N chr7 79625575 N DEL 13
SRR1766460.10637313 chr7 79625262 N chr7 79625577 N DEL 13
SRR1766457.3942266 chr7 79625263 N chr7 79625578 N DEL 12
SRR1766443.6212544 chr7 79625269 N chr7 79625584 N DEL 6
SRR1766449.1720211 chr7 79625579 N chr7 79625640 N DEL 2
SRR1766453.397342 chr7 79625282 N chr7 79625682 N DEL 9
SRR1766446.7835646 chr7 79625282 N chr7 79625682 N DEL 9
SRR1766465.7139258 chr7 79625585 N chr7 79625691 N DEL 4
SRR1766462.4258862 chr7 79625585 N chr7 79625691 N DEL 4
SRR1766482.641648 chr7 79625585 N chr7 79625691 N DEL 3
SRR1766469.1407303 chr7 79625585 N chr7 79625691 N DEL 2
SRR1766473.1050873 chr7 79625585 N chr7 79625691 N DEL 1
SRR1766455.769442 chr7 79625404 N chr7 79625731 N DEL 17
SRR1766458.3622690 chr7 79625404 N chr7 79625731 N DEL 17
SRR1766460.6574941 chr7 79625277 N chr7 79625743 N DEL 3
SRR1766485.3527106 chr7 79625267 N chr7 79625733 N DEL 13
SRR1766478.1821811 chr7 79625266 N chr7 79625732 N DEL 14
SRR1766442.32985031 chr7 79625404 N chr7 79625731 N DEL 20
SRR1766448.4254032 chr7 79625404 N chr7 79625731 N DEL 20
SRR1766442.8894332 chr7 79625289 N chr7 79625731 N DEL 20
SRR1766473.10770663 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766452.1963307 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766482.608962 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766485.7101525 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766475.5230133 chr7 79625731 N chr7 79625802 N DUP 20
SRR1766484.2449073 chr7 79625308 N chr7 79625982 N DEL 7
SRR1766452.6232821 chr7 79625265 N chr7 79625982 N DEL 7
SRR1766476.8620447 chr2 195568522 N chr2 195568699 N DUP 13
SRR1766486.3359303 chr2 195568522 N chr2 195568650 N DUP 9
SRR1766452.5552961 chr2 195568537 N chr2 195568714 N DUP 1
SRR1766444.965161 chr2 195568522 N chr2 195568699 N DUP 11
SRR1766482.10930402 chr2 195568575 N chr2 195568754 N DEL 5
SRR1766462.7625354 chrY 26648574 N chrY 26648723 N DUP 9
SRR1766453.8226183 chrY 26648578 N chrY 26648692 N DUP 5
SRR1766442.41109618 chrY 26648611 N chrY 26648667 N DEL 7
SRR1766476.4032404 chr9 65463226 N chr9 65463334 N DEL 5
SRR1766453.2346912 chr9 65463292 N chr9 65463351 N DUP 5
SRR1766486.6542628 chr9 65463386 N chr9 65463866 N DEL 1
SRR1766472.55170 chr9 65463290 N chr9 65463409 N DUP 10
SRR1766450.7261467 chr9 65463409 N chr9 65463685 N DEL 5
SRR1766464.1495322 chr9 65463292 N chr9 65463439 N DUP 5
SRR1766459.9681421 chr9 65463460 N chr9 65464337 N DEL 5
SRR1766484.8049098 chr9 65463482 N chr9 65464110 N DEL 2
SRR1766442.1743688 chr9 65463370 N chr9 65463921 N DUP 5
SRR1766484.3958210 chr9 65463297 N chr9 65463390 N DEL 5
SRR1766447.6990334 chr9 65463294 N chr9 65463471 N DUP 1
SRR1766463.9567618 chr9 65463538 N chr9 65464093 N DEL 8
SRR1766450.1631028 chr9 65463442 N chr9 65463656 N DUP 7
SRR1766447.10630000 chr9 65463266 N chr9 65463447 N DEL 4
SRR1766481.7352772 chr9 65463267 N chr9 65463448 N DEL 3
SRR1766451.7435671 chr9 65463450 N chr9 65463840 N DUP 1
SRR1766465.5267955 chr9 65463526 N chr9 65463585 N DUP 11
SRR1766479.3744136 chr9 65463656 N chr9 65463906 N DEL 5
SRR1766485.7920916 chr9 65463483 N chr9 65463570 N DEL 5
SRR1766453.898781 chr9 65463680 N chr9 65463857 N DEL 1
SRR1766478.6011591 chr9 65463690 N chr9 65463867 N DEL 4
SRR1766473.2785009 chr9 65463249 N chr9 65463703 N DUP 3
SRR1766467.1318371 chr9 65463334 N chr9 65463696 N DUP 5
SRR1766442.33096789 chr9 65463315 N chr9 65463638 N DEL 5
SRR1766475.2784622 chr9 65463464 N chr9 65463794 N DUP 6
SRR1766450.6875658 chr9 65463583 N chr9 65463713 N DEL 5
SRR1766482.2786916 chr9 65463295 N chr9 65463807 N DEL 5
SRR1766454.3071092 chr9 65463141 N chr9 65463915 N DUP 1
SRR1766486.191736 chr9 65463576 N chr9 65463822 N DEL 14
SRR1766454.4912392 chr9 65463861 N chr9 65463931 N DUP 5
SRR1766459.6140402 chr9 65463361 N chr9 65463955 N DUP 9
SRR1766476.11307616 chr9 65463354 N chr9 65463948 N DUP 4
SRR1766443.9767953 chr9 65463946 N chr9 65464239 N DEL 2
SRR1766450.29170 chr9 65463959 N chr9 65464078 N DEL 15
SRR1766457.4708208 chr9 65463897 N chr9 65463967 N DUP 5
SRR1766478.689726 chr9 65463156 N chr9 65463859 N DEL 5
SRR1766445.4150389 chr9 65463966 N chr9 65464085 N DEL 11
SRR1766449.975507 chr9 65463462 N chr9 65463983 N DUP 10
SRR1766475.7491234 chr9 65463987 N chr9 65464280 N DEL 2
SRR1766480.5921802 chr9 65464053 N chr9 65464346 N DEL 2
SRR1766445.9632079 chr9 65464053 N chr9 65464346 N DEL 5
SRR1766459.7350213 chr9 65463969 N chr9 65464260 N DUP 5
SRR1766479.10458781 chr9 65464053 N chr9 65464346 N DEL 5
SRR1766442.6528827 chr9 65463142 N chr9 65464092 N DUP 2
SRR1766470.9058213 chr9 65463924 N chr9 65464013 N DEL 6
SRR1766481.8034749 chr9 65463429 N chr9 65464128 N DUP 5
SRR1766486.10829293 chr9 65463466 N chr9 65464163 N DUP 4
SRR1766448.6874688 chr9 65464163 N chr9 65464342 N DEL 12
SRR1766451.1854065 chr9 65463917 N chr9 65464152 N DUP 3
SRR1766486.3184930 chr9 65463834 N chr9 65464142 N DUP 6
SRR1766449.5077095 chr9 65464070 N chr9 65464361 N DUP 5
SRR1766486.10722375 chr9 65463365 N chr9 65464094 N DEL 5
SRR1766479.3744136 chr9 65463310 N chr9 65464099 N DEL 5
SRR1766445.550523 chr9 65463917 N chr9 65464208 N DUP 1
SRR1766469.2135139 chr9 65463591 N chr9 65464146 N DEL 10
SRR1766462.5534147 chr9 65463999 N chr9 65464232 N DUP 10
SRR1766486.915269 chr9 65463446 N chr9 65464147 N DEL 5
SRR1766461.7998064 chr9 65463964 N chr9 65464199 N DEL 10
SRR1766469.2342132 chr9 65463957 N chr9 65464192 N DEL 5
SRR1766447.3478055 chr9 65463198 N chr9 65464206 N DEL 6
SRR1766444.1004140 chr9 65463999 N chr9 65464292 N DEL 20
SRR1766442.10577646 chr9 65463854 N chr9 65464278 N DEL 5
SRR1766442.20079269 chr20 59428211 N chr20 59428338 N DUP 1
SRR1766465.4839687 chr20 59428182 N chr20 59428371 N DEL 3
SRR1766485.10528812 chr20 59428184 N chr20 59428373 N DEL 1
SRR1766467.1586799 chr20 59428216 N chr20 59428393 N DEL 2
SRR1766473.11131901 chr18 5307811 N chr18 5308006 N DUP 4
SRR1766469.4208441 chr18 5307811 N chr18 5308006 N DUP 2
SRR1766474.5992460 chr18 5307846 N chr18 5307991 N DUP 10
SRR1766482.12475002 chr18 5307846 N chr18 5307991 N DUP 10
SRR1766467.19534 chr18 5307846 N chr18 5307991 N DUP 10
SRR1766467.5165606 chr18 5307846 N chr18 5307991 N DUP 10
SRR1766468.6569986 chr18 5307864 N chr18 5307991 N DUP 13
SRR1766459.7245454 chr18 5307844 N chr18 5307899 N DEL 10
SRR1766457.7471719 chr18 5307846 N chr18 5307901 N DEL 10
SRR1766464.7261643 chr18 5307848 N chr18 5307903 N DEL 10
SRR1766451.6833976 chr18 5307858 N chr18 5307913 N DEL 9
SRR1766443.956066 chr18 5307851 N chr18 5307906 N DEL 8
SRR1766486.9586748 chr18 5307858 N chr18 5307913 N DEL 7
SRR1766450.5314766 chr18 5307858 N chr18 5307913 N DEL 6
SRR1766463.2698492 chr18 5307858 N chr18 5307913 N DEL 6
SRR1766448.3490131 chr18 5307858 N chr18 5307913 N DEL 1
SRR1766482.10645815 chr18 5307860 N chr18 5307915 N DEL 4
SRR1766483.9165522 chr18 5307857 N chr18 5307912 N DEL 2
SRR1766458.3819816 chr18 5307856 N chr18 5307911 N DEL 3
SRR1766469.7513519 chr13 45507938 N chr13 45508249 N DUP 1
SRR1766454.6268504 chr19 1335176 N chr19 1335294 N DEL 5
SRR1766479.2213449 chr19 1335176 N chr19 1335294 N DEL 7
SRR1766465.1469268 chr19 1335176 N chr19 1335294 N DEL 7
SRR1766465.9284207 chr19 1335193 N chr19 1335310 N DUP 2
SRR1766451.8485256 chr19 1335193 N chr19 1335310 N DUP 2
SRR1766459.10463865 chr19 1335193 N chr19 1335310 N DUP 7
SRR1766484.2450542 chr19 1335199 N chr19 1335316 N DUP 4
SRR1766465.1046633 chr19 1335228 N chr19 1335465 N DEL 8
SRR1766442.7950695 chr7 153099455 N chr7 153099592 N DUP 14
SRR1766472.5737061 chr7 153099506 N chr7 153099610 N DUP 8
SRR1766447.10125988 chr7 153099506 N chr7 153099610 N DUP 6
SRR1766463.556198 chr7 153099506 N chr7 153099610 N DUP 6
SRR1766463.8056104 chr7 153099506 N chr7 153099610 N DUP 4
SRR1766458.4748583 chr7 153099506 N chr7 153099610 N DUP 12
SRR1766477.10462747 chr7 153099506 N chr7 153099610 N DUP 19
SRR1766471.259 chr7 153099510 N chr7 153099581 N DEL 17
SRR1766473.4535927 chr7 153099510 N chr7 153099581 N DEL 17
SRR1766455.8674197 chr7 153099510 N chr7 153099581 N DEL 16
SRR1766465.7834250 chr7 153099477 N chr7 153099581 N DEL 10
SRR1766460.2375924 chr7 153099477 N chr7 153099581 N DEL 10
SRR1766442.35288392 chr7 153099477 N chr7 153099581 N DEL 7
SRR1766484.1426707 chr7 153099477 N chr7 153099581 N DEL 7
SRR1766443.4296107 chr7 153099478 N chr7 153099582 N DEL 6
SRR1766442.17799100 chr7 153099479 N chr7 153099583 N DEL 5
SRR1766453.1673370 chr7 153099468 N chr7 153099607 N DEL 5
SRR1766477.502888 chr7 153099469 N chr7 153099608 N DEL 4
SRR1766458.4748583 chr7 153099471 N chr7 153099610 N DEL 2
SRR1766462.2134386 chr7 153099472 N chr7 153099611 N DEL 1
SRR1766454.1291260 chr21 8108183 N chr21 8108318 N DUP 5
SRR1766483.10532728 chr21 8108183 N chr21 8108318 N DUP 5
SRR1766481.12544080 chr21 8108184 N chr21 8108319 N DUP 5
SRR1766470.5027380 chr19 40377188 N chr19 40377495 N DEL 6
SRR1766460.4998436 chr19 40377071 N chr19 40377273 N DUP 5
SRR1766454.4028571 chr19 40377443 N chr19 40377511 N DUP 30
SRR1766465.8063457 chr19 40377376 N chr19 40377618 N DEL 5
SRR1766475.9761562 chr12 130844007 N chr12 130844070 N DEL 5
SRR1766464.3274854 chr12 130844007 N chr12 130844070 N DEL 5
SRR1766473.6584017 chr12 130844007 N chr12 130844070 N DEL 5
SRR1766474.1468128 chr12 130844007 N chr12 130844070 N DEL 5
SRR1766475.3782027 chr12 130844007 N chr12 130844070 N DEL 5
SRR1766460.1525966 chr12 130844007 N chr12 130844070 N DEL 5
SRR1766468.3105777 chr12 130844007 N chr12 130844070 N DEL 5
SRR1766442.6322403 chr12 130843991 N chr12 130844094 N DEL 34
SRR1766457.8128979 chr12 130843976 N chr12 130844070 N DEL 5
SRR1766446.1126221 chr12 130843945 N chr12 130844070 N DEL 5
SRR1766449.5325254 chr12 130843995 N chr12 130844098 N DEL 8
SRR1766460.1390015 chr12 130843991 N chr12 130844094 N DEL 14
SRR1766465.2507526 chr12 130843971 N chr12 130844105 N DEL 4
SRR1766486.9030550 chr12 130843877 N chr12 130844249 N DUP 4
SRR1766448.1798010 chr18 72700626 N chr18 72700713 N DEL 1
SRR1766464.3691464 chr18 72700626 N chr18 72700713 N DEL 5
SRR1766454.2855140 chr18 72700626 N chr18 72700713 N DEL 4
SRR1766482.10739218 chr18 72700618 N chr18 72700673 N DEL 1
SRR1766442.29247993 chr18 72700618 N chr18 72700673 N DEL 1
SRR1766486.3970704 chr18 72700595 N chr18 72700674 N DEL 17
SRR1766474.2729783 chr18 72700593 N chr18 72700644 N DUP 13
SRR1766486.3837591 chr18 72700593 N chr18 72700644 N DUP 10
SRR1766486.8019183 chr18 72700585 N chr18 72700676 N DUP 17
SRR1766450.7661405 chr18 72700585 N chr18 72700676 N DUP 17
SRR1766442.7020145 chr18 72700585 N chr18 72700676 N DUP 21
SRR1766475.3957081 chr18 72700595 N chr18 72700646 N DUP 10
SRR1766442.30657527 chr18 72700585 N chr18 72700676 N DUP 25
SRR1766448.3275279 chr18 72700585 N chr18 72700676 N DUP 25
SRR1766444.4425999 chr18 72700607 N chr18 72700728 N DUP 11
SRR1766470.8099070 chr18 72700585 N chr18 72700676 N DUP 25
SRR1766458.6652782 chr18 72700607 N chr18 72700728 N DUP 14
SRR1766449.10167784 chr18 72700607 N chr18 72700728 N DUP 14
SRR1766452.3049058 chr18 72700607 N chr18 72700728 N DUP 14
SRR1766455.8822209 chr18 72700607 N chr18 72700728 N DUP 14
SRR1766449.9388123 chr18 72700642 N chr18 72700775 N DUP 8
SRR1766482.6669758 chr18 72700714 N chr18 72700779 N DEL 17
SRR1766447.1740189 chr18 72700585 N chr18 72700676 N DUP 33
SRR1766459.6422557 chr18 72700619 N chr18 72700686 N DUP 6
SRR1766460.4229383 chr18 72700619 N chr18 72700686 N DUP 7
SRR1766465.5830632 chr18 72700619 N chr18 72700686 N DUP 7
SRR1766486.11203849 chr18 72700660 N chr18 72700717 N DEL 12
SRR1766486.8736913 chr18 72700713 N chr18 72700768 N DUP 21
SRR1766458.8526070 chr18 72700723 N chr18 72700812 N DUP 11
SRR1766446.5312837 chr18 72700723 N chr18 72700802 N DUP 20
SRR1766452.9140727 chr18 72700723 N chr18 72700802 N DUP 18
SRR1766447.1653752 chr18 72700586 N chr18 72700689 N DEL 16
SRR1766471.9090486 chr18 72700723 N chr18 72700802 N DUP 20
SRR1766455.4383246 chr18 72700586 N chr18 72700689 N DEL 15
SRR1766456.2661636 chr18 72700679 N chr18 72700800 N DUP 14
SRR1766455.451742 chr18 72700717 N chr18 72700808 N DUP 16
SRR1766452.3235652 chr18 72700569 N chr18 72700798 N DUP 3
SRR1766452.7514105 chr18 72700609 N chr18 72700806 N DUP 10
SRR1766443.9552656 chr18 72700716 N chr18 72700827 N DUP 9
SRR1766477.8502443 chr18 72700688 N chr18 72700759 N DUP 16
SRR1766473.4480261 chr18 72700713 N chr18 72700768 N DUP 24
SRR1766442.12898108 chr18 72700569 N chr18 72700820 N DUP 10
SRR1766475.5339645 chr18 72700649 N chr18 72700824 N DUP 27
SRR1766448.1798010 chr18 72700638 N chr18 72700839 N DUP 15
SRR1766479.4542296 chr18 72700618 N chr18 72700837 N DUP 6
SRR1766445.8678055 chr18 72700733 N chr18 72700822 N DUP 7
SRR1766480.7812158 chr18 72700739 N chr18 72700846 N DUP 19
SRR1766460.4303843 chr18 72700713 N chr18 72700768 N DUP 18
SRR1766442.44724368 chr18 72700791 N chr18 72700854 N DEL 14
SRR1766455.9733843 chr18 72700791 N chr18 72700854 N DEL 15
SRR1766466.1964496 chr18 72700724 N chr18 72700779 N DEL 10
SRR1766463.2524836 chr18 72700698 N chr18 72700785 N DEL 11
SRR1766486.8019183 chr18 72700698 N chr18 72700785 N DEL 11
SRR1766454.10850453 chr18 72700798 N chr18 72700851 N DEL 20
SRR1766442.1681150 chr18 72700798 N chr18 72700851 N DEL 24
SRR1766474.8554568 chr18 72700798 N chr18 72700851 N DEL 24
SRR1766483.12153215 chr18 72700798 N chr18 72700851 N DEL 22
SRR1766477.7121867 chr18 72700798 N chr18 72700851 N DEL 21
SRR1766443.10371014 chr18 72700788 N chr18 72700851 N DEL 24
SRR1766477.10723407 chr18 72700788 N chr18 72700851 N DEL 23
SRR1766476.4863783 chr18 72700788 N chr18 72700851 N DEL 24
SRR1766467.4006965 chr18 72700799 N chr18 72700852 N DEL 21
SRR1766480.5171341 chr18 72700644 N chr18 72700807 N DEL 9
SRR1766452.3317249 chr18 72700645 N chr18 72700808 N DEL 9
SRR1766486.2793190 chr18 72700794 N chr18 72700857 N DEL 24
SRR1766448.9225421 chr18 72700672 N chr18 72700851 N DEL 20
SRR1766473.585183 chr18 72700727 N chr18 72700856 N DEL 22
SRR1766474.2729783 chr18 72700648 N chr18 72700837 N DEL 16
SRR1766460.9078900 chr18 72700752 N chr18 72700851 N DEL 22
SRR1766465.1660947 chr18 72700752 N chr18 72700851 N DEL 21
SRR1766442.25737276 chr18 72700752 N chr18 72700851 N DEL 14
SRR1766481.3362828 chr18 72700752 N chr18 72700851 N DEL 14
SRR1766476.10545279 chr18 72700638 N chr18 72700865 N DEL 8
SRR1766447.1740189 chr18 72700638 N chr18 72700865 N DEL 7
SRR1766463.9147906 chr18 72700714 N chr18 72700853 N DEL 8
SRR1766442.30511607 chr18 72700594 N chr18 72700875 N DEL 9
SRR1766454.2383869 chr18 72700594 N chr18 72700875 N DEL 9
SRR1766477.11752535 chr18 72700614 N chr18 72700881 N DEL 5
SRR1766463.6122822 chr18 72700616 N chr18 72700883 N DEL 5
SRR1766473.470257 chr18 72700617 N chr18 72700884 N DEL 5
SRR1766473.783508 chr18 72700617 N chr18 72700884 N DEL 5
SRR1766465.7040589 chr17 79009271 N chr17 79009428 N DEL 5
SRR1766444.5777634 chr2 219217455 N chr2 219217749 N DEL 24
SRR1766484.2983321 chr9 123972080 N chr9 123972265 N DUP 4
SRR1766450.1830161 chr9 123972236 N chr9 123972305 N DUP 5
SRR1766448.5937264 chr3 126480906 N chr3 126481047 N DUP 2
SRR1766450.3832692 chr4 113340843 N chr4 113340998 N DEL 12
SRR1766468.5266684 chr4 113340858 N chr4 113340998 N DEL 10
SRR1766479.10477188 chr13 104352717 N chr13 104352827 N DEL 5
SRR1766453.7864303 chr18 56600438 N chr18 56600643 N DEL 2
SRR1766482.9820345 chr18 56600438 N chr18 56600643 N DEL 2
SRR1766479.9645793 chr18 56600438 N chr18 56600643 N DEL 5
SRR1766477.9889776 chr18 56600438 N chr18 56600643 N DEL 5
SRR1766470.8593486 chr18 56600438 N chr18 56600643 N DEL 5
SRR1766466.10861152 chr18 56600438 N chr18 56600643 N DEL 5
SRR1766442.31217042 chr18 56600456 N chr18 56600729 N DEL 12
SRR1766442.41083980 chr18 56600477 N chr18 56600546 N DEL 5
SRR1766466.8081937 chr18 56600477 N chr18 56600750 N DEL 10
SRR1766468.1832756 chr18 56600524 N chr18 56600729 N DEL 5
SRR1766457.2333732 chr18 56600477 N chr18 56600546 N DEL 5
SRR1766464.10391499 chr18 56600592 N chr18 56600729 N DEL 5
SRR1766467.3765105 chr18 56600490 N chr18 56600559 N DEL 2
SRR1766482.3069028 chr18 56600477 N chr18 56600682 N DEL 12
SRR1766466.10075382 chr18 56600477 N chr18 56600682 N DEL 5
SRR1766463.5474017 chr18 56600456 N chr18 56600729 N DEL 10
SRR1766442.40438631 chr18 56600483 N chr18 56600756 N DEL 4
SRR1766471.9599803 chr18 56600490 N chr18 56600763 N DEL 2
SRR1766446.1359248 chr13 112913059 N chr13 112913114 N DEL 2
SRR1766468.2214364 chr13 112913096 N chr13 112913290 N DEL 16
SRR1766482.1615913 chr13 112912925 N chr13 112913136 N DUP 10
SRR1766485.1254717 chr13 112912925 N chr13 112913136 N DUP 10
SRR1766454.9352715 chr13 112913046 N chr13 112913472 N DUP 2
SRR1766444.937925 chr13 112913168 N chr13 112913367 N DEL 26
SRR1766469.6957938 chr13 112913171 N chr13 112913417 N DUP 5
SRR1766468.1245468 chr13 112913196 N chr13 112913485 N DUP 13
SRR1766460.9256776 chr13 112913023 N chr13 112913319 N DUP 9
SRR1766465.580634 chr13 112913023 N chr13 112913319 N DUP 9
SRR1766459.3967336 chr13 112913319 N chr13 112913376 N DEL 9
SRR1766442.21004947 chr13 112913230 N chr13 112913441 N DUP 12
SRR1766445.9258250 chr13 112913319 N chr13 112913376 N DEL 9
SRR1766471.10374421 chr13 112913319 N chr13 112913376 N DEL 9
SRR1766477.11772392 chr13 112913030 N chr13 112913230 N DEL 10
SRR1766478.4786746 chr13 112912940 N chr13 112913261 N DEL 10
SRR1766464.9335565 chr13 112913037 N chr13 112913285 N DEL 5
SRR1766469.2555346 chr13 112913333 N chr13 112913440 N DUP 5
SRR1766479.5159318 chr13 112912952 N chr13 112913412 N DEL 1
SRR1766467.7379286 chrX 2478754 N chrX 2478843 N DEL 5
SRR1766472.1862328 chrX 2478837 N chrX 2479035 N DUP 10
SRR1766481.8035858 chrX 2479253 N chrX 2480015 N DEL 5
SRR1766459.2464684 chrX 2478778 N chrX 2479517 N DUP 5
SRR1766466.6429593 chrX 2479502 N chrX 2479824 N DEL 10
SRR1766479.10144879 chrX 2479510 N chrX 2479832 N DEL 4
SRR1766455.6917523 chrX 2479453 N chrX 2479773 N DUP 5
SRR1766483.6659664 chrX 2479341 N chrX 2479494 N DEL 5
SRR1766477.4567019 chrX 2479489 N chrX 2479811 N DEL 5
SRR1766467.372297 chrX 2479508 N chrX 2479830 N DEL 15
SRR1766442.11822571 chr1 191824847 N chr1 191824945 N DUP 6
SRR1766447.6647937 chr1 191824847 N chr1 191824945 N DUP 6
SRR1766449.9297277 chr1 191824863 N chr1 191824961 N DEL 1
SRR1766446.3714889 chr2 883725 N chr2 883911 N DEL 5
SRR1766485.8998984 chr2 883725 N chr2 883911 N DEL 5
SRR1766442.41055716 chr2 883800 N chr2 883949 N DEL 4
SRR1766450.7217391 chr1 4332501 N chr1 4332995 N DEL 5
SRR1766445.783593 chr1 4332511 N chr1 4332570 N DEL 5
SRR1766476.4598130 chr1 4332511 N chr1 4332570 N DEL 5
SRR1766456.2953573 chr1 4332511 N chr1 4332570 N DEL 9
SRR1766474.4875424 chr1 4332511 N chr1 4332570 N DEL 10
SRR1766485.7883323 chr1 4332511 N chr1 4332570 N DEL 10
SRR1766443.2662307 chr1 4332502 N chr1 4333170 N DEL 5
SRR1766471.1229517 chr1 4332511 N chr1 4332570 N DEL 17
SRR1766447.2595331 chr1 4332511 N chr1 4332570 N DEL 19
SRR1766452.5371918 chr1 4332502 N chr1 4332590 N DEL 20
SRR1766479.6270613 chr1 4332515 N chr1 4333359 N DEL 5
SRR1766471.6661709 chr1 4332511 N chr1 4332570 N DEL 10
SRR1766442.25037148 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766480.789992 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766483.8087285 chr1 4332556 N chr1 4333518 N DEL 16
SRR1766469.1790376 chr1 4332556 N chr1 4332992 N DEL 22
SRR1766471.256383 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766465.10568007 chr1 4332511 N chr1 4332918 N DEL 15
SRR1766443.3753855 chr1 4332556 N chr1 4333518 N DEL 20
SRR1766471.8142180 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766450.6375570 chr1 4332511 N chr1 4332570 N DEL 20
SRR1766478.7511124 chr1 4332511 N chr1 4332570 N DEL 10
SRR1766454.9133928 chr1 4332614 N chr1 4333427 N DUP 10
SRR1766443.11094727 chr1 4332570 N chr1 4332627 N DUP 15
SRR1766479.12282309 chr1 4332511 N chr1 4332570 N DEL 12
SRR1766452.3110424 chr1 4332523 N chr1 4332582 N DEL 3
SRR1766467.5353285 chr1 4332523 N chr1 4332582 N DEL 3
SRR1766466.3535845 chr1 4332690 N chr1 4332777 N DEL 13
SRR1766448.9216519 chr1 4332529 N chr1 4332588 N DEL 5
SRR1766462.4078557 chr1 4332645 N chr1 4332936 N DEL 10
SRR1766477.3445356 chr1 4332536 N chr1 4332595 N DEL 5
SRR1766476.6614264 chr1 4332701 N chr1 4333576 N DEL 5
SRR1766482.9931920 chr1 4332729 N chr1 4333136 N DEL 6
SRR1766449.3611427 chr1 4332615 N chr1 4332991 N DUP 11
SRR1766478.828829 chr1 4332671 N chr1 4333517 N DEL 14
SRR1766485.2259402 chr1 4332570 N chr1 4332627 N DUP 10
SRR1766456.2953573 chr1 4332614 N chr1 4333048 N DUP 10
SRR1766467.849919 chr1 4333225 N chr1 4333491 N DEL 8
SRR1766470.8163488 chr1 4332614 N chr1 4332758 N DUP 5
SRR1766471.256383 chr1 4332570 N chr1 4332685 N DUP 5
SRR1766471.6661709 chr1 4332599 N chr1 4332743 N DUP 5
SRR1766481.8647723 chr1 4332592 N chr1 4332823 N DUP 5
SRR1766474.4875424 chr1 4332526 N chr1 4332614 N DEL 5
SRR1766472.7361104 chr1 4332520 N chr1 4332607 N DEL 7
SRR1766476.6614264 chr1 4332700 N chr1 4333194 N DEL 5
SRR1766471.1229517 chr1 4332614 N chr1 4332990 N DUP 10
SRR1766448.9216519 chr1 4332743 N chr1 4332976 N DEL 10
SRR1766443.9513170 chr1 4332570 N chr1 4332714 N DUP 5
SRR1766460.5584371 chr1 4332700 N chr1 4333194 N DEL 10
SRR1766447.1486885 chr1 4332686 N chr1 4332743 N DUP 5
SRR1766449.2220687 chr1 4332681 N chr1 4333088 N DEL 8
SRR1766464.1642681 chr1 4333001 N chr1 4333584 N DUP 10
SRR1766481.11062883 chr1 4332535 N chr1 4333582 N DUP 2
SRR1766463.8403608 chr1 4332614 N chr1 4333576 N DEL 10
SRR1766450.2795016 chr1 4333020 N chr1 4333489 N DEL 15
SRR1766459.7560099 chr1 4333049 N chr1 4333371 N DEL 10
SRR1766460.4685531 chr1 4332532 N chr1 4332997 N DEL 5
SRR1766444.5549244 chr1 4333240 N chr1 4333448 N DEL 10
SRR1766453.2633158 chr1 4333066 N chr1 4333359 N DEL 5
SRR1766443.2989947 chr1 4333182 N chr1 4333448 N DEL 10
SRR1766465.7261728 chr1 4332556 N chr1 4333460 N DEL 10
SRR1766462.9770067 chr1 4333053 N chr1 4333112 N DEL 6
SRR1766460.2024603 chr1 4332962 N chr1 4333077 N DUP 5
SRR1766454.10890745 chr1 4333054 N chr1 4333523 N DEL 10
SRR1766479.6270613 chr1 4333021 N chr1 4333575 N DUP 15
SRR1766484.9888651 chr1 4332515 N chr1 4333448 N DEL 15
SRR1766443.2989947 chr1 4332533 N chr1 4333085 N DEL 5
SRR1766485.286538 chr1 4332520 N chr1 4333453 N DEL 5
SRR1766442.34626457 chr1 4332533 N chr1 4333085 N DEL 5
SRR1766448.1485734 chr1 4332565 N chr1 4333146 N DEL 10
SRR1766478.5981531 chr1 4332545 N chr1 4333097 N DEL 3
SRR1766473.11281022 chr1 4333252 N chr1 4333489 N DEL 9
SRR1766472.7361104 chr1 4332631 N chr1 4333448 N DEL 12
SRR1766484.1814950 chr1 4333124 N chr1 4333448 N DEL 5
SRR1766486.5451510 chr1 4332936 N chr1 4333167 N DUP 15
SRR1766442.16759186 chr1 4332527 N chr1 4333108 N DEL 5
SRR1766444.2797920 chr1 4333112 N chr1 4333256 N DUP 10
SRR1766470.9585706 chr1 4332614 N chr1 4333108 N DEL 10
SRR1766474.1748250 chr1 4332556 N chr1 4333460 N DEL 5
SRR1766463.4639370 chr1 4333165 N chr1 4333489 N DEL 5
SRR1766483.4148876 chr1 4333053 N chr1 4333112 N DEL 5
SRR1766472.10639638 chr1 4333133 N chr1 4333457 N DEL 10
SRR1766442.8407769 chr1 4332874 N chr1 4333136 N DEL 5
SRR1766466.6107027 chr1 4332562 N chr1 4333085 N DEL 10
SRR1766474.1894881 chr1 4332556 N chr1 4333137 N DEL 10
SRR1766475.9062244 chr1 4333053 N chr1 4333609 N DEL 9
SRR1766466.10153244 chr1 4332642 N chr1 4333136 N DEL 12
SRR1766467.849919 chr1 4333166 N chr1 4333310 N DUP 10
SRR1766471.1670898 chr1 4333085 N chr1 4333142 N DUP 5
SRR1766464.5114633 chr1 4333053 N chr1 4333141 N DEL 12
SRR1766472.9786426 chr1 4333037 N chr1 4333448 N DEL 5
SRR1766450.2795016 chr1 4333170 N chr1 4333550 N DUP 5
SRR1766470.9585706 chr1 4332652 N chr1 4333175 N DEL 6
SRR1766449.8726051 chr1 4333066 N chr1 4333448 N DEL 5
SRR1766467.1043592 chr1 4333053 N chr1 4333493 N DEL 12
SRR1766460.10628435 chr1 4332556 N chr1 4333166 N DEL 5
SRR1766442.32457730 chr1 4332614 N chr1 4333222 N DUP 10
SRR1766459.7560099 chr1 4332590 N chr1 4333169 N DUP 10
SRR1766481.10704111 chr1 4332566 N chr1 4333147 N DEL 5
SRR1766481.11062883 chr1 4332590 N chr1 4333169 N DUP 10
SRR1766442.16313221 chr1 4332502 N chr1 4333226 N DUP 10
SRR1766462.1269920 chr1 4332560 N chr1 4333170 N DEL 10
SRR1766471.1038908 chr1 4333252 N chr1 4333489 N DEL 10
SRR1766474.1894881 chr1 4333170 N chr1 4333227 N DUP 5
SRR1766469.3524751 chr1 4333066 N chr1 4333359 N DEL 10
SRR1766449.8726051 chr1 4333252 N chr1 4333489 N DEL 10
SRR1766466.3741585 chr1 4333223 N chr1 4333489 N DEL 10
SRR1766481.3825966 chr1 4333240 N chr1 4333448 N DEL 10
SRR1766450.792823 chr1 4333085 N chr1 4333229 N DUP 10
SRR1766442.20683542 chr1 4332560 N chr1 4333170 N DEL 10
SRR1766461.10140590 chr1 4333002 N chr1 4333119 N DEL 4
SRR1766442.16313221 chr1 4333170 N chr1 4333227 N DUP 5
SRR1766476.5789993 chr1 4333024 N chr1 4333170 N DEL 5
SRR1766483.11597062 chr1 4332992 N chr1 4333165 N DUP 10
SRR1766477.6080896 chr1 4332531 N chr1 4333170 N DEL 5
SRR1766455.6174278 chr1 4332671 N chr1 4333223 N DEL 20
SRR1766483.8250848 chr1 4333228 N chr1 4333285 N DUP 10
SRR1766444.3208028 chr1 4332992 N chr1 4333194 N DUP 5
SRR1766483.8250848 chr1 4332595 N chr1 4333176 N DEL 9
SRR1766469.8345969 chr1 4333223 N chr1 4333489 N DEL 10
SRR1766455.8779410 chr1 4333057 N chr1 4333232 N DEL 5
SRR1766478.11806826 chr1 4333252 N chr1 4333634 N DEL 5
SRR1766452.9231973 chr1 4333252 N chr1 4333634 N DEL 5
SRR1766447.620163 chr1 4333165 N chr1 4333489 N DEL 6
SRR1766458.7649016 chr1 4333049 N chr1 4333371 N DEL 10
SRR1766452.9231973 chr1 4332555 N chr1 4333604 N DEL 5
SRR1766454.4261401 chr1 4333256 N chr1 4333522 N DEL 5
SRR1766469.677256 chr1 4332555 N chr1 4333604 N DEL 10
SRR1766442.13032733 chr1 4333169 N chr1 4333228 N DEL 5
SRR1766465.3335790 chr1 4333252 N chr1 4333634 N DEL 5
SRR1766474.8228594 chr1 4332538 N chr1 4333349 N DUP 7
SRR1766442.37408697 chr1 4333217 N chr1 4333361 N DUP 5
SRR1766483.7481342 chr1 4333169 N chr1 4333493 N DEL 10
SRR1766442.8407769 chr1 4333240 N chr1 4333359 N DEL 10
SRR1766467.1043592 chr1 4333275 N chr1 4333361 N DUP 5
SRR1766464.5741593 chr1 4333285 N chr1 4333464 N DEL 12
SRR1766442.34375501 chr1 4333053 N chr1 4333464 N DEL 14
SRR1766445.186957 chr1 4333021 N chr1 4333399 N DUP 5
SRR1766468.3127432 chr1 4333135 N chr1 4333397 N DUP 5
SRR1766458.5654430 chr1 4333289 N chr1 4333553 N DUP 2
SRR1766461.7475944 chr1 4332528 N chr1 4333575 N DUP 4
SRR1766459.2363648 chr1 4332564 N chr1 4333613 N DEL 5
SRR1766453.10705774 chr1 4333358 N chr1 4333415 N DUP 5
SRR1766442.46233639 chr1 4333227 N chr1 4333433 N DEL 10
SRR1766442.46233639 chr1 4332531 N chr1 4333433 N DEL 5
SRR1766468.1790849 chr1 4333182 N chr1 4333448 N DEL 7
SRR1766455.9480667 chr1 4332556 N chr1 4333460 N DEL 8
SRR1766443.3753855 chr1 4332564 N chr1 4333468 N DEL 12
SRR1766467.9049772 chr1 4333326 N chr1 4333447 N DEL 12
SRR1766485.286538 chr1 4332564 N chr1 4333468 N DEL 12
SRR1766474.7774313 chr1 4333136 N chr1 4333489 N DEL 10
SRR1766442.33298095 chr1 4332557 N chr1 4333461 N DEL 7
SRR1766442.43738499 chr1 4332556 N chr1 4333021 N DEL 5
SRR1766449.7436817 chr1 4333053 N chr1 4333493 N DEL 7
SRR1766459.3730973 chr1 4332615 N chr1 4333461 N DEL 7
SRR1766466.10153244 chr1 4332642 N chr1 4333136 N DEL 15
SRR1766478.4413525 chr1 4332502 N chr1 4333255 N DUP 10
SRR1766479.4063835 chr1 4332561 N chr1 4333465 N DEL 5
SRR1766463.4639370 chr1 4332614 N chr1 4333545 N DUP 5
SRR1766459.2363648 chr1 4332563 N chr1 4333086 N DEL 5
SRR1766466.3741585 chr1 4332875 N chr1 4333489 N DEL 10
SRR1766450.2510119 chr1 4333136 N chr1 4333489 N DEL 10
SRR1766445.9931266 chr1 4333240 N chr1 4333448 N DEL 6
SRR1766445.9931266 chr1 4333428 N chr1 4333489 N DEL 7
SRR1766480.5203697 chr1 4332963 N chr1 4333575 N DUP 2
SRR1766453.3374479 chr1 4332512 N chr1 4333120 N DUP 2
SRR1766469.8345969 chr1 4332540 N chr1 4333121 N DEL 2
SRR1766446.9867708 chr1 4333428 N chr1 4333489 N DEL 6
SRR1766442.38347614 chr1 4332600 N chr1 4333065 N DEL 4
SRR1766473.3704186 chr1 4332555 N chr1 4332614 N DEL 5
SRR1766473.3704186 chr1 4332614 N chr1 4333545 N DUP 10
SRR1766457.4261973 chr1 4333153 N chr1 4333448 N DEL 5
SRR1766481.12841215 chr1 4332874 N chr1 4333459 N DEL 15
SRR1766465.2185972 chr1 4332562 N chr1 4333085 N DEL 10
SRR1766480.5203697 chr1 4333165 N chr1 4333489 N DEL 5
SRR1766479.6994666 chr1 4333053 N chr1 4333522 N DEL 10
SRR1766447.620163 chr1 4333240 N chr1 4333448 N DEL 10
SRR1766458.7649016 chr1 4333136 N chr1 4333576 N DEL 5
SRR1766447.2251398 chr1 4333090 N chr1 4333731 N DUP 10
SRR1766480.8000657 chr1 4332874 N chr1 4333517 N DEL 10
SRR1766465.2185972 chr1 4333078 N chr1 4333489 N DEL 10
SRR1766467.9049772 chr1 4333547 N chr1 4333691 N DUP 10
SRR1766481.6779784 chr1 4333092 N chr1 4333588 N DUP 10
SRR1766469.3524751 chr1 4333124 N chr1 4333448 N DEL 5
SRR1766447.5845708 chr1 4333136 N chr1 4333460 N DEL 5
SRR1766465.7261728 chr1 4333371 N chr1 4333575 N DUP 10
SRR1766463.4878448 chr1 4332553 N chr1 4333515 N DEL 3
SRR1766482.2700706 chr1 4332541 N chr1 4333503 N DEL 1
SRR1766479.1262570 chr1 4332541 N chr1 4333503 N DEL 1
SRR1766459.6990454 chr1 4333020 N chr1 4333108 N DEL 1
SRR1766442.41634223 chr1 4332642 N chr1 4333517 N DEL 5
SRR1766481.7225112 chr1 4332992 N chr1 4333575 N DUP 6
SRR1766442.38347614 chr1 4333179 N chr1 4333503 N DEL 5
SRR1766483.4148876 chr1 4333166 N chr1 4333575 N DUP 12
SRR1766479.2559879 chr1 4332879 N chr1 4333493 N DEL 10
SRR1766465.5208960 chr1 4332544 N chr1 4333448 N DEL 10
SRR1766446.4553163 chr1 4333460 N chr1 4333575 N DUP 5
SRR1766446.8172668 chr1 4332613 N chr1 4333517 N DEL 5
SRR1766455.346619 chr1 4333053 N chr1 4333522 N DEL 10
SRR1766472.1021449 chr1 4333518 N chr1 4333575 N DUP 5
SRR1766455.9480667 chr1 4332556 N chr1 4333518 N DEL 5
SRR1766479.1262570 chr1 4333460 N chr1 4333575 N DUP 5
SRR1766459.3730973 chr1 4332544 N chr1 4333448 N DEL 5
SRR1766458.7629482 chr1 4333460 N chr1 4333575 N DUP 10
SRR1766469.10592314 chr1 4333371 N chr1 4333575 N DUP 10
SRR1766474.8228594 chr1 4332999 N chr1 4333172 N DUP 10
SRR1766483.4585195 chr1 4332622 N chr1 4333468 N DEL 5
SRR1766482.1670418 chr1 4332544 N chr1 4333448 N DEL 10
SRR1766449.1687719 chr1 4333310 N chr1 4333460 N DEL 15
SRR1766484.3692511 chr1 4333170 N chr1 4333579 N DUP 10
SRR1766460.9406510 chr1 4332556 N chr1 4332963 N DEL 20
SRR1766468.4864345 chr1 4332875 N chr1 4333576 N DEL 10
SRR1766442.40835555 chr1 4332556 N chr1 4333460 N DEL 4
SRR1766442.4939146 chr1 4332598 N chr1 4333473 N DEL 8
SRR1766474.670863 chr1 4332556 N chr1 4333460 N DEL 10
SRR1766465.9274606 chr1 4332560 N chr1 4333170 N DEL 10
SRR1766458.7629482 chr1 4332556 N chr1 4333460 N DEL 10
SRR1766459.6990454 chr1 4332562 N chr1 4333553 N DEL 5
SRR1766486.5451510 chr1 4332943 N chr1 4333174 N DUP 5
SRR1766471.1670898 chr1 4332562 N chr1 4333085 N DEL 9
SRR1766481.12841215 chr1 4333020 N chr1 4333576 N DEL 5
SRR1766484.4761812 chr1 4333048 N chr1 4333604 N DEL 10
SRR1766442.33298095 chr1 4333518 N chr1 4333633 N DUP 5
SRR1766442.43738499 chr1 4333048 N chr1 4333604 N DEL 10
SRR1766476.9274028 chr1 4332618 N chr1 4333257 N DEL 5
SRR1766453.5992314 chr1 4332560 N chr1 4333609 N DEL 5
SRR1766444.1054712 chr1 4332556 N chr1 4333460 N DEL 10
SRR1766442.40835555 chr1 4333488 N chr1 4333603 N DUP 5
SRR1766454.10890745 chr1 4333053 N chr1 4333141 N DEL 15
SRR1766486.10288154 chr1 4333140 N chr1 4333667 N DEL 5
SRR1766448.6090716 chr1 4333140 N chr1 4333667 N DEL 5
SRR1766485.2358435 chr1 4333227 N chr1 4333667 N DEL 6
SRR1766450.8707403 chr1 4332552 N chr1 4333717 N DEL 5
SRR1766467.11823516 chr20 39587209 N chr20 39587258 N DUP 7
SRR1766462.8971630 chr20 39587209 N chr20 39587258 N DUP 13
SRR1766461.3632346 chr20 39587214 N chr20 39587263 N DUP 7
SRR1766457.4544417 chr20 39587209 N chr20 39587258 N DUP 16
SRR1766468.154946 chr2 16394934 N chr2 16395048 N DEL 11
SRR1766443.1433892 chr2 16394776 N chr2 16395021 N DUP 1
SRR1766475.2546903 chr2 16394879 N chr2 16395028 N DUP 5
SRR1766477.6539397 chr2 16394881 N chr2 16395065 N DUP 3
SRR1766482.5551912 chr16 30168670 N chr16 30168827 N DEL 1
SRR1766478.3064759 chr16 30168723 N chr16 30168880 N DEL 9
SRR1766472.3984521 chr16 30168723 N chr16 30168880 N DEL 12
SRR1766455.543757 chr16 30168726 N chr16 30168883 N DEL 5
SRR1766469.1566859 chr1 240562926 N chr1 240563269 N DEL 5
SRR1766454.8041988 chr1 240562858 N chr1 240563056 N DUP 17
SRR1766468.7033252 chr1 240562859 N chr1 240563099 N DUP 10
SRR1766479.6932056 chr1 240562858 N chr1 240563108 N DUP 6
SRR1766456.5164934 chr1 240563111 N chr1 240563249 N DEL 5
SRR1766466.8439118 chr1 240562859 N chr1 240563115 N DUP 16
SRR1766468.4875062 chr1 240563121 N chr1 240563285 N DEL 15
SRR1766459.8035047 chr1 240563111 N chr1 240563293 N DUP 5
SRR1766468.352914 chr1 240562954 N chr1 240563160 N DEL 5
SRR1766483.6409062 chr1 240562883 N chr1 240563169 N DEL 3
SRR1766476.1165897 chr1 240562959 N chr1 240563220 N DEL 1
SRR1766458.7703655 chr1 240562882 N chr1 240563235 N DEL 15
SRR1766453.912378 chr1 240562873 N chr1 240563318 N DEL 11
SRR1766447.4676141 chr1 1971362 N chr1 1971465 N DUP 1
SRR1766446.2314478 chr5 2082060 N chr5 2082754 N DEL 10
SRR1766464.834586 chr5 2082074 N chr5 2082201 N DEL 5
SRR1766461.5392737 chr5 2082124 N chr5 2082692 N DEL 5
SRR1766443.8121442 chr5 2082119 N chr5 2082246 N DEL 3
SRR1766476.8349894 chr5 2082074 N chr5 2082201 N DEL 3
SRR1766455.148065 chr5 2082133 N chr5 2082197 N DEL 5
SRR1766442.15028508 chr5 2082122 N chr5 2082249 N DEL 5
SRR1766458.1347836 chr5 2082119 N chr5 2082750 N DEL 5
SRR1766460.973177 chr5 2082097 N chr5 2082728 N DEL 5
SRR1766459.1812272 chr5 2082119 N chr5 2082750 N DEL 5
SRR1766476.5724190 chr5 2082097 N chr5 2082350 N DEL 10
SRR1766478.10028038 chr5 2082132 N chr5 2082196 N DEL 5
SRR1766460.4549354 chr5 2082119 N chr5 2082624 N DEL 5
SRR1766462.2130872 chr5 2082119 N chr5 2082624 N DEL 5
SRR1766469.9201828 chr5 2082160 N chr5 2082665 N DEL 5
SRR1766465.9617330 chr5 2082132 N chr5 2082196 N DEL 15
SRR1766466.6979812 chr5 2082119 N chr5 2082624 N DEL 5
SRR1766451.2121864 chr5 2082182 N chr5 2082750 N DEL 10
SRR1766454.1259899 chr5 2082132 N chr5 2082196 N DEL 10
SRR1766466.7929962 chr5 2082212 N chr5 2082906 N DEL 5
SRR1766452.7887974 chr5 2082212 N chr5 2082906 N DEL 5
SRR1766460.4549354 chr5 2082112 N chr5 2082174 N DUP 3
SRR1766453.6838218 chr5 2082191 N chr5 2082255 N DEL 10
SRR1766459.7030901 chr5 2082166 N chr5 2082354 N DUP 5
SRR1766473.3659979 chr5 2082245 N chr5 2082750 N DEL 5
SRR1766461.9627156 chr5 2082245 N chr5 2082750 N DEL 5
SRR1766451.9412735 chr5 2082245 N chr5 2082750 N DEL 5
SRR1766459.8540435 chr5 2082249 N chr5 2082754 N DEL 5
SRR1766472.11871052 chr5 2082196 N chr5 2082258 N DUP 10
SRR1766467.6948079 chr5 2082192 N chr5 2082254 N DUP 5
SRR1766442.36890550 chr5 2082196 N chr5 2082258 N DUP 5
SRR1766484.1156189 chr5 2082196 N chr5 2082447 N DUP 9
SRR1766453.704886 chr5 2082196 N chr5 2082951 N DUP 20
SRR1766456.182501 chr5 2082197 N chr5 2082385 N DUP 11
SRR1766446.2080380 chr5 2082201 N chr5 2082704 N DUP 5
SRR1766443.1616175 chr5 2082209 N chr5 2082964 N DUP 16
SRR1766469.5317302 chr5 2082227 N chr5 2082478 N DUP 10
SRR1766478.6279524 chr5 2082196 N chr5 2082258 N DUP 5
SRR1766481.1004632 chr5 2082250 N chr5 2082879 N DUP 10
SRR1766484.8580938 chr5 2082196 N chr5 2082258 N DUP 5
SRR1766455.4480380 chr5 2082142 N chr5 2082206 N DEL 5
SRR1766483.10367560 chr5 2082211 N chr5 2082966 N DUP 7
SRR1766476.8382786 chr5 2082212 N chr5 2082967 N DUP 6
SRR1766459.5443341 chr5 2082209 N chr5 2082964 N DUP 10
SRR1766450.5480536 chr5 2082209 N chr5 2082964 N DUP 12
SRR1766466.7925634 chr5 2082209 N chr5 2082964 N DUP 9
SRR1766481.11384315 chr5 2082161 N chr5 2082286 N DUP 10
SRR1766446.1595698 chr5 2082196 N chr5 2082258 N DUP 5
SRR1766475.6634289 chr5 2082209 N chr5 2082964 N DUP 10
SRR1766446.4595964 chr5 2082100 N chr5 2082227 N DEL 5
SRR1766469.10290856 chr5 2082196 N chr5 2082258 N DUP 7
SRR1766460.842661 chr5 2082228 N chr5 2082920 N DUP 5
SRR1766469.8755837 chr5 2082229 N chr5 2082921 N DUP 5
SRR1766484.4042638 chr5 2082232 N chr5 2082924 N DUP 5
SRR1766481.1004632 chr5 2082236 N chr5 2082928 N DUP 2
SRR1766450.954317 chr5 2082237 N chr5 2082929 N DUP 1
SRR1766450.1585522 chr5 2082032 N chr5 2082346 N DUP 1
SRR1766469.964652 chr5 2082032 N chr5 2082346 N DUP 1
SRR1766450.5453203 chr5 2082308 N chr5 2082750 N DEL 10
SRR1766483.8801681 chr5 2082164 N chr5 2082352 N DUP 5
SRR1766473.3085682 chr5 2082227 N chr5 2082352 N DUP 5
SRR1766468.3596826 chr5 2082251 N chr5 2082376 N DUP 5
SRR1766450.7750657 chr5 2082227 N chr5 2082352 N DUP 5
SRR1766481.8880086 chr5 2082227 N chr5 2082352 N DUP 5
SRR1766475.6634289 chr5 2082227 N chr5 2082478 N DUP 10
SRR1766481.7799500 chr5 2082227 N chr5 2082352 N DUP 5
SRR1766477.3744741 chr5 2082227 N chr5 2082352 N DUP 5
SRR1766469.8755837 chr5 2082290 N chr5 2082352 N DUP 5
SRR1766459.6845459 chr5 2082287 N chr5 2082790 N DUP 5
SRR1766465.4384166 chr5 2082287 N chr5 2082790 N DUP 5
SRR1766466.5686427 chr5 2082227 N chr5 2082352 N DUP 5
SRR1766473.5306008 chr5 2082196 N chr5 2082321 N DUP 5
SRR1766482.9760780 chr5 2082227 N chr5 2082352 N DUP 5
SRR1766468.3596826 chr5 2082223 N chr5 2082287 N DEL 5
SRR1766482.10649015 chr5 2082290 N chr5 2082352 N DUP 5
SRR1766451.9412735 chr5 2082258 N chr5 2082700 N DEL 6
SRR1766450.9142505 chr5 2082290 N chr5 2082352 N DUP 8
SRR1766469.8761440 chr5 2082227 N chr5 2082352 N DUP 5
SRR1766466.6979812 chr5 2082098 N chr5 2082288 N DEL 5
SRR1766460.1427802 chr5 2082290 N chr5 2082352 N DUP 5
SRR1766458.8142029 chr5 2082293 N chr5 2082355 N DUP 5
SRR1766459.4591209 chr5 2082294 N chr5 2082356 N DUP 5
SRR1766453.5955092 chr5 2082169 N chr5 2082296 N DEL 5
SRR1766458.1347836 chr5 2082291 N chr5 2082353 N DUP 9
SRR1766467.8752444 chr5 2082173 N chr5 2082300 N DEL 2
SRR1766480.5386032 chr5 2082196 N chr5 2082384 N DUP 5
SRR1766450.1104214 chr5 2082380 N chr5 2082822 N DEL 5
SRR1766482.875934 chr5 2082380 N chr5 2082822 N DEL 5
SRR1766477.11119298 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766463.2581591 chr5 2082075 N chr5 2082452 N DUP 3
SRR1766444.3096530 chr5 2082164 N chr5 2082352 N DUP 10
SRR1766449.7154566 chr5 2082196 N chr5 2082447 N DUP 5
SRR1766468.4036633 chr5 2082075 N chr5 2082452 N DUP 5
SRR1766453.3350555 chr5 2082196 N chr5 2082447 N DUP 10
SRR1766477.11550512 chr5 2082227 N chr5 2082478 N DUP 10
SRR1766442.22977030 chr5 2082227 N chr5 2082478 N DUP 15
SRR1766444.669476 chr5 2082249 N chr5 2082500 N DUP 5
SRR1766469.5618666 chr5 2082350 N chr5 2082475 N DUP 10
SRR1766445.9402365 chr5 2082061 N chr5 2082438 N DUP 5
SRR1766442.537461 chr5 2082311 N chr5 2082438 N DEL 5
SRR1766470.6372347 chr5 2082075 N chr5 2082263 N DUP 13
SRR1766442.30431816 chr5 2082061 N chr5 2082438 N DUP 5
SRR1766474.531252 chr5 2082196 N chr5 2082510 N DUP 3
SRR1766485.8949923 chr5 2082075 N chr5 2082452 N DUP 5
SRR1766445.10020896 chr5 2082500 N chr5 2082627 N DEL 5
SRR1766458.9248811 chr5 2082196 N chr5 2082510 N DUP 4
SRR1766456.3171398 chr5 2082077 N chr5 2082454 N DUP 5
SRR1766482.9383632 chr5 2082104 N chr5 2082355 N DUP 9
SRR1766449.2189563 chr5 2082209 N chr5 2082964 N DUP 34
SRR1766442.34745321 chr5 2082152 N chr5 2082216 N DEL 5
SRR1766459.10980685 chr5 2082196 N chr5 2082447 N DUP 20
SRR1766453.3543145 chr5 2082192 N chr5 2082254 N DUP 10
SRR1766484.1156189 chr5 2082209 N chr5 2082964 N DUP 20
SRR1766478.1860006 chr5 2082209 N chr5 2082964 N DUP 30
SRR1766450.2008726 chr5 2082209 N chr5 2082964 N DUP 30
SRR1766459.1812272 chr5 2082172 N chr5 2082297 N DUP 4
SRR1766443.610151 chr5 2082209 N chr5 2082964 N DUP 22
SRR1766485.4625684 chr5 2082136 N chr5 2082200 N DEL 10
SRR1766474.531252 chr5 2082209 N chr5 2082964 N DUP 13
SRR1766464.791940 chr5 2082226 N chr5 2082981 N DUP 2
SRR1766469.5618666 chr5 2082231 N chr5 2082293 N DUP 5
SRR1766479.3504639 chr5 2082290 N chr5 2082352 N DUP 5
SRR1766474.7242484 chr5 2082290 N chr5 2082352 N DUP 5
SRR1766457.7272215 chr5 2082321 N chr5 2082700 N DEL 5
SRR1766478.6279524 chr5 2082321 N chr5 2082700 N DEL 5
SRR1766485.8949923 chr5 2082447 N chr5 2082700 N DEL 15
SRR1766452.7887974 chr5 2082673 N chr5 2082924 N DUP 2
SRR1766484.4042638 chr5 2082321 N chr5 2082700 N DEL 5
SRR1766450.954317 chr5 2082321 N chr5 2082700 N DEL 5
SRR1766469.1366315 chr5 2082258 N chr5 2082700 N DEL 5
SRR1766484.8580938 chr5 2082135 N chr5 2082703 N DEL 5
SRR1766450.5255427 chr5 2082196 N chr5 2082384 N DUP 11
SRR1766485.4625684 chr5 2082136 N chr5 2082704 N DEL 5
SRR1766469.1366315 chr5 2082136 N chr5 2082704 N DEL 5
SRR1766480.3532710 chr5 2082137 N chr5 2082705 N DEL 5
SRR1766442.36890550 chr5 2082291 N chr5 2082733 N DEL 10
SRR1766461.9669304 chr5 2082731 N chr5 2082793 N DUP 10
SRR1766461.2408665 chr5 2082353 N chr5 2082793 N DUP 5
SRR1766451.8830020 chr5 2082249 N chr5 2082878 N DUP 8
SRR1766465.4384166 chr5 2082226 N chr5 2082353 N DEL 10
SRR1766467.11307747 chr5 2082316 N chr5 2082821 N DEL 10
SRR1766470.6948601 chr5 2082262 N chr5 2082830 N DEL 5
SRR1766455.148065 chr5 2082190 N chr5 2082821 N DEL 15
SRR1766442.25830866 chr5 2082316 N chr5 2082821 N DEL 18
SRR1766453.4739312 chr5 2082378 N chr5 2082820 N DEL 5
SRR1766456.182501 chr5 2082378 N chr5 2082820 N DEL 5
SRR1766468.1486245 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766457.7798515 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766442.35123216 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766456.2077572 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766466.7925634 chr5 2082378 N chr5 2082820 N DEL 5
SRR1766478.10028038 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766481.6592463 chr5 2082380 N chr5 2082822 N DEL 15
SRR1766453.9884496 chr5 2082196 N chr5 2082888 N DUP 10
SRR1766471.5912184 chr5 2082135 N chr5 2082829 N DEL 8
SRR1766461.5710385 chr5 2082338 N chr5 2082906 N DEL 15
SRR1766461.4353759 chr5 2082198 N chr5 2082953 N DUP 5
SRR1766466.5686427 chr5 2082341 N chr5 2082909 N DEL 5
SRR1766450.2008726 chr5 2082464 N chr5 2082906 N DEL 5
SRR1766479.12825593 chr5 2082906 N chr5 2082968 N DUP 5
SRR1766486.2088918 chr5 2082317 N chr5 2082885 N DEL 10
SRR1766459.10980685 chr5 2082906 N chr5 2082968 N DUP 9
SRR1766446.2988791 chr5 2082906 N chr5 2082968 N DUP 10
SRR1766458.9252244 chr5 2082906 N chr5 2082968 N DUP 18
SRR1766473.7429139 chr5 2082172 N chr5 2082866 N DEL 3
SRR1766471.8172915 chr5 2082474 N chr5 2082916 N DEL 10
SRR1766485.7238556 chr5 2082906 N chr5 2082968 N DUP 21
SRR1766481.5992998 chr17 81432869 N chr17 81432992 N DEL 8
SRR1766468.6448089 chr7 132647055 N chr7 132647160 N DEL 5
SRR1766444.4837942 chr7 132647014 N chr7 132647345 N DEL 55
SRR1766447.4250475 chr7 132646995 N chr7 132647208 N DUP 10
SRR1766467.7397862 chr7 132647328 N chr7 132647445 N DEL 1
SRR1766450.5524231 chr7 132647045 N chr7 132647490 N DEL 5
SRR1766455.6214342 chr7 132647157 N chr7 132647498 N DEL 5
SRR1766458.847579 chr12 82639286 N chr12 82639412 N DUP 5
SRR1766455.560933 chr12 82639292 N chr12 82639600 N DUP 5
SRR1766471.10617810 chr12 82639304 N chr12 82639361 N DUP 5
SRR1766471.10331568 chr12 82639354 N chr12 82639935 N DUP 5
SRR1766453.7361038 chr12 82639653 N chr12 82639736 N DUP 5
SRR1766442.37684280 chr12 82640372 N chr12 82640563 N DEL 14
SRR1766461.10673178 chr12 82639946 N chr12 82640282 N DEL 16
SRR1766457.3600 chr12 82639946 N chr12 82640282 N DEL 15
SRR1766454.7802014 chr12 82640266 N chr12 82640401 N DUP 13
SRR1766442.10124210 chr12 82640203 N chr12 82640312 N DEL 5
SRR1766452.142368 chr12 82639421 N chr12 82640417 N DEL 1
SRR1766464.7757806 chr12 82639694 N chr12 82640413 N DEL 5
SRR1766462.8806091 chr4 38880239 N chr4 38880295 N DEL 18
SRR1766459.10336075 chr4 38880239 N chr4 38880295 N DEL 20
SRR1766463.5569745 chr4 189413752 N chr4 189413842 N DEL 5
SRR1766449.10020969 chr4 189413874 N chr4 189414053 N DEL 5
SRR1766466.1781678 chr4 189413789 N chr4 189413968 N DEL 5
SRR1766474.9514344 chr4 189413802 N chr4 189413981 N DEL 2
SRR1766445.5113819 chr4 189413820 N chr4 189413999 N DEL 5
SRR1766480.6249173 chr4 189413856 N chr4 189414035 N DEL 6
SRR1766469.6736847 chr4 189413856 N chr4 189414035 N DEL 5
SRR1766464.6001581 chr16 83617573 N chr16 83617628 N DUP 2
SRR1766473.4127737 chr16 83617573 N chr16 83617628 N DUP 2
SRR1766463.4207033 chr16 83617573 N chr16 83617628 N DUP 5
SRR1766455.730428 chr16 83617573 N chr16 83617628 N DUP 5
SRR1766470.3446292 chr16 83617587 N chr16 83617644 N DEL 5
SRR1766461.9637774 chr16 83617588 N chr16 83617645 N DEL 5
SRR1766442.7108494 chr16 83617591 N chr16 83617648 N DEL 5
SRR1766475.10911978 chr16 83617600 N chr16 83617657 N DEL 1
SRR1766478.9929418 chr16 83617600 N chr16 83617657 N DEL 1
SRR1766462.4400180 chr14 104527464 N chr14 104527754 N DEL 5
SRR1766480.1944846 chr14 104527334 N chr14 104527479 N DUP 2
SRR1766446.1317252 chr14 104527361 N chr14 104527416 N DEL 2
SRR1766467.11216392 chr14 104527474 N chr14 104527593 N DUP 5
SRR1766483.10278979 chr14 104527482 N chr14 104527770 N DUP 1
SRR1766462.1575328 chr14 104527491 N chr14 104527914 N DUP 9
SRR1766449.3849837 chr14 104527334 N chr14 104527768 N DUP 1
SRR1766468.2074319 chr2 206104325 N chr2 206104473 N DEL 44
SRR1766453.10124286 chr7 56268615 N chr7 56268680 N DEL 1
SRR1766456.5791334 chr1 169273385 N chr1 169273788 N DEL 14
SRR1766455.6740250 chr1 169273544 N chr1 169273947 N DEL 5
SRR1766454.7421730 chr1 169273377 N chr1 169273780 N DEL 10
SRR1766464.9403336 chr1 169273389 N chr1 169273792 N DEL 9
SRR1766466.8733007 chr5 144847782 N chr5 144848047 N DEL 10
SRR1766486.9950591 chr7 40377351 N chr7 40377404 N DEL 46
SRR1766478.7707663 chr7 40377351 N chr7 40377404 N DEL 46
SRR1766458.9347111 chr7 40377326 N chr7 40377404 N DEL 42
SRR1766467.4403153 chr12 110867120 N chr12 110867348 N DEL 1
SRR1766479.11080116 chr12 110867472 N chr12 110867649 N DEL 10
SRR1766478.498748 chr12 110867070 N chr12 110867472 N DUP 5
SRR1766474.7752301 chr12 110867025 N chr12 110867603 N DUP 4
SRR1766477.10916460 chr12 110867070 N chr12 110867648 N DUP 1
SRR1766446.6387964 chr12 110867070 N chr12 110867472 N DUP 5
SRR1766476.6082857 chr12 110867073 N chr12 110867653 N DEL 5
SRR1766454.3643285 chr12 110867070 N chr12 110867472 N DUP 5
SRR1766477.3735648 chr12 110867070 N chr12 110867472 N DUP 5
SRR1766481.3652032 chr12 110867099 N chr12 110867677 N DUP 5
SRR1766453.9246010 chr12 110867070 N chr12 110867472 N DUP 5
SRR1766468.578644 chr12 110867194 N chr12 110867459 N DEL 5
SRR1766442.25827805 chr12 110867120 N chr12 110867747 N DUP 11
SRR1766475.8541565 chr12 110867098 N chr12 110867676 N DUP 1
SRR1766452.4317184 chr12 110867029 N chr12 110867204 N DUP 2
SRR1766453.3528027 chr12 110867101 N chr12 110867278 N DUP 5
SRR1766452.3582707 chr12 110867038 N chr12 110867215 N DEL 5
SRR1766468.5788729 chr12 110867074 N chr12 110867300 N DUP 5
SRR1766478.5240337 chr12 110867148 N chr12 110867374 N DUP 5
SRR1766482.10856527 chr12 110867148 N chr12 110867374 N DUP 5
SRR1766444.418453 chr12 110867205 N chr12 110867431 N DUP 5
SRR1766462.7066876 chr12 110867205 N chr12 110867431 N DUP 5
SRR1766473.10508484 chr12 110867116 N chr12 110867469 N DUP 5
SRR1766458.7799853 chr12 110867395 N chr12 110867748 N DEL 5
SRR1766442.25204273 chr12 110867395 N chr12 110867748 N DEL 5
SRR1766480.4873267 chr12 110867009 N chr12 110867086 N DUP 5
SRR1766466.2645213 chr12 110867266 N chr12 110867494 N DEL 5
SRR1766486.5346696 chr12 110867266 N chr12 110867494 N DEL 5
SRR1766482.11152785 chr12 110867494 N chr12 110867845 N DUP 5
SRR1766462.7066876 chr12 110867266 N chr12 110867494 N DEL 5
SRR1766486.5346696 chr12 110867266 N chr12 110867494 N DEL 10
SRR1766449.8393221 chr12 110867266 N chr12 110867494 N DEL 5
SRR1766480.6170934 chr12 110867266 N chr12 110867494 N DEL 10
SRR1766442.10523014 chr12 110867266 N chr12 110867494 N DEL 5
SRR1766459.9475523 chr12 110867135 N chr12 110867539 N DEL 5
SRR1766446.4737884 chr12 110867510 N chr12 110867861 N DUP 4
SRR1766448.3276346 chr12 110867285 N chr12 110867512 N DEL 7
SRR1766475.6125733 chr12 110867109 N chr12 110867562 N DEL 10
SRR1766473.4120718 chr12 110867109 N chr12 110867562 N DEL 5
SRR1766450.4354291 chr12 110867014 N chr12 110867592 N DUP 5
SRR1766467.3543220 chr12 110867113 N chr12 110867566 N DEL 5
SRR1766453.693926 chr12 110867014 N chr12 110867592 N DUP 5
SRR1766473.5176837 chr12 110867278 N chr12 110867678 N DUP 5
SRR1766444.4674284 chr12 110867350 N chr12 110867652 N DUP 5
SRR1766482.5260876 chr12 110867014 N chr12 110867592 N DUP 5
SRR1766470.7426955 chr12 110867014 N chr12 110867592 N DUP 5
SRR1766460.164932 chr12 110867014 N chr12 110867592 N DUP 5
SRR1766466.9048096 chr12 110867019 N chr12 110867597 N DUP 5
SRR1766448.6070695 chr12 110867036 N chr12 110867616 N DEL 5
SRR1766464.4061348 chr12 110867472 N chr12 110867649 N DEL 5
SRR1766454.9696847 chr12 110867075 N chr12 110867653 N DUP 4
SRR1766442.15290632 chr12 110867073 N chr12 110867653 N DEL 5
SRR1766464.3133171 chr12 110867073 N chr12 110867653 N DEL 5
SRR1766460.164932 chr12 110867073 N chr12 110867653 N DEL 5
SRR1766471.9667961 chr12 110867073 N chr12 110867653 N DEL 5
SRR1766451.6830640 chr12 110867078 N chr12 110867658 N DEL 5
SRR1766450.1529907 chr12 110867144 N chr12 110867723 N DEL 7
SRR1766454.9696847 chr12 110867155 N chr12 110867383 N DEL 5
SRR1766471.3801521 chr12 110867119 N chr12 110867748 N DEL 5
SRR1766444.5139845 chr9 125623367 N chr9 125623678 N DUP 5
SRR1766477.431558 chr9 125623549 N chr9 125623664 N DUP 1
SRR1766471.7077942 chr9 125623558 N chr9 125623633 N DUP 3
SRR1766465.8775750 chr9 125623453 N chr9 125623805 N DUP 2
SRR1766451.8692874 chr9 125623854 N chr9 125623951 N DUP 5
SRR1766486.7937904 chr3 198076499 N chr3 198076566 N DEL 15
SRR1766463.1352146 chr1 227741089 N chr1 227741284 N DUP 5
SRR1766451.5195573 chr3 181926025 N chr3 181926339 N DUP 1
SRR1766442.603612 chr22 41316229 N chr22 41316911 N DEL 5
SRR1766463.2959732 chr22 41316254 N chr22 41316555 N DUP 5
SRR1766468.5656870 chr22 41316443 N chr22 41316746 N DEL 5
SRR1766486.695665 chr4 36484994 N chr4 36485105 N DEL 19
SRR1766469.7818746 chr4 36484995 N chr4 36485106 N DEL 14
SRR1766474.716550 chr4 36485001 N chr4 36485112 N DEL 8
SRR1766475.3842078 chr4 36485002 N chr4 36485113 N DEL 7
SRR1766471.6738478 chr4 36485005 N chr4 36485116 N DEL 4
SRR1766462.9877296 chr2 86833656 N chr2 86833717 N DEL 5
SRR1766446.8250341 chr9 118675594 N chr9 118675735 N DUP 5
SRR1766456.1621067 chr17 77829034 N chr17 77829244 N DUP 5
SRR1766457.989236 chr17 77828939 N chr17 77829039 N DEL 5
SRR1766485.12098834 chr17 77829019 N chr17 77829172 N DUP 5
SRR1766463.5807244 chr17 77828945 N chr17 77829273 N DUP 5
SRR1766460.6147325 chr2 164818738 N chr2 164818797 N DEL 6
SRR1766454.8862485 chr2 164818738 N chr2 164818797 N DEL 9
SRR1766443.2206782 chr2 164818738 N chr2 164818797 N DEL 10
SRR1766463.6435315 chr13 103600738 N chr13 103600889 N DEL 5
SRR1766457.5854277 chr13 103600738 N chr13 103600889 N DEL 5
SRR1766445.8277886 chr13 103600675 N chr13 103600754 N DEL 5
SRR1766466.10313350 chr13 103600758 N chr13 103600907 N DUP 5
SRR1766442.40114078 chr13 103600760 N chr13 103600909 N DUP 5
SRR1766455.6766269 chr13 103600761 N chr13 103600910 N DUP 4
SRR1766450.8427630 chr13 103600761 N chr13 103600910 N DUP 4
SRR1766486.4613960 chr2 87092042 N chr2 87092141 N DUP 5
SRR1766463.5271076 chr2 87092042 N chr2 87092141 N DUP 5
SRR1766451.4231903 chr2 87092057 N chr2 87092158 N DEL 5
SRR1766472.10090472 chr12 130055053 N chr12 130055191 N DUP 6
SRR1766467.3610157 chr12 130055314 N chr12 130055455 N DEL 10
SRR1766455.5570942 chr12 130055276 N chr12 130055438 N DEL 10
SRR1766467.739141 chr12 130055532 N chr12 130055663 N DUP 13
SRR1766467.5596904 chr12 130055704 N chr12 130055772 N DEL 5
SRR1766445.10450722 chr16 22939832 N chr16 22939986 N DEL 5
SRR1766459.4947587 chr16 22939832 N chr16 22939986 N DEL 15
SRR1766458.6881922 chr16 22939832 N chr16 22939986 N DEL 5
SRR1766471.9068161 chr16 22939832 N chr16 22939986 N DEL 15
SRR1766474.342384 chr16 22939832 N chr16 22939986 N DEL 5
SRR1766464.6009955 chr16 22939878 N chr16 22940083 N DEL 5
SRR1766442.20254737 chr16 22939878 N chr16 22940083 N DEL 5
SRR1766445.3124665 chr16 22939889 N chr16 22940247 N DEL 1
SRR1766465.11114509 chr16 22939906 N chr16 22939958 N DEL 2
SRR1766480.5689529 chr16 22939878 N chr16 22940083 N DEL 5
SRR1766476.11080999 chr16 22939878 N chr16 22940083 N DEL 9
SRR1766485.4627710 chr16 22939878 N chr16 22940083 N DEL 14
SRR1766467.1384458 chr16 22939939 N chr16 22940042 N DEL 10
SRR1766449.5204186 chr16 22939935 N chr16 22940395 N DEL 25
SRR1766473.8981300 chr16 22939921 N chr16 22940075 N DEL 5
SRR1766446.8457225 chr16 22940023 N chr16 22940075 N DEL 3
SRR1766442.24138589 chr16 22939938 N chr16 22940039 N DUP 5
SRR1766484.4375114 chr16 22940023 N chr16 22940075 N DEL 5
SRR1766482.8020261 chr16 22940023 N chr16 22940075 N DEL 5
SRR1766449.2813098 chr16 22940037 N chr16 22940395 N DEL 5
SRR1766457.6908869 chr16 22939832 N chr16 22939986 N DEL 10
SRR1766466.8348564 chr16 22939832 N chr16 22939986 N DEL 10
SRR1766453.3983640 chr16 22940083 N chr16 22940339 N DEL 5
SRR1766470.5536249 chr16 22940075 N chr16 22940125 N DUP 5
SRR1766476.3892989 chr16 22939992 N chr16 22940093 N DUP 5
SRR1766445.7186460 chr16 22939972 N chr16 22940075 N DEL 5
SRR1766474.8870799 chr16 22939992 N chr16 22940144 N DUP 1
SRR1766459.4947587 chr16 22939931 N chr16 22940085 N DEL 5
SRR1766443.1096478 chr16 22940075 N chr16 22940176 N DUP 10
SRR1766464.5020783 chr16 22939824 N chr16 22940131 N DEL 1
SRR1766476.11080999 chr16 22940039 N chr16 22940193 N DEL 5
SRR1766442.13450978 chr16 22940292 N chr16 22940395 N DEL 5
SRR1766468.3553453 chr16 22939903 N chr16 22940210 N DEL 5
SRR1766471.9068161 chr16 22939856 N chr16 22940214 N DEL 5
SRR1766459.1470423 chr16 22939824 N chr16 22940233 N DEL 1
SRR1766451.4714494 chr16 22940033 N chr16 22940289 N DEL 5
SRR1766442.17547546 chr16 22940084 N chr16 22940338 N DUP 5
SRR1766473.6722629 chr16 22940084 N chr16 22940338 N DUP 5
SRR1766442.5186914 chr16 22939931 N chr16 22940289 N DEL 5
SRR1766465.11114509 chr16 22940084 N chr16 22940338 N DUP 5
SRR1766458.6881922 chr16 22939933 N chr16 22940291 N DEL 5
SRR1766445.3124665 chr16 22939981 N chr16 22940339 N DEL 10
SRR1766442.20254737 chr16 22939972 N chr16 22940330 N DEL 5
SRR1766450.10621546 chr16 22940054 N chr16 22940361 N DEL 5
SRR1766449.5204186 chr16 22939863 N chr16 22940374 N DEL 2
SRR1766483.2116312 chr16 22940176 N chr16 22940432 N DEL 5
SRR1766486.8558441 chr16 22940059 N chr16 22940417 N DEL 10
SRR1766443.7356166 chr16 22939859 N chr16 22940472 N DEL 10
SRR1766471.299641 chr16 22939837 N chr16 22940450 N DEL 3
SRR1766451.9705334 chr2 203066848 N chr2 203067192 N DEL 1
SRR1766444.4080153 chr2 203066954 N chr2 203067184 N DEL 7
SRR1766480.3534626 chr2 203066889 N chr2 203067157 N DUP 5
SRR1766447.6177243 chr2 203067006 N chr2 203067157 N DEL 2
SRR1766470.4958127 chr2 203067117 N chr2 203067192 N DEL 1
SRR1766475.7297021 chr2 203067146 N chr2 203067218 N DEL 12
SRR1766453.10854310 chr2 203067006 N chr2 203067226 N DUP 5
SRR1766460.2929372 chr2 203067006 N chr2 203067226 N DUP 5
SRR1766442.8466988 chr2 203067024 N chr2 203067246 N DEL 1
SRR1766480.1189412 chr14 85847829 N chr14 85848674 N DEL 5
SRR1766485.43942 chr14 85847716 N chr14 85847797 N DEL 17
SRR1766452.5001147 chr14 85847716 N chr14 85847797 N DEL 17
SRR1766452.6262241 chr14 85847716 N chr14 85847797 N DEL 17
SRR1766460.2025712 chr14 85847842 N chr14 85848173 N DEL 26
SRR1766467.11107955 chr14 85847842 N chr14 85848173 N DEL 26
SRR1766482.7098379 chr14 85847842 N chr14 85848173 N DEL 20
SRR1766448.8686377 chr14 85847842 N chr14 85848173 N DEL 14
SRR1766464.3307051 chr14 85847831 N chr14 85848304 N DUP 5
SRR1766479.5509182 chr14 85847831 N chr14 85848304 N DUP 5
SRR1766484.6081919 chr14 85847718 N chr14 85847841 N DEL 9
SRR1766447.7863724 chr14 85847718 N chr14 85847841 N DEL 9
SRR1766474.1578178 chr14 85847718 N chr14 85847841 N DEL 9
SRR1766457.2890363 chr14 85847718 N chr14 85847841 N DEL 9
SRR1766442.6395756 chr14 85847980 N chr14 85848143 N DEL 7
SRR1766442.18764324 chr14 85847980 N chr14 85848143 N DEL 7
SRR1766471.213505 chr14 85847853 N chr14 85848012 N DUP 9
SRR1766479.9491425 chr14 85848012 N chr14 85848143 N DEL 1
SRR1766467.3561983 chr14 85847853 N chr14 85848012 N DUP 9
SRR1766471.10228021 chr14 85847853 N chr14 85848012 N DUP 9
SRR1766485.1450157 chr14 85848012 N chr14 85848143 N DEL 2
SRR1766448.11086691 chr14 85847980 N chr14 85848143 N DEL 4
SRR1766480.1189412 chr14 85847980 N chr14 85848143 N DEL 6
SRR1766447.548212 chr14 85847853 N chr14 85847980 N DUP 9
SRR1766479.3017748 chr14 85847853 N chr14 85847980 N DUP 9
SRR1766447.1682721 chr14 85847853 N chr14 85847980 N DUP 9
SRR1766479.5317535 chr14 85847853 N chr14 85847980 N DUP 9
SRR1766457.4905689 chr14 85847853 N chr14 85847980 N DUP 9
SRR1766485.8613481 chr14 85847853 N chr14 85847980 N DUP 9
SRR1766459.5049270 chr14 85847980 N chr14 85848205 N DEL 9
SRR1766475.513567 chr14 85847980 N chr14 85848239 N DEL 11
SRR1766484.10538475 chr14 85847853 N chr14 85848202 N DUP 7
SRR1766468.5553988 chr14 85847980 N chr14 85848239 N DEL 13
SRR1766477.3232805 chr14 85847948 N chr14 85848239 N DEL 20
SRR1766480.6845697 chr14 85847853 N chr14 85848202 N DUP 7
SRR1766450.201548 chr14 85847853 N chr14 85848202 N DUP 7
SRR1766449.7372603 chr14 85847853 N chr14 85848202 N DUP 7
SRR1766473.7152043 chr14 85847850 N chr14 85848205 N DEL 7
SRR1766472.5219863 chr14 85847850 N chr14 85848205 N DEL 7
SRR1766485.1450157 chr14 85847850 N chr14 85848205 N DEL 7
SRR1766456.615286 chr14 85847948 N chr14 85848239 N DEL 14
SRR1766477.7886641 chr14 85847850 N chr14 85848205 N DEL 7
SRR1766454.6404747 chr14 85847852 N chr14 85848207 N DEL 7
SRR1766460.9172 chr14 85847948 N chr14 85848239 N DEL 14
SRR1766486.4783513 chr14 85847948 N chr14 85848239 N DEL 14
SRR1766479.4721047 chr14 85847855 N chr14 85848210 N DEL 7
SRR1766474.5834590 chr14 85847857 N chr14 85848212 N DEL 7
SRR1766479.8146751 chr14 85847916 N chr14 85848239 N DEL 14
SRR1766459.10919837 chr14 85847850 N chr14 85848239 N DEL 14
SRR1766461.4501618 chr14 85847850 N chr14 85848239 N DEL 14
SRR1766442.5325705 chr14 85848358 N chr14 85848425 N DEL 4
SRR1766466.974042 chr14 85848185 N chr14 85848252 N DEL 2
SRR1766476.7988844 chr14 85848184 N chr14 85848251 N DEL 3
SRR1766476.6646398 chr14 85848411 N chr14 85848480 N DUP 3
SRR1766442.41278438 chr14 85847888 N chr14 85848393 N DEL 5
SRR1766442.10830330 chr14 85847858 N chr14 85848397 N DEL 9
SRR1766474.1540014 chr14 85847831 N chr14 85848674 N DUP 1
SRR1766475.8544493 chr14 85847831 N chr14 85848674 N DUP 5
SRR1766456.4477421 chr14 85847853 N chr14 85848698 N DEL 5
SRR1766450.8090954 chr14 85847853 N chr14 85848698 N DEL 5
SRR1766482.2091417 chr1 39093455 N chr1 39093631 N DUP 1
SRR1766451.2657643 chr13 113980377 N chr13 113980504 N DEL 9
SRR1766460.11113442 chr13 113980361 N chr13 113980486 N DEL 2
SRR1766445.6889230 chr16 88798349 N chr16 88798495 N DUP 10
SRR1766447.4960551 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766451.1294356 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766480.6458147 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766448.7728452 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766476.10535936 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766471.3981639 chr3 84516444 N chr3 84516521 N DUP 3
SRR1766483.6685656 chr2 194048799 N chr2 194048858 N DUP 5
SRR1766469.10217048 chr2 194048797 N chr2 194048856 N DUP 5
SRR1766485.4770490 chr7 56758204 N chr7 56758256 N DUP 9
SRR1766446.5048959 chr7 56758269 N chr7 56758328 N DUP 10
SRR1766456.5651620 chr7 56758157 N chr7 56758232 N DEL 7
SRR1766442.28069048 chr7 56758189 N chr7 56758299 N DEL 6
SRR1766452.5143620 chr7 56758159 N chr7 56758299 N DEL 5
SRR1766474.5652012 chr7 56758246 N chr7 56758300 N DEL 5
SRR1766446.1673506 chr7 56758249 N chr7 56758303 N DEL 5
SRR1766473.5150155 chr9 10323351 N chr9 10323437 N DEL 8
SRR1766473.8006928 chrX 41507258 N chrX 41507388 N DUP 19
SRR1766446.9253113 chrX 41507250 N chrX 41507504 N DUP 4
SRR1766449.9886848 chr18 41577544 N chr18 41577603 N DEL 7
SRR1766471.11093861 chr18 41577544 N chr18 41577603 N DEL 7
SRR1766444.673217 chr18 41577546 N chr18 41577601 N DUP 7
SRR1766464.51547 chr18 41577546 N chr18 41577601 N DUP 7
SRR1766462.8335824 chr18 41577546 N chr18 41577601 N DUP 7
SRR1766477.8194992 chr18 41577546 N chr18 41577601 N DUP 7
SRR1766442.26236837 chr18 41577546 N chr18 41577601 N DUP 7
SRR1766482.6273841 chr18 41577546 N chr18 41577601 N DUP 7
SRR1766461.9587488 chr18 41577546 N chr18 41577601 N DUP 7
SRR1766459.3109839 chr18 41577578 N chr18 41577669 N DUP 17
SRR1766480.2690849 chr18 41577484 N chr18 41577551 N DEL 9
SRR1766468.7427780 chr18 41577485 N chr18 41577552 N DEL 8
SRR1766479.11271671 chr18 41577483 N chr18 41577564 N DEL 7
SRR1766484.4335905 chr18 41577533 N chr18 41577604 N DEL 3
SRR1766467.1751958 chr18 41577521 N chr18 41577616 N DEL 7
SRR1766473.7966644 chr18 41577521 N chr18 41577616 N DEL 7
SRR1766463.1418286 chr16 33174144 N chr16 33174199 N DUP 1
SRR1766479.567655 chr1 191089530 N chr1 191089689 N DEL 5
SRR1766446.8869254 chr1 191089479 N chr1 191089531 N DUP 5
SRR1766446.8869254 chr1 191089479 N chr1 191089531 N DUP 6
SRR1766447.9364277 chr1 191089479 N chr1 191089531 N DUP 9
SRR1766448.356980 chr1 191089495 N chr1 191089549 N DEL 10
SRR1766476.6334867 chr1 191089497 N chr1 191089551 N DEL 8
SRR1766442.20149232 chr1 191089419 N chr1 191089665 N DUP 5
SRR1766466.3560216 chr8 142991125 N chr8 142991313 N DUP 6
SRR1766442.27113742 chr8 142991218 N chr8 142991274 N DEL 5
SRR1766465.9799946 chr8 142991129 N chr8 142991326 N DEL 13
SRR1766449.3814756 chr17 83172608 N chr17 83173590 N DEL 6
SRR1766475.2455562 chr17 83172590 N chr17 83172665 N DUP 5
SRR1766476.3608551 chr17 83172588 N chr17 83172663 N DUP 5
SRR1766459.10714832 chr17 83172596 N chr17 83173121 N DUP 5
SRR1766442.15018479 chr17 83172628 N chr17 83172965 N DUP 5
SRR1766451.1754076 chr17 83172625 N chr17 83172776 N DEL 10
SRR1766452.4099532 chr17 83172538 N chr17 83172725 N DUP 15
SRR1766445.132210 chr17 83172598 N chr17 83172749 N DEL 10
SRR1766486.3638211 chr17 83172560 N chr17 83172749 N DEL 13
SRR1766450.6781346 chr17 83172625 N chr17 83172814 N DEL 7
SRR1766443.5260056 chr17 83172788 N chr17 83172863 N DUP 10
SRR1766481.8658521 chr17 83172625 N chr17 83172776 N DEL 10
SRR1766482.8305591 chr17 83172784 N chr17 83173538 N DUP 11
SRR1766474.8876135 chr17 83173214 N chr17 83173669 N DEL 19
SRR1766485.329596 chr17 83172521 N chr17 83172860 N DUP 14
SRR1766470.10254926 chr17 83172693 N chr17 83173447 N DEL 1
SRR1766457.459335 chr17 83173069 N chr17 83173295 N DUP 5
SRR1766472.9689428 chr17 83172619 N chr17 83172694 N DUP 19
SRR1766453.8373625 chr17 83173101 N chr17 83173555 N DUP 9
SRR1766442.30436134 chr17 83172580 N chr17 83173069 N DEL 16
SRR1766448.9952925 chr17 83172689 N chr17 83173481 N DEL 28
SRR1766463.7038479 chr17 83172689 N chr17 83173367 N DEL 20
SRR1766458.5118080 chr17 83172651 N chr17 83173367 N DEL 5
SRR1766467.7585776 chr17 83172708 N chr17 83173690 N DEL 8
SRR1766451.251250 chr17 83172715 N chr17 83173697 N DEL 6
SRR1766460.9694844 chr17 83173540 N chr17 83173691 N DEL 9
SRR1766450.1975808 chr8 14847784 N chr8 14847891 N DUP 5
SRR1766442.8424595 chr10 46136053 N chr10 46136184 N DEL 5
SRR1766485.10379071 chr10 46136090 N chr10 46136189 N DEL 1
SRR1766463.8855270 chr10 46136056 N chr10 46136105 N DUP 10
SRR1766452.2129119 chr10 46136056 N chr10 46136105 N DUP 12
SRR1766455.4201587 chr10 46136103 N chr10 46136168 N DEL 15
SRR1766455.1355315 chr10 46136090 N chr10 46136153 N DEL 11
SRR1766463.5064477 chr10 46136090 N chr10 46136153 N DEL 13
SRR1766470.1464109 chr10 46136090 N chr10 46136153 N DEL 13
SRR1766446.2336436 chr10 46136103 N chr10 46136168 N DEL 21
SRR1766444.3439636 chr10 46136092 N chr10 46136155 N DUP 9
SRR1766486.3944116 chr10 46136069 N chr10 46136200 N DUP 7
SRR1766451.2805452 chr10 46136131 N chr10 46136200 N DUP 11
SRR1766465.9136980 chr10 46136136 N chr10 46136205 N DUP 16
SRR1766472.7832035 chr10 46136116 N chr10 46136177 N DEL 3
SRR1766462.1010556 chr10 46136116 N chr10 46136177 N DEL 3
SRR1766469.10406037 chr8 144620132 N chr8 144620334 N DEL 5
SRR1766470.6016246 chr8 144620276 N chr8 144620353 N DUP 5
SRR1766474.10273409 chr13 18943421 N chr13 18944062 N DEL 5
SRR1766474.8206167 chr13 18943575 N chr13 18944435 N DEL 5
SRR1766472.192973 chr13 18943999 N chr13 18944435 N DEL 4
SRR1766483.6151220 chr13 18943482 N chr13 18943907 N DEL 5
SRR1766458.6546707 chr13 18943522 N chr13 18943947 N DEL 1
SRR1766455.6065868 chr13 18943468 N chr13 18944110 N DEL 2
SRR1766467.8816434 chr13 18944057 N chr13 18944691 N DUP 3
SRR1766480.3435731 chr13 18944234 N chr13 18944452 N DEL 1
SRR1766468.4257555 chr13 18944234 N chr13 18944452 N DEL 2
SRR1766447.4947984 chr13 18944260 N chr13 18944476 N DUP 5
SRR1766442.4284622 chr13 18944429 N chr13 18945058 N DUP 5
SRR1766471.10465404 chr13 18944211 N chr13 18944429 N DEL 10
SRR1766472.6005983 chr13 18943782 N chr13 18944431 N DEL 5
SRR1766465.8064377 chr13 18944529 N chr13 18945170 N DEL 20
SRR1766446.2587259 chr13 18943452 N chr13 18944939 N DUP 5
SRR1766445.8252043 chr19 16215328 N chr19 16215501 N DEL 6
SRR1766478.11923371 chr19 16215328 N chr19 16215501 N DEL 8
SRR1766446.8225216 chrX 46395879 N chrX 46396105 N DEL 5
SRR1766448.274281 chrX 46395879 N chrX 46396105 N DEL 5
SRR1766479.11267620 chrX 46395879 N chrX 46396105 N DEL 9
SRR1766442.12326902 chrX 46395797 N chrX 46395974 N DEL 4
SRR1766446.8225216 chrX 46395846 N chrX 46396072 N DEL 5
SRR1766457.2094111 chrX 46395780 N chrX 46396177 N DUP 1
SRR1766473.1106268 chrX 46396009 N chrX 46396181 N DUP 2
SRR1766465.1776203 chrX 46395854 N chrX 46396251 N DUP 5
SRR1766467.6239920 chrX 46395854 N chrX 46396251 N DUP 5
SRR1766485.9812571 chrX 46396353 N chrX 46396474 N DEL 2
SRR1766451.567230 chrX 46395877 N chrX 46396276 N DEL 1
SRR1766448.274281 chrX 46396346 N chrX 46396465 N DUP 5
SRR1766452.10157088 chrX 46396389 N chrX 46396508 N DUP 5
SRR1766484.10734055 chrX 46396389 N chrX 46396508 N DUP 5
SRR1766470.9742582 chr2 129735706 N chr2 129735776 N DEL 5
SRR1766459.8489642 chr2 129735711 N chr2 129735781 N DEL 5
SRR1766478.3136656 chr2 129735714 N chr2 129735784 N DEL 5
SRR1766485.5811589 chr2 129735720 N chr2 129735994 N DUP 13
SRR1766479.5661079 chr2 129735983 N chr2 129736036 N DUP 3
SRR1766482.1963407 chr5 175050953 N chr5 175051008 N DUP 25
SRR1766449.1821551 chr5 175050953 N chr5 175051008 N DUP 36
SRR1766482.12957866 chr5 175050969 N chr5 175051024 N DUP 27
SRR1766455.3355411 chr5 175050969 N chr5 175051024 N DUP 27
SRR1766442.39217338 chr5 175050953 N chr5 175051008 N DUP 37
SRR1766461.5058047 chr5 175050953 N chr5 175051008 N DUP 37
SRR1766475.3288234 chr5 175050955 N chr5 175051037 N DUP 26
SRR1766454.8584461 chr5 175050955 N chr5 175051037 N DUP 28
SRR1766467.11469131 chr5 175050955 N chr5 175051037 N DUP 24
SRR1766459.7085575 chr5 175050955 N chr5 175051037 N DUP 30
SRR1766458.4133442 chr5 175050945 N chr5 175051029 N DUP 34
SRR1766442.35734643 chr5 175050945 N chr5 175051029 N DUP 46
SRR1766445.504216 chr5 175050945 N chr5 175051029 N DUP 45
SRR1766447.4007054 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766447.9114426 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766448.4957899 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766448.7792711 chr5 175050955 N chr5 175051037 N DUP 39
SRR1766452.10321710 chr5 175050945 N chr5 175051029 N DUP 38
SRR1766455.553817 chr5 175050953 N chr5 175051008 N DUP 42
SRR1766455.6790559 chr5 175050953 N chr5 175051008 N DUP 31
SRR1766463.148498 chr5 175050945 N chr5 175051029 N DUP 43
SRR1766471.6238285 chr5 175050945 N chr5 175051029 N DUP 40
SRR1766472.4827124 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766479.9037325 chr5 175050945 N chr5 175051029 N DUP 38
SRR1766481.11873666 chr5 175050945 N chr5 175051029 N DUP 36
SRR1766483.8909131 chr5 175050944 N chr5 175051028 N DUP 41
SRR1766447.4007054 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766451.1959023 chr5 175050945 N chr5 175051029 N DUP 38
SRR1766454.6574963 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766456.4092508 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766457.8785463 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766463.602383 chr5 175050945 N chr5 175051029 N DUP 41
SRR1766466.2065916 chr5 175050945 N chr5 175051029 N DUP 45
SRR1766469.4497478 chr5 175050945 N chr5 175051029 N DUP 46
SRR1766470.7788759 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766471.6698630 chr5 175050945 N chr5 175051029 N DUP 46
SRR1766472.2327221 chr5 175050955 N chr5 175051037 N DUP 38
SRR1766447.413892 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766452.6976528 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766457.4840642 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766470.7313587 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766478.6602309 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766484.10286372 chr5 175050944 N chr5 175051028 N DUP 33
SRR1766442.35734643 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766450.5203004 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766461.5058047 chr5 175050945 N chr5 175051029 N DUP 39
SRR1766455.1892458 chr5 175050945 N chr5 175051029 N DUP 34
SRR1766472.39408 chr5 175050945 N chr5 175051029 N DUP 34
SRR1766480.8347342 chr5 175050945 N chr5 175051029 N DUP 34
SRR1766461.7579894 chr5 175050953 N chr5 175051008 N DUP 25
SRR1766451.8483047 chr5 175050944 N chr5 175051028 N DUP 34
SRR1766447.9114426 chr5 175050953 N chr5 175051008 N DUP 24
SRR1766462.9281737 chr5 175050953 N chr5 175051008 N DUP 24
SRR1766466.9559969 chr5 175050953 N chr5 175051008 N DUP 48
SRR1766467.2137023 chr5 175050953 N chr5 175051008 N DUP 30
SRR1766469.8261633 chr5 175050944 N chr5 175051028 N DUP 34
SRR1766474.9737249 chr5 175050944 N chr5 175051028 N DUP 29
SRR1766465.10918318 chr5 175050945 N chr5 175051029 N DUP 47
SRR1766474.3466537 chr5 175050945 N chr5 175051029 N DUP 47
SRR1766461.2177190 chr5 175050945 N chr5 175051029 N DUP 48
SRR1766475.5285578 chr5 175050945 N chr5 175051029 N DUP 48
SRR1766484.7853826 chr5 175050944 N chr5 175051028 N DUP 48
SRR1766486.8999378 chr5 175050945 N chr5 175051029 N DUP 48
SRR1766474.3490832 chr5 175050953 N chr5 175051008 N DUP 48
SRR1766457.579844 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766457.9467093 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766466.11002212 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766461.3594756 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766476.2840754 chr5 175050945 N chr5 175051029 N DUP 49
SRR1766482.5844 chr5 175050953 N chr5 175051008 N DUP 41
SRR1766483.5615626 chr5 175051170 N chr5 175051227 N DEL 12
SRR1766485.11013878 chr4 6660670 N chr4 6660831 N DEL 9
SRR1766463.10813359 chr4 6660608 N chr4 6660664 N DEL 5
SRR1766479.11296806 chr4 6660576 N chr4 6660827 N DUP 5
SRR1766468.2271377 chr4 6660609 N chr4 6660807 N DEL 5
SRR1766481.8242543 chr4 6660783 N chr4 6660866 N DEL 9
SRR1766442.26737790 chr4 6660610 N chr4 6660878 N DEL 3
SRR1766452.9684565 chr4 6660611 N chr4 6660937 N DEL 14
SRR1766482.777608 chr4 6660609 N chr4 6660959 N DEL 4
SRR1766475.10855387 chr4 6660603 N chr4 6660990 N DEL 2
SRR1766453.555705 chr4 6660633 N chr4 6660989 N DEL 2
SRR1766486.5451939 chr4 6660615 N chr4 6660997 N DEL 6
SRR1766448.2424079 chr4 6660615 N chr4 6660997 N DEL 6
SRR1766444.1691075 chr4 6660615 N chr4 6660997 N DEL 6
SRR1766448.5226856 chr16 88672116 N chr16 88672290 N DUP 5
SRR1766444.896964 chr7 2502238 N chr7 2502412 N DEL 8
SRR1766443.3545412 chr7 2502240 N chr7 2502311 N DEL 5
SRR1766442.30452748 chr3 29864960 N chr3 29865259 N DEL 4
SRR1766483.4463568 chr3 29865086 N chr3 29865247 N DEL 8
SRR1766454.7436088 chr3 29864966 N chr3 29865131 N DUP 4
SRR1766471.2666047 chr3 29865016 N chr3 29865170 N DUP 5
SRR1766446.5129797 chr3 29865051 N chr3 29865111 N DEL 9
SRR1766450.1184413 chr3 29865124 N chr3 29865275 N DUP 9
SRR1766482.12279354 chr3 29865037 N chr3 29865141 N DEL 5
SRR1766468.7009829 chr3 29864986 N chr3 29865147 N DEL 8
SRR1766477.5929666 chr3 29865132 N chr3 29865253 N DEL 8
SRR1766446.6575174 chr3 29864976 N chr3 29865263 N DEL 8
SRR1766473.2455928 chr9 65825571 N chr9 65825760 N DEL 13
SRR1766481.8013694 chr9 65825571 N chr9 65825760 N DEL 18
SRR1766455.5832948 chr17 79827460 N chr17 79827583 N DEL 7
SRR1766470.1526337 chr17 79827460 N chr17 79827583 N DEL 12
SRR1766477.6147934 chr17 79827460 N chr17 79827583 N DEL 12
SRR1766455.3741851 chr17 79827499 N chr17 79827604 N DUP 5
SRR1766459.7159435 chr16 89196407 N chr16 89196489 N DEL 3
SRR1766442.2526109 chr16 89196420 N chr16 89196502 N DEL 2
SRR1766446.1917798 chr16 89196419 N chr16 89196501 N DEL 3
SRR1766442.34887238 chr16 89196416 N chr16 89196498 N DEL 6
SRR1766478.6220677 chr16 89196419 N chr16 89196501 N DEL 3
SRR1766468.7190526 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766475.10314943 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766453.5373669 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766468.82812 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766450.6205861 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.8470335 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766470.4308219 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.46260196 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.17570005 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766453.9692498 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.11277883 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766463.7644666 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766442.43724364 chr16 89196502 N chr16 89196608 N DEL 29
SRR1766454.10340797 chr16 89196426 N chr16 89196613 N DEL 10
SRR1766446.2875471 chr14 48710753 N chr14 48710986 N DUP 22
SRR1766450.2967389 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766472.10603905 chr14 48710753 N chr14 48710986 N DUP 23
SRR1766481.2252587 chr14 48710815 N chr14 48710876 N DUP 5
SRR1766474.4587026 chr14 48710863 N chr14 48710946 N DEL 11
SRR1766483.6730716 chr14 48710845 N chr14 48710959 N DEL 19
SRR1766484.3931912 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766462.3532246 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766454.10212117 chr14 48710815 N chr14 48710876 N DUP 5
SRR1766470.3292467 chr14 48710863 N chr14 48710946 N DEL 11
SRR1766463.5167162 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766484.11328190 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766445.5006 chr14 48710815 N chr14 48710876 N DUP 12
SRR1766481.2252587 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766448.3439606 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766476.7842206 chr14 48710753 N chr14 48710904 N DUP 19
SRR1766479.9829555 chr14 48710891 N chr14 48710946 N DEL 3
SRR1766472.5072988 chr14 48710815 N chr14 48710876 N DUP 5
SRR1766473.5600841 chr14 48710891 N chr14 48710946 N DEL 5
SRR1766457.4773511 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766442.36294710 chr14 48710753 N chr14 48710904 N DUP 19
SRR1766457.4441503 chr14 48710863 N chr14 48710946 N DEL 11
SRR1766472.5072988 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766479.13419391 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766470.5542698 chr14 48710815 N chr14 48710876 N DUP 19
SRR1766476.5459174 chr14 48710753 N chr14 48710904 N DUP 19
SRR1766483.6730716 chr14 48710815 N chr14 48710876 N DUP 5
SRR1766448.3881858 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766468.4399353 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766478.689995 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766462.2861715 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766445.4807957 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766471.7338370 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766463.5102635 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766482.383305 chr14 48710815 N chr14 48710876 N DUP 16
SRR1766471.6801776 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766475.11458987 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766466.11132086 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766468.719585 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766457.2583891 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766448.974867 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766442.14276195 chr14 48710753 N chr14 48710876 N DUP 11
SRR1766465.9454850 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766471.2565241 chr14 48710815 N chr14 48710876 N DUP 5
SRR1766454.1977085 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766461.7484242 chr14 48710815 N chr14 48710876 N DUP 10
SRR1766475.496564 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766479.2762163 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766470.3974219 chr14 48710815 N chr14 48710876 N DUP 9
SRR1766457.5768050 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766445.2414144 chr14 48710815 N chr14 48710876 N DUP 8
SRR1766448.5798599 chr14 48710753 N chr14 48710904 N DUP 12
SRR1766484.1647397 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766442.17306690 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766479.7892122 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766443.6859543 chr14 48710753 N chr14 48710986 N DUP 20
SRR1766472.187545 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766454.8148945 chr14 48710815 N chr14 48710876 N DUP 5
SRR1766442.12775010 chr14 48710815 N chr14 48710876 N DUP 5
SRR1766467.3508269 chr14 48710753 N chr14 48710904 N DUP 19
SRR1766442.26609313 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766467.5431639 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766446.3022653 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766442.38357669 chr14 48710753 N chr14 48710811 N DUP 19
SRR1766470.5233128 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766470.1748001 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766480.5891804 chr14 48710815 N chr14 48710876 N DUP 5
SRR1766458.4095278 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766467.5431639 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766481.9557509 chr14 48710753 N chr14 48710814 N DUP 11
SRR1766457.2534100 chr14 48710757 N chr14 48710818 N DUP 11
SRR1766446.7779737 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766474.1258087 chr14 48710782 N chr14 48710840 N DUP 5
SRR1766483.3811038 chr14 48710753 N chr14 48710986 N DUP 24
SRR1766458.3453112 chr14 48710782 N chr14 48710840 N DUP 7
SRR1766469.531006 chr14 48710782 N chr14 48710840 N DUP 10
SRR1766462.8067962 chr14 48710758 N chr14 48710994 N DUP 9
SRR1766457.5768050 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766467.3768663 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766448.2507356 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766442.31012994 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766463.5102635 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766470.5233128 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766483.7327647 chr14 48710845 N chr14 48710959 N DEL 26
SRR1766453.10379217 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766445.3167664 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766460.6129341 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766474.1487035 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766485.2389651 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766468.5267218 chr14 48710814 N chr14 48710959 N DEL 26
SRR1766479.2762163 chr14 48710814 N chr14 48710959 N DEL 25
SRR1766444.107791 chr14 48710784 N chr14 48710960 N DEL 6
SRR1766473.5600841 chr14 48710783 N chr14 48710959 N DEL 15
SRR1766453.9529119 chr14 48710792 N chr14 48710968 N DEL 5
SRR1766480.2668754 chr4 48104393 N chr4 48104685 N DEL 2
SRR1766464.5503426 chr4 48104390 N chr4 48104682 N DEL 3
SRR1766479.11219911 chr4 48104411 N chr4 48104534 N DEL 5
SRR1766468.6160003 chr4 48104399 N chr4 48104652 N DEL 1
SRR1766465.8550235 chr4 48104359 N chr4 48104417 N DUP 7
SRR1766459.5346174 chr4 48104399 N chr4 48104652 N DEL 3
SRR1766449.6067038 chr4 48104431 N chr4 48104684 N DEL 16
SRR1766466.8418436 chr4 48104421 N chr4 48104514 N DEL 18
SRR1766452.9985132 chr4 48104421 N chr4 48104514 N DEL 21
SRR1766451.311775 chr4 48104421 N chr4 48104514 N DEL 22
SRR1766479.11186786 chr4 48104465 N chr4 48104714 N DEL 9
SRR1766464.5030637 chr4 48104368 N chr4 48104462 N DUP 11
SRR1766448.7504018 chr4 48104464 N chr4 48104691 N DEL 17
SRR1766456.6177428 chr4 48104356 N chr4 48104442 N DUP 18
SRR1766450.6373742 chr4 48104464 N chr4 48104691 N DEL 19
SRR1766442.15647221 chr4 48104420 N chr4 48104625 N DEL 23
SRR1766442.32996336 chr4 48104464 N chr4 48104691 N DEL 21
SRR1766476.10020416 chr4 48104420 N chr4 48104625 N DEL 24
SRR1766486.5629839 chr4 48104464 N chr4 48104691 N DEL 24
SRR1766454.1951430 chr4 48104420 N chr4 48104625 N DEL 27
SRR1766451.821205 chr4 48104420 N chr4 48104625 N DEL 28
SRR1766477.5593298 chr4 48104464 N chr4 48104691 N DEL 27
SRR1766453.3320851 chr4 48104464 N chr4 48104691 N DEL 27
SRR1766471.6344989 chr4 48104422 N chr4 48104488 N DEL 9
SRR1766450.9514644 chr4 48104367 N chr4 48104632 N DUP 14
SRR1766470.2954518 chr4 48104422 N chr4 48104488 N DEL 9
SRR1766454.7123705 chr4 48104412 N chr4 48104645 N DUP 9
SRR1766454.6132757 chr4 48104392 N chr4 48104544 N DEL 1
SRR1766452.4658940 chr4 48104365 N chr4 48104651 N DUP 13
SRR1766478.2343450 chr4 48104365 N chr4 48104651 N DUP 18
SRR1766459.2554158 chr4 48104420 N chr4 48104625 N DEL 27
SRR1766481.10027804 chr4 48104420 N chr4 48104625 N DEL 26
SRR1766445.4609705 chr4 48104383 N chr4 48104518 N DUP 12
SRR1766442.26239820 chr4 48104464 N chr4 48104691 N DEL 33
SRR1766442.36144754 chr4 48104464 N chr4 48104691 N DEL 33
SRR1766482.7192643 chr4 48104638 N chr4 48104715 N DUP 10
SRR1766456.1433357 chr4 48104417 N chr4 48104684 N DEL 28
SRR1766456.955390 chr4 48104682 N chr4 48104739 N DUP 20
SRR1766482.3702258 chr4 48104403 N chr4 48104702 N DEL 15
SRR1766482.3483891 chr4 48104436 N chr4 48104691 N DEL 14
SRR1766477.6422413 chr4 48104399 N chr4 48104693 N DEL 11
SRR1766442.24635555 chr4 48104403 N chr4 48104702 N DEL 17
SRR1766468.5239912 chr4 48104403 N chr4 48104702 N DEL 17
SRR1766481.13074124 chr4 48104406 N chr4 48104705 N DEL 12
SRR1766463.9799838 chr4 48104408 N chr4 48104707 N DEL 10
SRR1766476.9873913 chr4 48104635 N chr4 48104703 N DEL 3
SRR1766479.6438310 chr4 48104635 N chr4 48104703 N DEL 3
SRR1766485.2960717 chr4 48104636 N chr4 48104704 N DEL 2
SRR1766471.5996994 chr4 48104399 N chr4 48104733 N DEL 6
SRR1766469.6442650 chr11 86732187 N chr11 86732537 N DEL 2
SRR1766482.1708237 chr11 86732120 N chr11 86732235 N DUP 6
SRR1766478.7668797 chr11 86732120 N chr11 86732235 N DUP 7
SRR1766482.7251140 chr11 86732246 N chr11 86732325 N DUP 7
SRR1766453.3820474 chr11 86732132 N chr11 86732248 N DEL 9
SRR1766442.32012255 chr11 86732135 N chr11 86732251 N DEL 7
SRR1766442.496214 chr11 86732407 N chr11 86732741 N DUP 20
SRR1766461.8010174 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766449.134392 chr17 77562775 N chr17 77562882 N DEL 18
SRR1766472.6600386 chr17 77562838 N chr17 77563008 N DEL 8
SRR1766453.1980992 chr17 77562776 N chr17 77562934 N DUP 10
SRR1766461.1225806 chr17 77562790 N chr17 77562895 N DUP 1
SRR1766449.2517215 chr17 77562775 N chr17 77562882 N DEL 16
SRR1766463.9843627 chr17 77562763 N chr17 77562870 N DEL 10
SRR1766480.7103607 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766481.4453507 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766470.2058659 chr17 77562769 N chr17 77562876 N DEL 10
SRR1766464.9796395 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766477.2284814 chr17 77562763 N chr17 77562870 N DEL 10
SRR1766448.4375654 chr17 77562775 N chr17 77562882 N DEL 15
SRR1766442.12186364 chr17 77562717 N chr17 77562877 N DEL 3
SRR1766453.2539701 chr17 77562716 N chr17 77562876 N DEL 4
SRR1766454.10232245 chr17 77562728 N chr17 77563004 N DEL 6
SRR1766485.7907791 chr7 125569331 N chr7 125569448 N DUP 1
SRR1766443.8109916 chr7 125569331 N chr7 125569448 N DUP 5
SRR1766486.11170887 chr7 125569328 N chr7 125569449 N DUP 7
SRR1766442.28393003 chr7 125569498 N chr7 125569603 N DEL 2
SRR1766471.10707284 chr4 1412089 N chr4 1412150 N DEL 5
SRR1766473.3896575 chr4 1412089 N chr4 1412150 N DEL 5
SRR1766463.2700460 chr4 1412089 N chr4 1412150 N DEL 5
SRR1766482.3322447 chr4 1412089 N chr4 1412150 N DEL 5
SRR1766467.725646 chr4 1412089 N chr4 1412150 N DEL 5
SRR1766451.9203647 chr4 1412089 N chr4 1412150 N DEL 5
SRR1766471.7885683 chr4 1412089 N chr4 1412150 N DEL 5
SRR1766456.6422111 chr4 1412089 N chr4 1412210 N DEL 5
SRR1766447.2968816 chr4 1412089 N chr4 1412210 N DEL 5
SRR1766476.1470523 chr4 1412145 N chr4 1412206 N DEL 5
SRR1766460.5915513 chr4 1412115 N chr4 1412174 N DUP 5
SRR1766477.5833728 chrY 11027124 N chrY 11027215 N DEL 11
SRR1766484.2408070 chr2 203206997 N chr2 203207154 N DEL 3
SRR1766460.7628273 chr2 203206997 N chr2 203207154 N DEL 5
SRR1766478.7868750 chr2 203206999 N chr2 203207076 N DEL 5
SRR1766485.12001774 chr2 203206999 N chr2 203207076 N DEL 8
SRR1766462.10109056 chr2 203207020 N chr2 203207095 N DUP 5
SRR1766469.8495504 chr2 203207140 N chr2 203207374 N DEL 9
SRR1766474.3526728 chr2 203207076 N chr2 203207155 N DUP 3
SRR1766462.7164651 chr2 203207007 N chr2 203207164 N DEL 5
SRR1766456.4422699 chr2 203207094 N chr2 203207175 N DEL 5
SRR1766475.383348 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766480.6669082 chr6 106542757 N chr6 106543132 N DEL 8
SRR1766464.10825663 chr6 106543004 N chr6 106543386 N DEL 5
SRR1766479.6208372 chr6 106543004 N chr6 106543386 N DEL 5
SRR1766464.5401786 chr6 106543028 N chr6 106543410 N DEL 4
SRR1766462.11093355 chr6 106542757 N chr6 106543137 N DEL 2
SRR1766481.23690 chr6 106542757 N chr6 106543132 N DEL 3
SRR1766480.8268083 chr6 106542757 N chr6 106543137 N DEL 9
SRR1766454.9040902 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766484.5579563 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766443.7825574 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766484.1915601 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766450.8357767 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766480.6669082 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766442.4901217 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766446.4301961 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766486.2854498 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766484.4024732 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766482.3149900 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766455.1044501 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766474.2176121 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766482.6394426 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766447.8510608 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766477.1943205 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766442.38150251 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766454.1763559 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766454.6799396 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766452.8968949 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766484.1915601 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766446.9023220 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766442.9013655 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766467.9667718 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766453.10777787 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766477.4797036 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766482.282476 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766461.8985552 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766463.1766339 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766459.165027 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766442.28691290 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766475.1115337 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766451.9399581 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766450.1020368 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766456.6118378 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766442.8908181 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766457.3041478 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766474.8798753 chr6 106542757 N chr6 106543132 N DEL 10
SRR1766460.6682335 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766473.5338326 chr6 106542757 N chr6 106543137 N DEL 15
SRR1766481.2458626 chr6 106542759 N chr6 106543134 N DEL 10
SRR1766443.1400077 chr6 106542760 N chr6 106543135 N DEL 10
SRR1766485.9907970 chr6 106542769 N chr6 106543144 N DEL 3
SRR1766443.1655505 chr6 106542769 N chr6 106543144 N DEL 3
SRR1766459.5064670 chr6 106542770 N chr6 106543145 N DEL 2
SRR1766446.7998013 chr6 106542773 N chr6 106543183 N DEL 4
SRR1766448.5757365 chr6 106542773 N chr6 106543183 N DEL 4
SRR1766475.974681 chr6 106542776 N chr6 106543186 N DEL 1
SRR1766443.2010814 chr6 106542847 N chr6 106543229 N DEL 5
SRR1766442.9721449 chr6 106542847 N chr6 106543229 N DEL 5
SRR1766442.35302490 chr6 106542847 N chr6 106543229 N DEL 5
SRR1766442.375974 chr6 106542987 N chr6 106543367 N DUP 1
SRR1766483.9491190 chr2 57548080 N chr2 57548145 N DUP 11
SRR1766463.4045534 chr2 57548108 N chr2 57548161 N DEL 51
SRR1766477.9656294 chr2 57548108 N chr2 57548161 N DEL 29
SRR1766442.19056028 chr2 57548108 N chr2 57548161 N DEL 27
SRR1766470.6887218 chr2 57548108 N chr2 57548161 N DEL 24
SRR1766448.6682300 chr2 57548108 N chr2 57548161 N DEL 17
SRR1766482.7022931 chr2 57548066 N chr2 57548178 N DEL 5
SRR1766477.791051 chr2 57548069 N chr2 57548181 N DEL 5
SRR1766469.9087748 chrX 136451023 N chrX 136451222 N DUP 5
SRR1766469.4726991 chrX 136451242 N chrX 136451293 N DUP 5
SRR1766463.326785 chrX 136451242 N chrX 136451293 N DUP 5
SRR1766454.6806192 chrX 136451176 N chrX 136451305 N DUP 19
SRR1766462.10334310 chrX 136451220 N chrX 136451269 N DUP 21
SRR1766458.8746635 chrX 136451149 N chrX 136451220 N DEL 14
SRR1766464.8944529 chrX 136451220 N chrX 136451269 N DUP 19
SRR1766443.1096536 chrX 136451149 N chrX 136451220 N DEL 14
SRR1766449.7977451 chrX 136451114 N chrX 136451303 N DUP 18
SRR1766461.361617 chrX 136451222 N chrX 136451295 N DUP 12
SRR1766455.7313870 chrX 136451258 N chrX 136451319 N DUP 13
SRR1766442.43014644 chrX 136451145 N chrX 136451256 N DEL 18
SRR1766472.8105755 chrX 136451145 N chrX 136451256 N DEL 17
SRR1766456.952375 chrX 136451145 N chrX 136451256 N DEL 16
SRR1766451.6994936 chr5 180296973 N chr5 180297076 N DEL 8
SRR1766467.6367734 chr5 180296973 N chr5 180297076 N DEL 8
SRR1766477.8076387 chr5 180296973 N chr5 180297076 N DEL 8
SRR1766451.5315885 chr5 180297012 N chr5 180297105 N DEL 24
SRR1766486.800966 chr5 180296973 N chr5 180297076 N DEL 8
SRR1766472.5620055 chr5 180297012 N chr5 180297105 N DEL 23
SRR1766475.6730123 chr5 180296980 N chr5 180297083 N DEL 9
SRR1766451.9477798 chr5 180297004 N chr5 180297107 N DEL 1
SRR1766484.7177136 chr5 180297004 N chr5 180297107 N DEL 1
SRR1766446.8654432 chr5 180297008 N chr5 180297111 N DEL 1
SRR1766445.3010205 chr5 180297008 N chr5 180297111 N DEL 1
SRR1766463.7868411 chr5 180297014 N chr5 180297105 N DEL 19
SRR1766474.1965311 chr5 180297010 N chr5 180297113 N DEL 1
SRR1766450.8133446 chr5 180296924 N chr5 180297117 N DEL 3
SRR1766449.7751472 chr1 143258312 N chr1 143258458 N DUP 12
SRR1766462.5000713 chr1 143258260 N chr1 143258335 N DEL 5
SRR1766480.2207946 chr9 19434255 N chr9 19434449 N DEL 5
SRR1766483.2285478 chr9 19434284 N chr9 19434476 N DUP 5
SRR1766444.6093577 chr9 19434264 N chr9 19434341 N DEL 5
SRR1766471.5914594 chr9 19434298 N chr9 19434455 N DEL 3
SRR1766460.11155852 chr9 19434273 N chr9 19434467 N DEL 5
SRR1766442.3777574 chr9 19434223 N chr9 19434496 N DEL 1
SRR1766462.7149598 chr16 7229912 N chr16 7230179 N DUP 25
SRR1766452.2071920 chr16 7229912 N chr16 7230179 N DUP 25
SRR1766453.10549147 chr16 7230002 N chr16 7230179 N DUP 20
SRR1766458.9142567 chr16 7229929 N chr16 7230002 N DEL 5
SRR1766475.10773090 chr16 7229895 N chr16 7230004 N DEL 13
SRR1766452.9703534 chr16 7230042 N chr16 7230097 N DEL 5
SRR1766478.9213620 chr16 7230025 N chr16 7230080 N DEL 5
SRR1766460.1739809 chr16 7230117 N chr16 7230170 N DUP 5
SRR1766464.21270 chr16 7229935 N chr16 7230204 N DEL 5
SRR1766445.7225047 chr16 7229935 N chr16 7230204 N DEL 5
SRR1766453.2802284 chr16 7229750 N chr16 7230204 N DEL 5
SRR1766470.7208139 chr16 7229863 N chr16 7230208 N DEL 6
SRR1766443.3863348 chr16 7229798 N chr16 7230210 N DEL 5
SRR1766455.8383980 chr16 7229801 N chr16 7230213 N DEL 5
SRR1766442.37383857 chr16 7229803 N chr16 7230215 N DEL 4
SRR1766471.7267974 chr16 7229803 N chr16 7230215 N DEL 4
SRR1766449.5409877 chr14 89567530 N chr14 89567663 N DEL 5
SRR1766471.8222310 chr14 89567530 N chr14 89567663 N DEL 5
SRR1766468.4869278 chr14 89567530 N chr14 89567663 N DEL 5
SRR1766475.9081550 chr14 89567530 N chr14 89567663 N DEL 5
SRR1766477.5389434 chr14 89567530 N chr14 89567663 N DEL 5
SRR1766482.4017194 chr14 89567530 N chr14 89567663 N DEL 5
SRR1766474.4227927 chr14 89567556 N chr14 89567720 N DUP 7
SRR1766461.1387860 chr14 89567556 N chr14 89567720 N DUP 8
SRR1766475.306879 chr14 89567556 N chr14 89567720 N DUP 13
SRR1766442.1922502 chr14 89567556 N chr14 89567720 N DUP 27
SRR1766473.6022383 chr14 89567556 N chr14 89567654 N DUP 27
SRR1766460.9566402 chr14 89567589 N chr14 89567654 N DUP 30
SRR1766449.3225221 chr14 89567589 N chr14 89567654 N DUP 30
SRR1766449.4399257 chr14 89567556 N chr14 89567654 N DUP 25
SRR1766454.6520794 chr14 89567556 N chr14 89567654 N DUP 25
SRR1766458.3737403 chr14 89567556 N chr14 89567654 N DUP 25
SRR1766442.43692910 chr14 89567621 N chr14 89567688 N DEL 30
SRR1766458.8628337 chr15 55926122 N chr15 55926203 N DUP 3
SRR1766484.10906861 chr15 55926115 N chr15 55926216 N DUP 5
SRR1766443.221338 chr15 55926115 N chr15 55926216 N DUP 5
SRR1766468.5221580 chr15 55926115 N chr15 55926216 N DUP 5
SRR1766478.11494322 chr15 55926129 N chr15 55926232 N DEL 1
SRR1766442.43901911 chr6 22836799 N chr6 22836928 N DEL 10
SRR1766443.5421022 chr6 22836800 N chr6 22836929 N DEL 5
SRR1766461.1534938 chr6 22836945 N chr6 22837373 N DEL 6
SRR1766451.2477563 chr6 22836918 N chr6 22837221 N DUP 5
SRR1766457.769618 chr6 22837027 N chr6 22837377 N DEL 10
SRR1766474.6762309 chr6 22836737 N chr6 22837089 N DUP 10
SRR1766482.12278866 chr6 22836769 N chr6 22837121 N DUP 1
SRR1766483.6957947 chr6 22836780 N chr6 22837036 N DEL 3
SRR1766447.1367030 chr6 22836755 N chr6 22837060 N DEL 9
SRR1766456.6461724 chr6 22836863 N chr6 22837341 N DEL 5
SRR1766444.1238974 chr6 22837027 N chr6 22837377 N DEL 5
SRR1766467.8717218 chr6 22836899 N chr6 22837377 N DEL 5
SRR1766466.3864747 chr6 22836899 N chr6 22837377 N DEL 5
SRR1766477.11342266 chr6 22836908 N chr6 22837386 N DEL 5
SRR1766463.6793580 chr6 22836784 N chr6 22837389 N DEL 3
SRR1766484.8161991 chr6 22836830 N chr6 22837435 N DEL 5
SRR1766450.3228494 chr6 22836833 N chr6 22837438 N DEL 5
SRR1766471.9581985 chr6 22837326 N chr6 22837454 N DEL 1
SRR1766465.10260035 chr6 8403466 N chr6 8403567 N DEL 1
SRR1766481.7561205 chr11 2042289 N chr11 2042380 N DEL 5
SRR1766465.6558305 chr11 2042240 N chr11 2042386 N DEL 7
SRR1766460.1538195 chr14 73023400 N chr14 73023455 N DEL 6
SRR1766442.31154963 chr14 73023333 N chr14 73023471 N DUP 9
SRR1766473.7352866 chr14 73023364 N chr14 73023473 N DUP 10
SRR1766484.7356431 chr14 73023333 N chr14 73023471 N DUP 12
SRR1766451.1833916 chr14 73023333 N chr14 73023471 N DUP 13
SRR1766475.449926 chr14 73023333 N chr14 73023471 N DUP 13
SRR1766442.34510338 chr14 73023333 N chr14 73023471 N DUP 15
SRR1766448.9732904 chr14 73023333 N chr14 73023471 N DUP 17
SRR1766484.7564148 chr14 73023400 N chr14 73023455 N DEL 17
SRR1766444.2549652 chr14 73023401 N chr14 73023454 N DUP 13
SRR1766469.5986209 chr14 73023401 N chr14 73023454 N DUP 13
SRR1766483.1305459 chr14 73023401 N chr14 73023454 N DUP 13
SRR1766464.9278956 chr14 73023401 N chr14 73023454 N DUP 15
SRR1766463.7845313 chr14 73023401 N chr14 73023454 N DUP 15
SRR1766446.7593408 chr14 73023401 N chr14 73023454 N DUP 15
SRR1766443.9294079 chr14 73023401 N chr14 73023454 N DUP 15
SRR1766464.880577 chr14 73023333 N chr14 73023525 N DUP 4
SRR1766446.1327521 chr14 73023400 N chr14 73023455 N DEL 15
SRR1766446.7965769 chr14 73023400 N chr14 73023455 N DEL 15
SRR1766442.22081457 chr14 73023400 N chr14 73023455 N DEL 15
SRR1766458.1247687 chr14 73023400 N chr14 73023455 N DEL 15
SRR1766447.6500876 chr14 73023400 N chr14 73023455 N DEL 14
SRR1766452.3441462 chr14 73023400 N chr14 73023455 N DEL 13
SRR1766472.976719 chr14 73023387 N chr14 73023469 N DEL 1
SRR1766456.2016791 chr14 73023347 N chr14 73023539 N DEL 9
SRR1766456.4352145 chr14 73023347 N chr14 73023539 N DEL 9
SRR1766469.4768275 chr14 73023379 N chr14 73023542 N DEL 9
SRR1766442.31733825 chr12 124416670 N chr12 124416722 N DUP 6
SRR1766457.4836368 chr12 124416701 N chr12 124416880 N DEL 16
SRR1766462.6891396 chr12 124416670 N chr12 124416758 N DUP 5
SRR1766476.4800941 chr12 124416743 N chr12 124416957 N DEL 10
SRR1766480.7016293 chr6 47015895 N chr6 47016044 N DUP 2
SRR1766454.4652776 chr5 142075334 N chr5 142075517 N DEL 5
SRR1766461.3752135 chr5 142075334 N chr5 142075517 N DEL 5
SRR1766465.9171882 chr5 142075359 N chr5 142075542 N DEL 3
SRR1766485.4578163 chr5 142075394 N chr5 142075878 N DEL 5
SRR1766448.321931 chr5 142075359 N chr5 142075542 N DEL 7
SRR1766448.8697066 chr5 142075359 N chr5 142075542 N DEL 3
SRR1766452.4302792 chr5 142075446 N chr5 142075623 N DUP 14
SRR1766467.5489135 chr5 142075495 N chr5 142076377 N DEL 5
SRR1766456.5769900 chr5 142075513 N chr5 142075792 N DUP 4
SRR1766473.9003948 chr5 142075511 N chr5 142076518 N DUP 5
SRR1766446.9078262 chr5 142075507 N chr5 142076514 N DUP 5
SRR1766458.5423 chr5 142075507 N chr5 142075635 N DUP 5
SRR1766458.8424448 chr5 142075507 N chr5 142075635 N DUP 5
SRR1766482.4457438 chr5 142075413 N chr5 142075518 N DEL 4
SRR1766483.3363944 chr5 142075778 N chr5 142076052 N DUP 9
SRR1766473.3496839 chr5 142075436 N chr5 142075613 N DUP 5
SRR1766476.1934713 chr5 142075584 N chr5 142076060 N DUP 5
SRR1766446.1260415 chr5 142075632 N chr5 142075932 N DEL 5
SRR1766472.7189654 chr5 142075576 N chr5 142075779 N DEL 2
SRR1766474.438999 chr5 142075576 N chr5 142075779 N DEL 1
SRR1766471.10491058 chr5 142075446 N chr5 142075623 N DUP 3
SRR1766478.11736947 chr5 142075446 N chr5 142075623 N DUP 5
SRR1766484.4528833 chr5 142075637 N chr5 142075937 N DEL 10
SRR1766480.7340283 chr5 142075637 N chr5 142075937 N DEL 10
SRR1766472.4059986 chr5 142075627 N chr5 142076458 N DEL 5
SRR1766473.2427472 chr5 142075634 N chr5 142076465 N DEL 5
SRR1766449.4389187 chr5 142075666 N chr5 142076546 N DEL 5
SRR1766474.5598418 chr5 142075654 N chr5 142075757 N DEL 5
SRR1766460.8835584 chr5 142075666 N chr5 142076093 N DEL 5
SRR1766472.6419271 chr5 142075446 N chr5 142075623 N DUP 10
SRR1766473.1898952 chr5 142075656 N chr5 142075759 N DEL 5
SRR1766468.2833133 chr5 142075664 N chr5 142075965 N DEL 11
SRR1766475.2519650 chr5 142075666 N chr5 142075868 N DEL 4
SRR1766442.13700379 chr5 142075662 N chr5 142075962 N DEL 11
SRR1766467.10704287 chr5 142075767 N chr5 142076495 N DUP 13
SRR1766462.3291751 chr5 142075473 N chr5 142075650 N DUP 9
SRR1766456.3761382 chr5 142075461 N chr5 142075589 N DEL 3
SRR1766460.5921866 chr5 142075615 N chr5 142075714 N DUP 1
SRR1766454.5424195 chr5 142075406 N chr5 142075640 N DEL 3
SRR1766465.1585521 chr5 142075668 N chr5 142075770 N DUP 7
SRR1766461.3811885 chr5 142075724 N chr5 142075823 N DUP 12
SRR1766482.11441581 chr5 142075690 N chr5 142076521 N DEL 2
SRR1766442.23039326 chr5 142075621 N chr5 142075724 N DEL 12
SRR1766473.9003948 chr5 142075621 N chr5 142075724 N DEL 12
SRR1766448.1539612 chr5 142075629 N chr5 142075731 N DEL 11
SRR1766461.3811885 chr5 142075724 N chr5 142075823 N DUP 18
SRR1766473.6757673 chr5 142075722 N chr5 142075774 N DEL 13
SRR1766464.4547729 chr5 142075440 N chr5 142075725 N DEL 16
SRR1766479.5747455 chr5 142075460 N chr5 142075688 N DEL 1
SRR1766458.4332305 chr5 142075715 N chr5 142075767 N DEL 18
SRR1766481.4728186 chr5 142075767 N chr5 142075817 N DUP 4
SRR1766478.4332944 chr5 142075421 N chr5 142075757 N DEL 11
SRR1766450.4901598 chr5 142075763 N chr5 142076311 N DUP 9
SRR1766451.9203540 chr5 142075437 N chr5 142075865 N DUP 12
SRR1766452.9835353 chr5 142075493 N chr5 142075774 N DEL 2
SRR1766460.5641364 chr5 142075671 N chr5 142075872 N DEL 9
SRR1766447.7767453 chr5 142075509 N chr5 142075936 N DUP 2
SRR1766448.8697066 chr5 142075434 N chr5 142075867 N DEL 16
SRR1766473.10887337 chr5 142075434 N chr5 142075867 N DEL 16
SRR1766469.3578124 chr5 142075434 N chr5 142075867 N DEL 16
SRR1766476.1049434 chr5 142075435 N chr5 142075868 N DEL 14
SRR1766483.3797013 chr5 142075473 N chr5 142075951 N DEL 1
SRR1766442.20535769 chr5 142075417 N chr5 142075950 N DEL 2
SRR1766452.832518 chr5 142075415 N chr5 142075948 N DEL 4
SRR1766456.3761382 chr5 142075484 N chr5 142075962 N DEL 5
SRR1766469.3578124 chr5 142075507 N chr5 142075983 N DUP 10
SRR1766444.4694678 chr5 142075485 N chr5 142075963 N DEL 5
SRR1766476.2082872 chr5 142075991 N chr5 142076344 N DUP 5
SRR1766482.2601077 chr5 142075610 N chr5 142076011 N DEL 16
SRR1766471.2889692 chr5 142075610 N chr5 142076011 N DEL 16
SRR1766471.10882051 chr5 142075510 N chr5 142076113 N DUP 4
SRR1766456.5633708 chr5 142076113 N chr5 142076290 N DEL 5
SRR1766481.10070634 chr5 142075461 N chr5 142076113 N DUP 1
SRR1766460.8244418 chr5 142075461 N chr5 142076113 N DUP 5
SRR1766442.40426246 chr5 142075461 N chr5 142076113 N DUP 5
SRR1766485.9762040 chr5 142075756 N chr5 142076128 N DUP 10
SRR1766465.9802791 chr5 142075461 N chr5 142076113 N DUP 5
SRR1766474.438999 chr5 142075461 N chr5 142076113 N DUP 5
SRR1766460.10172022 chr5 142075461 N chr5 142076113 N DUP 5
SRR1766462.8520247 chr5 142075461 N chr5 142076113 N DUP 5
SRR1766442.15328908 chr5 142076113 N chr5 142076469 N DEL 5
SRR1766472.4059986 chr5 142075937 N chr5 142076112 N DUP 5
SRR1766457.328021 chr5 142075757 N chr5 142076129 N DUP 5
SRR1766446.7746122 chr5 142075937 N chr5 142076112 N DUP 5
SRR1766450.3596382 chr5 142075621 N chr5 142076144 N DUP 1
SRR1766461.7536071 chr5 142075348 N chr5 142076045 N DEL 2
SRR1766474.8456588 chr5 142075868 N chr5 142076142 N DUP 7
SRR1766450.10488860 chr5 142075765 N chr5 142076137 N DUP 5
SRR1766442.7403132 chr5 142076148 N chr5 142076377 N DEL 5
SRR1766442.28041839 chr5 142075446 N chr5 142076098 N DUP 5
SRR1766455.13450 chr5 142075480 N chr5 142076085 N DEL 5
SRR1766452.2516129 chr5 142075336 N chr5 142076207 N DUP 2
SRR1766454.10761406 chr5 142076148 N chr5 142076377 N DEL 5
SRR1766445.1884119 chr5 142075488 N chr5 142075966 N DEL 5
SRR1766484.170228 chr5 142075498 N chr5 142075976 N DEL 1
SRR1766480.7340283 chr5 142076203 N chr5 142076430 N DUP 5
SRR1766462.2882869 chr5 142076099 N chr5 142076377 N DEL 10
SRR1766471.7055014 chr5 142075635 N chr5 142076060 N DUP 7
SRR1766442.20535769 chr5 142075651 N chr5 142076354 N DEL 5
SRR1766465.9802791 chr5 142075421 N chr5 142076307 N DEL 6
SRR1766469.4624370 chr5 142076328 N chr5 142076377 N DUP 1
SRR1766446.212741 chr5 142076099 N chr5 142076327 N DEL 14
SRR1766474.10339830 chr5 142076099 N chr5 142076327 N DEL 9
SRR1766483.4753866 chr5 142076099 N chr5 142076327 N DEL 13
SRR1766470.7552634 chr5 142075500 N chr5 142076332 N DEL 5
SRR1766462.3291751 chr5 142075495 N chr5 142076377 N DEL 8
SRR1766465.2076561 chr5 142075605 N chr5 142075956 N DEL 10
SRR1766465.8121722 chr5 142075605 N chr5 142076484 N DUP 7
SRR1766484.1089274 chr5 142075605 N chr5 142076484 N DUP 3
SRR1766455.13450 chr5 142075482 N chr5 142076413 N DEL 5
SRR1766484.170228 chr5 142075465 N chr5 142076521 N DUP 2
SRR1766460.1780949 chr5 142075603 N chr5 142075757 N DEL 10
SRR1766466.661031 chr5 142076060 N chr5 142076465 N DEL 5
SRR1766450.3596382 chr5 142076060 N chr5 142076465 N DEL 5
SRR1766442.25418342 chr5 142076060 N chr5 142076465 N DEL 5
SRR1766481.10070634 chr5 142076060 N chr5 142076465 N DEL 5
SRR1766465.5207115 chr5 142075932 N chr5 142076560 N DUP 7
SRR1766464.10276757 chr5 142076289 N chr5 142076565 N DUP 5
SRR1766474.10339830 chr5 142075460 N chr5 142076565 N DUP 8
SRR1766477.8689244 chr5 142075474 N chr5 142076579 N DUP 6
SRR1766446.8048790 chr5 142076074 N chr5 142076479 N DEL 1
SRR1766442.38971932 chr5 142075587 N chr5 142076565 N DUP 4
SRR1766468.2803002 chr5 142075587 N chr5 142076565 N DUP 4
SRR1766447.9653765 chr5 142076331 N chr5 142076509 N DEL 5
SRR1766452.3788665 chr5 142075802 N chr5 142076580 N DEL 11
SRR1766469.718674 chr5 142075621 N chr5 142076552 N DEL 5
SRR1766464.889417 chr5 142075655 N chr5 142076584 N DEL 5
SRR1766450.5226772 chr2 240357809 N chr2 240357930 N DEL 17
SRR1766461.6529098 chr2 240357803 N chr2 240357936 N DEL 7
SRR1766445.5948862 chr2 240357804 N chr2 240357937 N DEL 7
SRR1766471.10069641 chr2 240357805 N chr2 240357938 N DEL 7
SRR1766467.4026215 chr2 240357802 N chr2 240357939 N DEL 6
SRR1766479.11882484 chr2 240357802 N chr2 240357939 N DEL 6
SRR1766467.5742111 chr2 240357804 N chr2 240357941 N DEL 4
SRR1766470.6801985 chr2 240357803 N chr2 240357944 N DEL 1
SRR1766452.5059440 chr6 41225575 N chr6 41225658 N DEL 1
SRR1766473.6339450 chr19 57019888 N chr19 57020218 N DUP 5
SRR1766486.10854292 chr12 122731874 N chr12 122732098 N DUP 14
SRR1766461.9885243 chr19 28114274 N chr19 28114347 N DEL 3
SRR1766458.1877385 chr19 28114274 N chr19 28114347 N DEL 5
SRR1766461.8102491 chr19 28114274 N chr19 28114347 N DEL 5
SRR1766461.3248928 chr19 28114274 N chr19 28114347 N DEL 5
SRR1766443.202890 chr19 28114314 N chr19 28114373 N DEL 3
SRR1766466.1350973 chr19 28114314 N chr19 28114373 N DEL 3
SRR1766459.11200037 chr19 28114323 N chr19 28114386 N DUP 17
SRR1766445.3464747 chr19 28114323 N chr19 28114386 N DUP 16
SRR1766479.6448928 chr19 28114241 N chr19 28114332 N DEL 6
SRR1766442.15591530 chr19 28114189 N chr19 28114337 N DEL 1
SRR1766450.2247666 chr19 28114244 N chr19 28114335 N DEL 3
SRR1766477.11694658 chr19 28114306 N chr19 28114395 N DEL 5
SRR1766469.3925652 chr19 28114303 N chr19 28114392 N DEL 8
SRR1766471.11539526 chr19 28114309 N chr19 28114398 N DEL 3
SRR1766465.4292348 chr8 116297695 N chr8 116297929 N DEL 12
SRR1766462.6420849 chr10 129070543 N chr10 129070709 N DUP 5
SRR1766484.8976712 chr10 75334163 N chr10 75334280 N DEL 5
SRR1766475.4128280 chr10 75333993 N chr10 75334110 N DEL 5
SRR1766460.9971632 chr10 75333993 N chr10 75334110 N DEL 2
SRR1766472.9166088 chr6 166955879 N chr6 166956030 N DEL 11
SRR1766483.8043546 chr2 239658804 N chr2 239659225 N DEL 5
SRR1766463.2727969 chr18 78839149 N chr18 78839218 N DUP 5
SRR1766479.6494928 chr18 78839036 N chr18 78839205 N DUP 7
SRR1766475.10800441 chr20 30292124 N chr20 30292395 N DUP 3
SRR1766452.4826438 chr9 85647606 N chr9 85647718 N DEL 5
SRR1766454.6063548 chr7 51827451 N chr7 51827502 N DUP 5
SRR1766454.9405089 chr15 57278879 N chr15 57278941 N DEL 5
SRR1766442.41158297 chr14 86443411 N chr14 86443576 N DEL 2
SRR1766482.4923603 chr14 86443411 N chr14 86443576 N DEL 6
SRR1766450.7533808 chr14 86443422 N chr14 86443494 N DEL 8
SRR1766470.347213 chr14 86443422 N chr14 86443494 N DEL 14
SRR1766475.9134706 chr14 86443422 N chr14 86443494 N DEL 20
SRR1766465.9250892 chr14 86443422 N chr14 86443494 N DEL 25
SRR1766460.8005540 chr14 86443460 N chr14 86443513 N DUP 24
SRR1766466.10372861 chr14 86443460 N chr14 86443513 N DUP 27
SRR1766463.2018673 chr14 86443460 N chr14 86443552 N DUP 41
SRR1766472.8052251 chr14 86443460 N chr14 86443552 N DUP 37
SRR1766442.7367609 chr14 86443460 N chr14 86443513 N DUP 33
SRR1766442.28998354 chr14 86443476 N chr14 86443573 N DUP 32
SRR1766442.21800567 chr14 86443460 N chr14 86443584 N DUP 45
SRR1766466.2280465 chr14 86443478 N chr14 86443548 N DUP 9
SRR1766470.1719124 chr14 86443478 N chr14 86443548 N DUP 9
SRR1766486.5411664 chr14 86443460 N chr14 86443513 N DUP 34
SRR1766452.10667945 chr14 86443460 N chr14 86443584 N DUP 41
SRR1766481.12920665 chr14 86443460 N chr14 86443513 N DUP 35
SRR1766448.2943442 chr14 86443460 N chr14 86443584 N DUP 36
SRR1766452.6550543 chr14 86443478 N chr14 86443548 N DUP 31
SRR1766470.5723466 chr14 86443460 N chr14 86443584 N DUP 36
SRR1766463.6288637 chr14 86443460 N chr14 86443584 N DUP 35
SRR1766475.4870310 chr14 86443478 N chr14 86443548 N DUP 30
SRR1766442.34630070 chr14 86443460 N chr14 86443513 N DUP 26
SRR1766474.2676307 chr14 86443460 N chr14 86443513 N DUP 48
SRR1766461.11011897 chr14 86443478 N chr14 86443548 N DUP 30
SRR1766470.611993 chr14 86443478 N chr14 86443548 N DUP 33
SRR1766442.7954196 chr14 86443478 N chr14 86443548 N DUP 34
SRR1766459.6923307 chr14 86443478 N chr14 86443548 N DUP 28
SRR1766467.7149342 chr14 86443460 N chr14 86443513 N DUP 23
SRR1766460.2752859 chr14 86443478 N chr14 86443548 N DUP 24
SRR1766464.2892468 chr14 86443478 N chr14 86443548 N DUP 25
SRR1766442.38756996 chr14 86443635 N chr14 86443737 N DEL 2
SRR1766484.2829057 chr14 86443635 N chr14 86443737 N DEL 3
SRR1766486.605216 chr14 86443635 N chr14 86443737 N DEL 4
SRR1766461.2890768 chr14 86443416 N chr14 86443576 N DEL 4
SRR1766481.9530921 chr14 86443487 N chr14 86443547 N DEL 3
SRR1766477.11133941 chr14 86443635 N chr14 86443737 N DEL 17
SRR1766457.8113491 chr14 86443635 N chr14 86443737 N DEL 17
SRR1766442.42952005 chr14 86443635 N chr14 86443737 N DEL 17
SRR1766454.1807925 chr14 86443635 N chr14 86443737 N DEL 29
SRR1766478.5238000 chr14 86443435 N chr14 86443685 N DEL 18
SRR1766462.2928365 chr14 86443577 N chr14 86443685 N DEL 22
SRR1766461.3674012 chr14 86443635 N chr14 86443737 N DEL 34
SRR1766483.3498350 chr14 86443635 N chr14 86443737 N DEL 34
SRR1766486.3612478 chr14 86443635 N chr14 86443737 N DEL 34
SRR1766483.407243 chr14 86443438 N chr14 86443688 N DEL 12
SRR1766450.8836247 chr14 86443661 N chr14 86443737 N DEL 16
SRR1766442.22992507 chr14 86443691 N chr14 86443767 N DEL 16
SRR1766479.4639488 chr14 86443661 N chr14 86443737 N DEL 11
SRR1766459.3077224 chr14 86443661 N chr14 86443737 N DEL 11
SRR1766463.349530 chr14 86443635 N chr14 86443737 N DEL 20
SRR1766474.8929750 chr14 86443661 N chr14 86443737 N DEL 11
SRR1766448.10153681 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766471.4194 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766449.8655581 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766454.4271292 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766473.9157197 chr14 86443753 N chr14 86443833 N DUP 40
SRR1766473.5821116 chr14 86443753 N chr14 86443833 N DUP 40
SRR1766482.7644767 chr14 86443753 N chr14 86443833 N DUP 39
SRR1766473.751926 chr14 86443763 N chr14 86443844 N DUP 24
SRR1766481.7212995 chr14 86443785 N chr14 86443840 N DEL 5
SRR1766473.8607299 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766452.7161305 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766485.2079904 chr14 86443785 N chr14 86443840 N DEL 5
SRR1766450.1632911 chr14 86443785 N chr14 86443840 N DEL 5
SRR1766482.5713540 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766469.2243889 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766484.2829057 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766442.24853383 chr14 86443813 N chr14 86443868 N DEL 15
SRR1766455.6036295 chr14 86443927 N chr14 86443999 N DUP 1
SRR1766469.783017 chr14 86443927 N chr14 86443999 N DUP 3
SRR1766478.6412690 chr14 86443927 N chr14 86443999 N DUP 3
SRR1766461.2890768 chr14 86443841 N chr14 86444015 N DUP 5
SRR1766477.11133941 chr14 86443841 N chr14 86444015 N DUP 5
SRR1766446.8464311 chr14 86443841 N chr14 86444015 N DUP 5
SRR1766471.11571761 chr14 86443841 N chr14 86444015 N DUP 5
SRR1766472.8052251 chr14 86443841 N chr14 86444015 N DUP 5
SRR1766481.9530921 chr14 86443841 N chr14 86444015 N DUP 5
SRR1766442.27934969 chr14 86443841 N chr14 86444015 N DUP 5
SRR1766478.5238000 chr14 86443841 N chr14 86444015 N DUP 5
SRR1766478.6937671 chr14 86444045 N chr14 86444143 N DEL 9
SRR1766451.2672792 chr14 86444057 N chr14 86444117 N DEL 15
SRR1766442.22992507 chr14 86444057 N chr14 86444117 N DEL 16
SRR1766463.349530 chr14 86443590 N chr14 86444058 N DUP 16
SRR1766454.2140418 chr14 86444059 N chr14 86444112 N DEL 16
SRR1766483.3498350 chr14 86444059 N chr14 86444112 N DEL 16
SRR1766476.939331 chr14 86444059 N chr14 86444112 N DEL 20
SRR1766455.6272504 chr14 86444085 N chr14 86444144 N DEL 7
SRR1766456.1128338 chr14 86444085 N chr14 86444144 N DEL 8
SRR1766472.10019288 chr14 86444085 N chr14 86444144 N DEL 8
SRR1766473.9157197 chr14 86443397 N chr14 86444095 N DUP 10
SRR1766470.2305340 chr14 86444059 N chr14 86444112 N DEL 23
SRR1766464.4151464 chr14 86444059 N chr14 86444112 N DEL 27
SRR1766442.7259017 chr14 86444059 N chr14 86444112 N DEL 33
SRR1766442.30329864 chr14 86444059 N chr14 86444112 N DEL 36
SRR1766461.6828702 chr14 86443959 N chr14 86444072 N DEL 19
SRR1766464.8581884 chr14 86443425 N chr14 86444072 N DEL 11
SRR1766479.10343351 chr14 86443425 N chr14 86444072 N DEL 10
SRR1766477.314063 chr14 86443779 N chr14 86444075 N DEL 5
SRR1766452.6844358 chr14 86443884 N chr14 86444112 N DEL 23
SRR1766447.6390002 chr14 86443884 N chr14 86444112 N DEL 23
SRR1766461.3674012 chr14 86443884 N chr14 86444112 N DEL 23
SRR1766459.3077224 chr14 86443423 N chr14 86444204 N DUP 5
SRR1766460.3863870 chr14 86443523 N chr14 86444112 N DEL 17
SRR1766442.6134313 chr14 86443525 N chr14 86444114 N DEL 13
SRR1766484.12607 chr14 86443418 N chr14 86444164 N DEL 8
SRR1766447.10177067 chr14 86443419 N chr14 86444165 N DEL 7
SRR1766484.11578735 chr14 86443438 N chr14 86444221 N DEL 5
SRR1766480.749636 chr12 127166359 N chr12 127166438 N DUP 5
SRR1766464.6305303 chr12 127166359 N chr12 127166438 N DUP 5
SRR1766445.8947762 chr12 127166345 N chr12 127166404 N DUP 16
SRR1766477.9796204 chr12 127166345 N chr12 127166404 N DUP 17
SRR1766467.4660244 chr12 127166345 N chr12 127166404 N DUP 19
SRR1766461.1350871 chr12 127166359 N chr12 127166438 N DUP 35
SRR1766482.4679794 chr12 127166345 N chr12 127166404 N DUP 29
SRR1766454.8431121 chr12 127166359 N chr12 127166438 N DUP 32
SRR1766464.783149 chr12 127166359 N chr12 127166438 N DUP 33
SRR1766472.51397 chr12 127166359 N chr12 127166468 N DUP 31
SRR1766473.4510760 chr12 127166395 N chr12 127166484 N DUP 10
SRR1766446.4228944 chr12 127166395 N chr12 127166484 N DUP 10
SRR1766458.124430 chr12 127166395 N chr12 127166484 N DUP 8
SRR1766472.3442793 chr12 127166395 N chr12 127166484 N DUP 5
SRR1766456.44351 chr18 48221103 N chr18 48221306 N DEL 4
SRR1766444.1787354 chr18 48221166 N chr18 48221227 N DEL 5
SRR1766484.4873416 chr18 48221251 N chr18 48221416 N DEL 5
SRR1766480.6313399 chr18 48221288 N chr18 48221536 N DEL 15
SRR1766470.8340052 chr18 48221199 N chr18 48221422 N DUP 5
SRR1766482.8137106 chr18 48221143 N chr18 48221449 N DEL 1
SRR1766483.6051766 chr18 48221516 N chr18 48221597 N DUP 5
SRR1766457.8812702 chr18 48221386 N chr18 48221676 N DUP 5
SRR1766442.28927115 chr18 48221530 N chr18 48221676 N DUP 5
SRR1766482.617237 chr18 48221530 N chr18 48221676 N DUP 5
SRR1766444.3414975 chr18 48221530 N chr18 48221676 N DUP 5
SRR1766479.254385 chr18 48221530 N chr18 48221676 N DUP 5
SRR1766475.2634042 chr18 48221530 N chr18 48221676 N DUP 5
SRR1766467.5822698 chr18 48221227 N chr18 48222027 N DUP 4
SRR1766463.2956149 chr18 48221130 N chr18 48222031 N DUP 5
SRR1766472.2279419 chr18 48221676 N chr18 48222147 N DEL 5
SRR1766447.10807702 chr5 174522591 N chr5 174522664 N DEL 9
SRR1766482.11101854 chr5 174522637 N chr5 174522704 N DEL 12
SRR1766443.2661640 chr5 174522603 N chr5 174522705 N DEL 10
SRR1766485.5863310 chr5 174522603 N chr5 174522707 N DEL 12
SRR1766470.10496663 chr5 174522568 N chr5 174522709 N DEL 7
SRR1766449.256505 chr5 174522610 N chr5 174522712 N DEL 4
SRR1766481.13096796 chr5 174522610 N chr5 174522712 N DEL 4
SRR1766456.1197074 chr5 174522611 N chr5 174522713 N DEL 6
SRR1766479.9137295 chr5 174522608 N chr5 174522712 N DEL 7
SRR1766474.9542019 chr16 87778546 N chr16 87778597 N DEL 6
SRR1766465.6323029 chr7 157778658 N chr7 157778766 N DUP 2
SRR1766486.8348504 chr2 16143476 N chr2 16145269 N DEL 5
SRR1766461.6664474 chr2 16143486 N chr2 16145263 N DEL 5
SRR1766476.6564664 chr2 16143492 N chr2 16145265 N DEL 5
SRR1766475.137651 chr2 16143496 N chr2 16145268 N DEL 5
SRR1766442.42802242 chr2 16143498 N chr2 16145266 N DEL 5
SRR1766470.8055520 chr2 16143505 N chr2 16145263 N DEL 5
SRR1766447.8212227 chr2 16143433 N chr2 16145283 N DUP 1
SRR1766446.7166010 chr2 16143549 N chr2 16145266 N DEL 5
SRR1766469.8122257 chr2 16143518 N chr2 16145313 N DUP 5
SRR1766483.639968 chr2 16143527 N chr2 16145283 N DUP 5
SRR1766463.9347421 chr2 16143597 N chr2 16145308 N DUP 5
SRR1766482.4800626 chr2 16143597 N chr2 16145308 N DUP 5
SRR1766442.43343682 chr2 16143597 N chr2 16145305 N DUP 5
SRR1766445.2145484 chr2 16143597 N chr2 16145298 N DUP 5
SRR1766475.4721310 chr2 16143671 N chr2 16145308 N DUP 10
SRR1766484.9596680 chr2 16143743 N chr2 16145263 N DEL 8
SRR1766446.9132315 chr2 16143762 N chr2 16145266 N DEL 8
SRR1766442.25173893 chr2 16143762 N chr2 16145266 N DEL 13
SRR1766464.8631971 chr2 16143775 N chr2 16145265 N DEL 8
SRR1766483.12279119 chr2 16143958 N chr2 16145266 N DEL 5
SRR1766465.7136545 chr2 16143983 N chr2 16145267 N DEL 5
SRR1766458.3621345 chr2 16143988 N chr2 16145263 N DEL 5
SRR1766455.4632081 chr2 16144001 N chr2 16145266 N DEL 5
SRR1766461.6664474 chr2 16144061 N chr2 16145266 N DEL 4
SRR1766478.6518221 chr2 16144013 N chr2 16145309 N DUP 13
SRR1766447.11063595 chr2 16144680 N chr2 16145265 N DEL 5
SRR1766446.9680897 chr2 16144888 N chr2 16145265 N DEL 5
SRR1766442.19880547 chr17 42123845 N chr17 42124168 N DUP 13
SRR1766465.327462 chr17 42123859 N chr17 42124485 N DEL 1
SRR1766474.1787146 chr17 42123859 N chr17 42124485 N DEL 1
SRR1766444.4321571 chrX 1493542 N chrX 1493622 N DEL 4
SRR1766453.2768409 chr3 93470409 N chr3 93470458 N DUP 43
SRR1766443.7451191 chr3 93470409 N chr3 93470458 N DUP 17
SRR1766479.12580237 chr3 93470409 N chr3 93470458 N DUP 37
SRR1766463.4981021 chr3 93470409 N chr3 93470458 N DUP 16
SRR1766475.5824442 chr3 93470409 N chr3 93470458 N DUP 18
SRR1766483.573341 chr3 93470409 N chr3 93470458 N DUP 38
SRR1766478.228532 chr3 93470409 N chr3 93470458 N DUP 38
SRR1766442.33326029 chr3 93470408 N chr3 93470457 N DUP 32
SRR1766448.8458862 chr3 93470409 N chr3 93470458 N DUP 30
SRR1766449.8704930 chr3 93470409 N chr3 93470458 N DUP 27
SRR1766450.6321970 chr3 93470409 N chr3 93470458 N DUP 39
SRR1766451.501006 chr6 11427439 N chr6 11427549 N DEL 6
SRR1766457.6842969 chr6 11427490 N chr6 11427583 N DUP 4
SRR1766480.3157736 chr19 49612047 N chr19 49612354 N DEL 10
SRR1766479.2753313 chr19 49611789 N chr19 49612089 N DEL 3
SRR1766486.2721101 chr19 49611792 N chr19 49612102 N DEL 5
SRR1766478.2680648 chr19 49611803 N chr19 49612113 N DEL 5
SRR1766442.29593571 chr19 49611877 N chr19 49612187 N DEL 5
SRR1766473.3911331 chr19 49611790 N chr19 49612391 N DEL 2
SRR1766456.5198627 chr20 38590560 N chr20 38590643 N DEL 8
SRR1766462.3856335 chr10 7378207 N chr10 7378315 N DUP 5
SRR1766470.9445773 chr10 7378213 N chr10 7378333 N DUP 5
SRR1766477.4097674 chr10 7378214 N chr10 7378280 N DUP 5
SRR1766449.2002767 chr10 7378181 N chr10 7378351 N DUP 5
SRR1766442.16666031 chr10 7378306 N chr10 7378355 N DUP 15
SRR1766442.22774063 chr10 7378306 N chr10 7378355 N DUP 12
SRR1766452.1763621 chr10 7378306 N chr10 7378355 N DUP 12
SRR1766471.565636 chr3 133425952 N chr3 133426187 N DEL 2
SRR1766455.2346304 chr3 133425952 N chr3 133426187 N DEL 2
SRR1766464.1520914 chr3 133425944 N chr3 133426179 N DEL 2
SRR1766473.8656906 chr3 133425941 N chr3 133426186 N DEL 3
SRR1766458.5063665 chr2 235999560 N chr2 235999675 N DUP 6
SRR1766483.7835706 chr2 235999552 N chr2 235999747 N DUP 5
SRR1766486.1874043 chr11 119780889 N chr11 119781032 N DEL 5
SRR1766469.4338266 chr11 119780889 N chr11 119781032 N DEL 5
SRR1766478.2576777 chr11 119780916 N chr11 119781026 N DEL 7
SRR1766453.6618849 chr15 66380729 N chr15 66381351 N DEL 5
SRR1766442.18312939 chr15 66381083 N chr15 66381712 N DEL 5
SRR1766461.4273248 chr15 66381083 N chr15 66381712 N DEL 5
SRR1766481.3892807 chr15 66381223 N chr15 66381852 N DEL 5
SRR1766484.9300895 chr15 66381480 N chr15 66382108 N DEL 1
SRR1766475.1516451 chr15 66381223 N chr15 66381852 N DEL 10
SRR1766459.846978 chr15 66381302 N chr15 66381931 N DEL 5
SRR1766485.9267945 chr15 66381307 N chr15 66381936 N DEL 5
SRR1766454.8122764 chr15 66381335 N chr15 66381964 N DEL 5
SRR1766442.32608465 chr2 239421632 N chr2 239421816 N DEL 10
SRR1766442.31053216 chr2 239421632 N chr2 239421816 N DEL 14
SRR1766444.1848128 chr2 239421591 N chr2 239421775 N DEL 13
SRR1766468.3852809 chr2 239421584 N chr2 239421768 N DEL 5
SRR1766482.5968863 chr4 155813832 N chr4 155813933 N DEL 2
SRR1766445.3333163 chr4 155813832 N chr4 155813933 N DEL 2
SRR1766469.2568791 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766463.9889289 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766445.9189130 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766457.8761368 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766467.6835347 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766485.3735642 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766455.8671205 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766470.3984863 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766479.10585143 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766445.8159518 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766476.4248384 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766448.8590730 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766477.1169820 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766445.3876841 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766484.7519642 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766452.545648 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766464.6119420 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766449.4772568 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766485.11179778 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766442.46053495 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766442.9740086 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766454.6528099 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766442.40790690 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766443.10154325 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766447.1813238 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766472.10207188 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766479.554003 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766450.6992825 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766485.10017543 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766483.8393435 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766456.614727 chr4 155813851 N chr4 155813902 N DEL 5
SRR1766473.7660680 chr4 155813699 N chr4 155813902 N DEL 5
SRR1766448.2306987 chr4 155813902 N chr4 155814001 N DUP 5
SRR1766461.3733233 chr4 155813902 N chr4 155814001 N DUP 5
SRR1766462.9418726 chr4 155813902 N chr4 155813951 N DUP 5
SRR1766454.8558290 chr4 155813902 N chr4 155813951 N DUP 5
SRR1766442.1431167 chr4 155813902 N chr4 155813951 N DUP 5
SRR1766483.2573074 chr4 155813902 N chr4 155813951 N DUP 5
SRR1766464.6838706 chr4 155813902 N chr4 155813951 N DUP 5
SRR1766473.9565909 chr4 155813902 N chr4 155813951 N DUP 5
SRR1766469.6222585 chr4 155813902 N chr4 155813951 N DUP 5
SRR1766482.1430303 chr4 155813699 N chr4 155813902 N DEL 5
SRR1766483.4150044 chr4 155813699 N chr4 155813902 N DEL 5
SRR1766481.11929080 chr4 155813701 N chr4 155813904 N DEL 5
SRR1766474.6317918 chr4 155813702 N chr4 155813905 N DEL 5
SRR1766448.4888377 chr4 155813706 N chr4 155813909 N DEL 5
SRR1766463.5801853 chr4 155813706 N chr4 155813909 N DEL 5
SRR1766477.5454927 chr4 155813708 N chr4 155813911 N DEL 5
SRR1766484.2558054 chr4 155813712 N chr4 155813915 N DEL 2
SRR1766445.3985009 chr4 155813713 N chr4 155813916 N DEL 1
SRR1766457.2240574 chr4 155813872 N chr4 155814047 N DUP 5
SRR1766446.2936681 chr4 155813872 N chr4 155814047 N DUP 5
SRR1766485.7572117 chr4 155813837 N chr4 155813964 N DEL 5
SRR1766453.3408308 chr4 155813675 N chr4 155813996 N DEL 2
SRR1766445.5324104 chr4 155813870 N chr4 155814047 N DEL 5
SRR1766481.7109412 chr4 155813769 N chr4 155813894 N DUP 5
SRR1766481.10553537 chr4 155813769 N chr4 155813894 N DUP 5
SRR1766449.7926828 chr4 155813769 N chr4 155813894 N DUP 5
SRR1766465.3186621 chr4 155813677 N chr4 155814074 N DEL 5
SRR1766474.11590493 chr4 155813832 N chr4 155813933 N DEL 4
SRR1766459.7497948 chr4 155813832 N chr4 155813933 N DEL 5
SRR1766468.910099 chr4 155813680 N chr4 155814077 N DEL 5
SRR1766467.8739756 chr4 155813734 N chr4 155814087 N DEL 4
SRR1766460.6510719 chr4 155813708 N chr4 155814087 N DEL 5
SRR1766475.11020464 chr4 155813894 N chr4 155814121 N DEL 5
SRR1766484.4912473 chr11 86862629 N chr11 86862741 N DUP 5
SRR1766453.8571909 chr11 86862818 N chr11 86863005 N DUP 6
SRR1766457.7857541 chr11 86862818 N chr11 86863005 N DUP 6
SRR1766485.1478883 chr11 86862818 N chr11 86863005 N DUP 6
SRR1766466.6829072 chr11 86862818 N chr11 86863005 N DUP 6
SRR1766465.8957514 chr2 239643044 N chr2 239643174 N DUP 5
SRR1766480.4569413 chr3 126978544 N chr3 126978655 N DUP 5
SRR1766446.547259 chr3 35748095 N chr3 35748324 N DEL 3
SRR1766459.10437719 chr3 35748095 N chr3 35748324 N DEL 5
SRR1766484.8535530 chr3 35748095 N chr3 35748324 N DEL 5
SRR1766446.4939025 chr3 35748095 N chr3 35748324 N DEL 5
SRR1766460.3406860 chr3 35748213 N chr3 35748434 N DEL 13
SRR1766451.1405939 chr3 35748259 N chr3 35748471 N DEL 9
SRR1766454.226758 chr3 35748372 N chr3 35748434 N DEL 2
SRR1766465.3682713 chr3 35748113 N chr3 35748280 N DEL 9
SRR1766462.5665021 chr3 35748113 N chr3 35748280 N DEL 10
SRR1766481.11643755 chr3 35748211 N chr3 35748440 N DEL 5
SRR1766442.6201418 chr3 35748432 N chr3 35748636 N DUP 10
SRR1766447.9867953 chr12 34301397 N chr12 34302239 N DEL 5
SRR1766465.1614826 chr12 34301593 N chr12 34301803 N DEL 3
SRR1766481.1776621 chr12 34301279 N chr12 34301699 N DUP 5
SRR1766486.1735191 chr12 34301311 N chr12 34301733 N DEL 15
SRR1766445.8880094 chr12 34301305 N chr12 34301727 N DEL 10
SRR1766485.9240589 chr12 34301349 N chr12 34302190 N DEL 12
SRR1766478.6052757 chr12 34301422 N chr12 34302475 N DEL 15
SRR1766460.1158988 chr7 67997661 N chr7 67997749 N DEL 5
SRR1766471.1733227 chr7 67997665 N chr7 67997749 N DEL 1
SRR1766443.3760953 chr7 67997665 N chr7 67997749 N DEL 2
SRR1766456.2063660 chr7 67997739 N chr7 67997811 N DEL 7
SRR1766477.895066 chr2 33911356 N chr2 33911419 N DEL 12
SRR1766486.7826877 chr11 2048095 N chr11 2048220 N DUP 5
SRR1766482.10136339 chr11 1628484 N chr11 1628549 N DUP 5
SRR1766443.9991109 chr11 1628484 N chr11 1628549 N DUP 5
SRR1766482.8865151 chr11 1628507 N chr11 1628574 N DEL 5
SRR1766461.7677152 chr11 1628535 N chr11 1628602 N DEL 5
SRR1766486.1635450 chr11 1628543 N chr11 1628610 N DEL 4
SRR1766462.3631852 chr1 220012868 N chr1 220012974 N DEL 9
SRR1766457.4849288 chr1 220012852 N chr1 220012956 N DUP 2
SRR1766480.8159475 chr1 220012938 N chr1 220013042 N DUP 16
SRR1766478.4506607 chr1 220012938 N chr1 220013042 N DUP 13
SRR1766457.8397286 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766450.7496326 chr1 220012938 N chr1 220013042 N DUP 14
SRR1766484.5501658 chr1 220012938 N chr1 220013042 N DUP 14
SRR1766461.2699270 chr1 220012938 N chr1 220013042 N DUP 11
SRR1766472.11486622 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766447.7842760 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766474.8348644 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766442.29118002 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766482.4618864 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766442.37559474 chr1 220012938 N chr1 220013042 N DUP 10
SRR1766464.1769644 chr1 220012916 N chr1 220013020 N DUP 5
SRR1766476.10057346 chr1 220012938 N chr1 220013042 N DUP 6
SRR1766472.232286 chr1 220012938 N chr1 220013042 N DUP 5
SRR1766467.8910960 chr1 220012938 N chr1 220013042 N DUP 5
SRR1766449.9105801 chr1 220012938 N chr1 220013042 N DUP 5
SRR1766446.9949506 chr1 220012938 N chr1 220013042 N DUP 5
SRR1766478.5541851 chr1 220012938 N chr1 220013042 N DUP 1
SRR1766451.4489784 chr1 220012938 N chr1 220013042 N DUP 5
SRR1766479.9545280 chr1 220012938 N chr1 220013042 N DUP 3
SRR1766459.741739 chr1 220012938 N chr1 220013042 N DUP 5
SRR1766450.3828786 chr1 220012938 N chr1 220013042 N DUP 5
SRR1766478.3735431 chr1 220012938 N chr1 220013042 N DUP 7
SRR1766454.5941028 chr1 220012938 N chr1 220013042 N DUP 5
SRR1766486.5171321 chr1 220012938 N chr1 220013042 N DUP 9
SRR1766447.1280491 chr1 220012938 N chr1 220013042 N DUP 11
SRR1766449.8955448 chr1 220012940 N chr1 220013044 N DUP 3
SRR1766466.5201590 chr1 220012938 N chr1 220013042 N DUP 11
SRR1766442.45625176 chr1 220012882 N chr1 220012988 N DEL 1
SRR1766485.7704134 chr1 11135798 N chr1 11136100 N DEL 14
SRR1766447.3532645 chr1 11135739 N chr1 11136041 N DEL 5
SRR1766485.4161943 chr1 11135790 N chr1 11136092 N DEL 5
SRR1766450.2134984 chr1 11135803 N chr1 11136105 N DEL 5
SRR1766469.8596490 chr7 138174569 N chr7 138174662 N DEL 13
SRR1766474.9648697 chr7 138174569 N chr7 138174662 N DEL 13
SRR1766442.23752160 chr7 138174569 N chr7 138174662 N DEL 13
SRR1766442.39213418 chr7 138174495 N chr7 138174669 N DEL 8
SRR1766473.3426607 chr7 138174498 N chr7 138174672 N DEL 5
SRR1766461.10141188 chr6 23802194 N chr6 23802291 N DEL 7
SRR1766472.8479695 chr6 23802191 N chr6 23802302 N DEL 12
SRR1766484.7172295 chr6 23802192 N chr6 23802303 N DEL 11
SRR1766477.8114459 chr6 23802234 N chr6 23802313 N DEL 1
SRR1766452.6476435 chr6 23802195 N chr6 23802306 N DEL 8
SRR1766465.4204474 chr6 23802194 N chr6 23802305 N DEL 9
SRR1766474.8638837 chr12 116652096 N chr12 116652175 N DUP 3
SRR1766445.1875357 chr12 116652096 N chr12 116652199 N DUP 13
SRR1766480.3500644 chr12 116652096 N chr12 116652199 N DUP 13
SRR1766476.2952469 chr12 116652002 N chr12 116652198 N DUP 12
SRR1766469.8966842 chr12 116652032 N chr12 116652178 N DEL 12
SRR1766470.878799 chr12 116652025 N chr12 116652175 N DEL 15
SRR1766462.7735033 chr12 116652114 N chr12 116652175 N DEL 17
SRR1766465.326487 chr12 116652110 N chr12 116652175 N DEL 15
SRR1766442.39744083 chr12 116652111 N chr12 116652184 N DEL 6
SRR1766442.1833073 chr12 116652025 N chr12 116652195 N DEL 4
SRR1766482.8648329 chr12 116652025 N chr12 116652195 N DEL 4
SRR1766478.2955197 chr12 116652110 N chr12 116652179 N DEL 11
SRR1766483.816841 chr12 116652016 N chr12 116652202 N DEL 4
SRR1766479.2916449 chr4 163894706 N chr4 163894774 N DUP 27
SRR1766482.8152960 chr4 163894706 N chr4 163894774 N DUP 27
SRR1766447.11446666 chr4 163894706 N chr4 163894774 N DUP 28
SRR1766471.5449216 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766478.1121405 chr4 163894706 N chr4 163894774 N DUP 34
SRR1766442.13216659 chr4 163894706 N chr4 163894774 N DUP 28
SRR1766442.23537322 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766459.9368097 chr4 163894706 N chr4 163894774 N DUP 34
SRR1766460.10824500 chr4 163894706 N chr4 163894774 N DUP 31
SRR1766467.6722339 chr4 163894706 N chr4 163894774 N DUP 30
SRR1766471.1311902 chr4 163894706 N chr4 163894774 N DUP 34
SRR1766471.6440397 chr4 163894706 N chr4 163894774 N DUP 33
SRR1766472.9948279 chr4 163894706 N chr4 163894774 N DUP 31
SRR1766478.767736 chr4 163894706 N chr4 163894774 N DUP 18
SRR1766479.8815481 chr4 163894706 N chr4 163894774 N DUP 34
SRR1766442.10322986 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766442.12261298 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766443.6385912 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766449.6458596 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766472.2736243 chr4 163894706 N chr4 163894774 N DUP 26
SRR1766449.6186756 chr4 163894706 N chr4 163894774 N DUP 27
SRR1766483.4538915 chr4 163894780 N chr4 163894840 N DEL 18
SRR1766486.11865358 chr4 163894780 N chr4 163894840 N DEL 18
SRR1766446.3686635 chr4 163894706 N chr4 163894774 N DUP 27
SRR1766447.771987 chr4 163894706 N chr4 163894774 N DUP 28
SRR1766446.2422617 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766471.1652729 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766477.9359985 chr4 163894706 N chr4 163894774 N DUP 30
SRR1766469.4720168 chr4 163894706 N chr4 163894774 N DUP 32
SRR1766469.6241735 chr4 163894706 N chr4 163894774 N DUP 32
SRR1766466.9190665 chr4 163894780 N chr4 163894840 N DEL 22
SRR1766457.4566415 chr4 163894706 N chr4 163894774 N DUP 29
SRR1766466.5281676 chr4 163894706 N chr4 163894774 N DUP 19
SRR1766479.8449256 chr4 163894706 N chr4 163894774 N DUP 19
SRR1766444.2914134 chr4 163894706 N chr4 163894774 N DUP 19
SRR1766468.5657479 chr4 163894780 N chr4 163894840 N DEL 27
SRR1766470.5628948 chr4 163894757 N chr4 163894840 N DEL 25
SRR1766463.1287744 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766464.10859506 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766469.5846318 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766455.3996277 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766442.2394403 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766469.5548198 chr4 163894757 N chr4 163894840 N DEL 22
SRR1766448.2239811 chr4 163894821 N chr4 163894904 N DUP 11
SRR1766480.4696999 chr4 163894786 N chr4 163894913 N DEL 8
SRR1766451.6251880 chr4 163894734 N chr4 163894840 N DEL 12
SRR1766485.2556431 chr4 163894734 N chr4 163894840 N DEL 9
SRR1766443.2916224 chr4 163894734 N chr4 163894840 N DEL 9
SRR1766463.8626599 chr4 163894713 N chr4 163894779 N DUP 16
SRR1766478.647037 chr4 163894738 N chr4 163894844 N DEL 9
SRR1766467.3053664 chr1 7995124 N chr1 7995236 N DUP 7
SRR1766468.704813 chr1 7995168 N chr1 7995240 N DUP 7
SRR1766453.6990199 chrX 57698243 N chrX 57698806 N DUP 15
SRR1766479.13431829 chrX 57697226 N chrX 57698256 N DEL 5
SRR1766478.4776782 chrX 57698325 N chrX 57698393 N DUP 9
SRR1766479.1250646 chrX 57698279 N chrX 57698704 N DEL 15
SRR1766447.11392507 chrX 57698303 N chrX 57698402 N DUP 17
SRR1766484.11020182 chrX 57698188 N chrX 57698702 N DUP 27
SRR1766472.11492922 chrX 57698191 N chrX 57698743 N DUP 19
SRR1766463.1756856 chrX 57698191 N chrX 57698743 N DUP 22
SRR1766480.8317691 chrX 57697517 N chrX 57698793 N DUP 16
SRR1766447.8639660 chrX 57698637 N chrX 57698711 N DUP 19
SRR1766455.3622714 chrX 57698385 N chrX 57698792 N DEL 11
SRR1766486.6530118 chrX 57698119 N chrX 57698711 N DEL 4
SRR1766464.6462547 chrX 57698325 N chrX 57698800 N DEL 15
SRR1766442.22382523 chrX 57698352 N chrX 57698793 N DEL 20
SRR1766485.4068355 chrX 57698336 N chrX 57698811 N DEL 9
SRR1766478.3119570 chr12 163288 N chr12 163350 N DEL 5
SRR1766452.7226477 chr12 163315 N chr12 163377 N DEL 5
SRR1766443.9148985 chr12 163361 N chr12 163520 N DUP 10
SRR1766444.7175308 chr12 163340 N chr12 163466 N DEL 3
SRR1766466.1062286 chr5 28597068 N chr5 28597165 N DUP 1
SRR1766483.3278211 chr5 28597094 N chr5 28597191 N DUP 5
SRR1766463.1360890 chr8 675298 N chr8 676149 N DEL 10
SRR1766442.23902793 chr8 675326 N chr8 676149 N DEL 4
SRR1766474.1508809 chr8 675377 N chr8 675871 N DUP 5
SRR1766470.10942897 chr8 675417 N chr8 676376 N DUP 5
SRR1766442.8484288 chr8 675381 N chr8 675490 N DUP 5
SRR1766459.2913150 chr8 675510 N chr8 676114 N DEL 5
SRR1766448.3331198 chr8 675381 N chr8 675545 N DUP 10
SRR1766452.6322525 chr8 675601 N chr8 676149 N DEL 8
SRR1766460.10552506 chr8 675326 N chr8 675546 N DEL 5
SRR1766442.32735876 chr8 675614 N chr8 676327 N DEL 1
SRR1766478.10319764 chr8 676022 N chr8 676600 N DEL 5
SRR1766450.2990230 chr8 675558 N chr8 676160 N DUP 5
SRR1766479.2164438 chr8 675397 N chr8 676136 N DUP 4
SRR1766486.7242873 chr8 675738 N chr8 676149 N DEL 5
SRR1766460.1098885 chr8 675381 N chr8 675545 N DUP 10
SRR1766453.1051698 chr8 675455 N chr8 676005 N DEL 1
SRR1766486.3205071 chr8 675279 N chr8 675524 N DUP 5
SRR1766471.265141 chr8 675875 N chr8 676149 N DEL 4
SRR1766443.4606196 chr8 675300 N chr8 676121 N DUP 5
SRR1766452.10317402 chr8 675867 N chr8 676060 N DEL 3
SRR1766466.1598569 chr8 675408 N chr8 675958 N DEL 5
SRR1766467.2112010 chr8 675299 N chr8 675958 N DEL 5
SRR1766486.7242873 chr8 675299 N chr8 675958 N DEL 5
SRR1766475.2074777 chr8 676020 N chr8 676598 N DEL 5
SRR1766466.833611 chr8 675950 N chr8 676113 N DUP 5
SRR1766452.9745485 chr8 675390 N chr8 675968 N DEL 5
SRR1766467.3787632 chr8 675902 N chr8 676040 N DEL 5
SRR1766459.10100389 chr8 675272 N chr8 676148 N DUP 5
SRR1766472.9457855 chr8 676177 N chr8 676312 N DUP 10
SRR1766442.17080050 chr8 675287 N chr8 676165 N DEL 4
SRR1766471.265141 chr8 676153 N chr8 676209 N DEL 10
SRR1766462.6195157 chr8 675877 N chr8 676206 N DEL 5
SRR1766467.8091979 chr8 675867 N chr8 676277 N DEL 5
SRR1766469.10085650 chr8 676153 N chr8 676290 N DEL 5
SRR1766480.6037195 chr8 675994 N chr8 676377 N DUP 5
SRR1766448.5518291 chr8 675994 N chr8 676377 N DUP 17
SRR1766479.6653007 chr8 675814 N chr8 676388 N DUP 10
SRR1766481.9376279 chr8 675873 N chr8 676339 N DEL 4
SRR1766448.10430876 chr8 675511 N chr8 676388 N DUP 13
SRR1766460.8211552 chr8 675511 N chr8 676388 N DUP 10
SRR1766476.703548 chr8 675873 N chr8 676422 N DEL 4
SRR1766471.10235038 chr8 676113 N chr8 676443 N DEL 8
SRR1766459.1254797 chr8 675620 N chr8 676114 N DEL 1
SRR1766477.3212384 chr8 675994 N chr8 676377 N DUP 17
SRR1766475.8708604 chr8 675872 N chr8 676476 N DEL 5
SRR1766454.2962923 chr8 675511 N chr8 676388 N DUP 12
SRR1766473.1928273 chr8 675876 N chr8 676480 N DEL 3
SRR1766451.5430175 chr8 675878 N chr8 676372 N DEL 4
SRR1766447.6296919 chr8 675867 N chr8 676637 N DEL 16
SRR1766442.36034255 chr7 2064807 N chr7 2065097 N DEL 6
SRR1766442.47010134 chr11 36202760 N chr11 36202812 N DUP 4
SRR1766449.6896906 chr11 36202760 N chr11 36202812 N DUP 5
SRR1766473.8452067 chr11 36202787 N chr11 36202841 N DEL 5
SRR1766443.3654201 chr11 36202787 N chr11 36202841 N DEL 5
SRR1766445.303264 chr11 36202787 N chr11 36202841 N DEL 5
SRR1766450.3218911 chr11 36202787 N chr11 36202841 N DEL 5
SRR1766460.1773016 chr11 36202787 N chr11 36202841 N DEL 5
SRR1766455.6657410 chr11 36202787 N chr11 36202841 N DEL 5
SRR1766456.3561354 chr11 36202787 N chr11 36202841 N DEL 5
SRR1766442.26630603 chr11 36202796 N chr11 36202850 N DEL 5
SRR1766461.7657361 chr20 61273107 N chr20 61273207 N DEL 5
SRR1766475.6201455 chr20 61272961 N chr20 61273235 N DUP 5
SRR1766466.7177960 chr15 82145145 N chr15 82145453 N DEL 9
SRR1766445.8177008 chr15 82145155 N chr15 82145466 N DUP 5
SRR1766486.5456397 chr16 22780342 N chr16 22780407 N DUP 2
SRR1766450.370449 chr16 22780295 N chr16 22780356 N DEL 1
SRR1766482.8277393 chr16 22780277 N chr16 22780404 N DEL 5
SRR1766466.9065571 chr16 22780312 N chr16 22780403 N DUP 9
SRR1766445.8520500 chr16 22780435 N chr16 22780564 N DUP 5
SRR1766468.5079575 chr16 22780434 N chr16 22780535 N DEL 9
SRR1766454.8905690 chr1 118319453 N chr1 118319548 N DUP 9
SRR1766454.4311037 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766442.23620487 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766444.1123921 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766461.3364703 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766474.11180459 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766474.4132836 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766477.5017017 chr1 118319485 N chr1 118319548 N DUP 15
SRR1766477.7916256 chr1 118319485 N chr1 118319548 N DUP 14
SRR1766454.5169580 chr1 118319452 N chr1 118319517 N DEL 5
SRR1766445.3090625 chr1 118319452 N chr1 118319517 N DEL 5
SRR1766460.4944063 chr1 118319452 N chr1 118319517 N DEL 5
SRR1766445.7842667 chr1 118319452 N chr1 118319517 N DEL 5
SRR1766442.3553134 chr1 118319460 N chr1 118319525 N DEL 5
SRR1766442.23755822 chr1 118319426 N chr1 118319523 N DEL 5
SRR1766466.9344091 chr1 118319431 N chr1 118319528 N DEL 4
SRR1766459.10495101 chr1 118319432 N chr1 118319529 N DEL 3
SRR1766479.10959502 chr1 118319593 N chr1 118319666 N DUP 1
SRR1766481.2045869 chr10 78613561 N chr10 78613730 N DUP 7
SRR1766474.7770053 chr2 131754152 N chr2 131754756 N DEL 8
SRR1766472.91195 chr2 131754162 N chr2 131754766 N DEL 5
SRR1766467.319842 chr2 131754091 N chr2 131754497 N DUP 5
SRR1766445.3799577 chr2 131754264 N chr2 131754869 N DEL 2
SRR1766485.982640 chr2 131754195 N chr2 131754385 N DUP 5
SRR1766445.4033811 chr2 131754323 N chr2 131754938 N DEL 5
SRR1766456.549129 chr2 131754323 N chr2 131754938 N DEL 5
SRR1766451.1865373 chr2 131754385 N chr2 131754798 N DEL 5
SRR1766467.3889060 chr2 131754385 N chr2 131754798 N DEL 5
SRR1766460.10224969 chr2 131754339 N chr2 131754952 N DUP 5
SRR1766471.7307468 chr2 131754341 N chr2 131754954 N DUP 3
SRR1766442.40045430 chr2 131754522 N chr2 131754918 N DEL 10
SRR1766448.3290773 chr2 131754542 N chr2 131755157 N DEL 1
SRR1766474.640842 chr2 131754646 N chr2 131755480 N DEL 15
SRR1766469.8960643 chr2 131754783 N chr2 131754986 N DEL 4
SRR1766449.2898239 chr2 131754937 N chr2 131755157 N DEL 5
SRR1766458.1347509 chr2 131754989 N chr2 131755209 N DEL 5
SRR1766448.5357778 chr2 131754971 N chr2 131755408 N DUP 5
SRR1766448.8849974 chr2 131755218 N chr2 131755438 N DEL 10
SRR1766442.6428061 chr2 131755223 N chr2 131755443 N DEL 5
SRR1766476.4843880 chr2 131755155 N chr2 131755375 N DEL 5
SRR1766463.147334 chr2 131754929 N chr2 131755149 N DEL 3
SRR1766448.3290773 chr2 131755189 N chr2 131755407 N DUP 5
SRR1766481.1627521 chr2 131753912 N chr2 131755349 N DUP 5
SRR1766486.956846 chr2 131755125 N chr2 131755343 N DUP 5
SRR1766471.5055056 chr2 131754091 N chr2 131755332 N DEL 14
SRR1766464.4352896 chr2 131754110 N chr2 131755354 N DEL 5
SRR1766446.2186628 chr2 131754023 N chr2 131755460 N DUP 2
SRR1766477.8390449 chr2 131754122 N chr2 131755366 N DEL 3
SRR1766442.8905190 chr2 131755410 N chr2 131755610 N DEL 5
SRR1766485.3276432 chr2 131755155 N chr2 131755375 N DEL 5
SRR1766462.8268510 chr2 131754562 N chr2 131755396 N DEL 10
SRR1766451.1949286 chr2 131754236 N chr2 131755480 N DUP 10
SRR1766445.8343522 chr2 131754041 N chr2 131755478 N DUP 20
SRR1766485.8599802 chr2 131755382 N chr2 131755582 N DEL 5
SRR1766458.7167720 chr2 131755382 N chr2 131755582 N DEL 5
SRR1766478.8628814 chr2 131754236 N chr2 131755679 N DUP 10
SRR1766452.10126581 chr2 131754561 N chr2 131755594 N DEL 3
SRR1766459.7886197 chr2 131755414 N chr2 131755614 N DEL 5
SRR1766453.4431327 chr2 131755366 N chr2 131755763 N DUP 5
SRR1766442.6002011 chr2 131755366 N chr2 131755763 N DUP 5
SRR1766445.4447575 chr2 131755366 N chr2 131755763 N DUP 5
SRR1766442.34828794 chr2 131755366 N chr2 131755763 N DUP 5
SRR1766464.6902198 chr20 48125024 N chr20 48125219 N DUP 5
SRR1766471.6202922 chr20 48125131 N chr20 48125415 N DEL 7
SRR1766442.35100020 chr20 48125032 N chr20 48125129 N DUP 7
SRR1766486.4764552 chr20 48125179 N chr20 48125463 N DEL 5
SRR1766442.21346585 chr20 48125179 N chr20 48125512 N DEL 5
SRR1766442.2446579 chr20 48125286 N chr20 48125383 N DUP 5
SRR1766483.3334794 chr20 48125041 N chr20 48125421 N DUP 5
SRR1766446.6741695 chr20 48125067 N chr20 48125351 N DEL 5
SRR1766483.2413574 chr20 48124971 N chr20 48125353 N DEL 5
SRR1766461.5217730 chr20 48125078 N chr20 48125362 N DEL 4
SRR1766446.5098337 chr20 48125013 N chr20 48125444 N DEL 4
SRR1766466.969770 chr17 8136052 N chr17 8136369 N DEL 5
SRR1766471.4998412 chr17 8136303 N chr17 8136618 N DUP 7
SRR1766450.4967247 chr17 8136303 N chr17 8136618 N DUP 7
SRR1766446.7113318 chr17 8136318 N chr17 8136635 N DEL 4
SRR1766483.8186047 chr17 8136318 N chr17 8136635 N DEL 4
SRR1766477.3335348 chr3 74984935 N chr3 74985096 N DEL 2
SRR1766484.1666974 chr3 74984935 N chr3 74985096 N DEL 2
SRR1766478.7593019 chr3 74984935 N chr3 74985096 N DEL 5
SRR1766459.8330245 chr3 74984935 N chr3 74985096 N DEL 5
SRR1766463.2670227 chr3 74984935 N chr3 74985096 N DEL 5
SRR1766485.11001027 chr3 74984935 N chr3 74985096 N DEL 5
SRR1766455.450447 chr3 74984952 N chr3 74985111 N DUP 5
SRR1766446.6536535 chr3 74984955 N chr3 74985114 N DUP 5
SRR1766482.8675257 chr3 74984956 N chr3 74985115 N DUP 5
SRR1766474.4846519 chr3 74984835 N chr3 74984964 N DEL 3
SRR1766467.7509102 chr3 74984966 N chr3 74985125 N DUP 1
SRR1766455.1617730 chr9 15642456 N chr9 15642507 N DUP 8
SRR1766457.563056 chr15 43580209 N chr15 43580346 N DEL 5
SRR1766449.10570729 chr8 128826802 N chr8 128827192 N DEL 5
SRR1766463.5331220 chr8 128826944 N chr8 128827019 N DUP 2
SRR1766459.2752207 chr8 128826797 N chr8 128827029 N DUP 5
SRR1766443.3967830 chr8 128826733 N chr8 128826982 N DEL 5
SRR1766443.8443962 chr8 128826926 N chr8 128827043 N DEL 5
SRR1766477.9897683 chr8 128826926 N chr8 128827043 N DEL 5
SRR1766442.32917741 chr8 128826813 N chr8 128827047 N DEL 4
SRR1766463.4408250 chr8 128826827 N chr8 128827217 N DEL 5
SRR1766477.7371702 chrY 10924331 N chrY 10924451 N DEL 8
SRR1766442.22223650 chrY 10924464 N chrY 10924553 N DUP 3
SRR1766467.7350027 chrY 10924559 N chrY 10924655 N DEL 2
SRR1766463.3710887 chrY 10924556 N chrY 10924652 N DEL 4
SRR1766479.6922269 chrY 10924556 N chrY 10924652 N DEL 5
SRR1766465.9780291 chrY 10924530 N chrY 10924666 N DEL 1
SRR1766442.438630 chrY 10924454 N chrY 10924538 N DUP 15
SRR1766473.11652537 chrY 10924492 N chrY 10924561 N DUP 9
SRR1766465.1310039 chrY 10924331 N chrY 10924466 N DEL 8
SRR1766464.1692850 chr22 43968417 N chr22 43968494 N DEL 8
SRR1766474.11222621 chr7 121088825 N chr7 121088942 N DUP 10
SRR1766479.9813574 chr9 129396731 N chr9 129396812 N DUP 5
SRR1766469.4071272 chr9 129396686 N chr9 129396899 N DUP 1
SRR1766442.35404240 chr4 3809314 N chr4 3809470 N DEL 12
SRR1766446.9714077 chr12 122973635 N chr12 122974117 N DEL 5
SRR1766464.9355145 chr12 122973576 N chr12 122973872 N DUP 5
SRR1766473.7969064 chr12 122973617 N chr12 122973915 N DEL 5
SRR1766466.3101809 chr12 122973465 N chr12 122973897 N DEL 5
SRR1766475.7743812 chr5 126784783 N chr5 126785415 N DEL 3
SRR1766443.2562577 chr5 126784809 N chr5 126785296 N DEL 2
SRR1766476.10384434 chr5 126784810 N chr5 126785630 N DEL 3
SRR1766486.1060408 chr5 126785223 N chr5 126785536 N DEL 1
SRR1766454.1002181 chr5 126785223 N chr5 126785536 N DEL 3
SRR1766452.5134650 chr5 126784923 N chr5 126785242 N DUP 6
SRR1766462.5594347 chr5 126785259 N chr5 126785572 N DEL 5
SRR1766473.9017380 chr5 126784820 N chr5 126785308 N DEL 3
SRR1766466.5930966 chr5 126784809 N chr5 126785444 N DUP 2
SRR1766445.353407 chr5 126785047 N chr5 126785372 N DEL 2
SRR1766476.7503955 chr1 218598632 N chr1 218598697 N DEL 5
SRR1766485.4772946 chr1 218598632 N chr1 218598697 N DEL 1
SRR1766474.775322 chr1 218598648 N chr1 218598711 N DUP 5
SRR1766442.30614974 chr1 218598825 N chr1 218598885 N DUP 5
SRR1766478.6250438 chr1 218598851 N chr1 218598911 N DUP 5
SRR1766465.10575103 chr16 90032570 N chr16 90032783 N DUP 5
SRR1766442.27773815 chr16 90032609 N chr16 90032719 N DEL 5
SRR1766447.4960551 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766451.1294356 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766480.6458147 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766448.7728452 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766476.10535936 chr3 84516437 N chr3 84516514 N DUP 5
SRR1766452.6457632 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766471.3981639 chr3 84516467 N chr3 84516544 N DUP 3
SRR1766445.10605601 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766479.3685808 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766464.2035149 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766481.122743 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766457.108051 chr3 84516444 N chr3 84516521 N DUP 5
SRR1766472.6183303 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766475.572756 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766442.21755581 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766454.6473201 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766455.9327672 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766443.7549029 chr3 84516444 N chr3 84516521 N DUP 5
SRR1766454.5017318 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766461.6654990 chr3 84516444 N chr3 84516521 N DUP 5
SRR1766460.4567726 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766477.723875 chr3 84516485 N chr3 84516564 N DEL 5
SRR1766470.9807630 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766453.1298845 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766443.5375404 chr3 84516491 N chr3 84516570 N DEL 5
SRR1766442.43446912 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766473.7594092 chr3 84516492 N chr3 84516571 N DEL 5
SRR1766467.10601920 chr3 84516492 N chr3 84516571 N DEL 5
SRR1766442.8079287 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766472.10160332 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766486.9040062 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766445.10675589 chr3 84516467 N chr3 84516544 N DUP 2
SRR1766460.3868142 chr3 84516508 N chr3 84516585 N DUP 5
SRR1766442.9048901 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766479.7344356 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766466.842296 chr3 84516514 N chr3 84516591 N DUP 2
SRR1766472.8888319 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766443.10394862 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766467.5469839 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766477.3393790 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766479.10083035 chr3 84516483 N chr3 84516560 N DUP 5
SRR1766442.46584708 chr3 84516454 N chr3 84516533 N DEL 4
SRR1766472.4524976 chr3 84516508 N chr3 84516585 N DUP 5
SRR1766465.726860 chr3 84516462 N chr3 84516695 N DUP 9
SRR1766451.10128570 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766449.8101899 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766473.5415678 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766452.5404735 chr3 84516482 N chr3 84516561 N DEL 5
SRR1766447.1095830 chr3 84516483 N chr3 84516562 N DEL 5
SRR1766454.5465673 chr3 84516486 N chr3 84516565 N DEL 5
SRR1766463.9162347 chr3 84516486 N chr3 84516565 N DEL 5
SRR1766449.1976117 chr3 84516451 N chr3 84516530 N DEL 5
SRR1766479.9674692 chr3 84516495 N chr3 84516574 N DEL 2
SRR1766475.6461909 chr3 84516504 N chr3 84516581 N DUP 1
SRR1766471.8139402 chr3 84516452 N chr3 84516702 N DUP 3
SRR1766481.6074095 chr3 84516452 N chr3 84516702 N DUP 4
SRR1766442.39109873 chr3 84516462 N chr3 84516695 N DUP 6
SRR1766466.6673304 chr3 84516482 N chr3 84516600 N DEL 5
SRR1766442.20777926 chr3 84516483 N chr3 84516601 N DEL 5
SRR1766482.3427920 chr3 84516490 N chr3 84516608 N DEL 5
SRR1766466.8611578 chr3 84516559 N chr3 84516737 N DUP 12
SRR1766467.2451381 chr3 84516559 N chr3 84516737 N DUP 12
SRR1766484.399139 chr3 84516559 N chr3 84516737 N DUP 12
SRR1766443.8950394 chr3 84516559 N chr3 84516737 N DUP 12
SRR1766458.4877101 chr3 84516629 N chr3 84516710 N DEL 7
SRR1766482.4537973 chr3 84516629 N chr3 84516710 N DEL 7
SRR1766447.9136130 chr3 84516629 N chr3 84516710 N DEL 7
SRR1766448.5861303 chr3 84516629 N chr3 84516710 N DEL 7
SRR1766462.10869914 chr3 84516629 N chr3 84516710 N DEL 7
SRR1766451.2327053 chr3 84516629 N chr3 84516710 N DEL 7
SRR1766484.2673446 chr3 84516590 N chr3 84516710 N DEL 7
SRR1766483.9073100 chr3 84516590 N chr3 84516710 N DEL 7
SRR1766478.7061796 chr3 84516729 N chr3 84516792 N DUP 16
SRR1766480.5945635 chr13 96400390 N chr13 96400441 N DUP 4
SRR1766448.571802 chr9 127746786 N chr9 127746922 N DEL 4
SRR1766462.6307534 chr10 126938917 N chr10 126938982 N DEL 5
SRR1766470.3809338 chr10 126938917 N chr10 126938982 N DEL 7
SRR1766469.8070109 chr10 126938917 N chr10 126938982 N DEL 8
SRR1766479.10019109 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766473.706836 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766485.912074 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766452.5053281 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766465.2700061 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766471.10810924 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766453.4648880 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766480.6438425 chr10 126938917 N chr10 126938982 N DEL 10
SRR1766464.1722466 chr10 126938916 N chr10 126939285 N DEL 5
SRR1766442.7414230 chr1 16284751 N chr1 16284886 N DUP 5
SRR1766452.59891 chr1 16284751 N chr1 16284886 N DUP 5
SRR1766462.10289388 chr1 16284751 N chr1 16284886 N DUP 5
SRR1766462.9410321 chr1 16284751 N chr1 16284886 N DUP 5
SRR1766462.11068409 chr1 16284751 N chr1 16284886 N DUP 5
SRR1766475.10565809 chr17 77920613 N chr17 77920751 N DEL 5
SRR1766485.2059701 chr17 77920548 N chr17 77920681 N DUP 15
SRR1766461.803893 chr9 128439918 N chr9 128440214 N DEL 20
SRR1766450.3464670 chrX 78175574 N chrX 78175633 N DUP 5
SRR1766484.3812985 chrX 78175514 N chrX 78175625 N DEL 4
SRR1766464.8179054 chr10 445379 N chr10 445507 N DEL 1
SRR1766471.3108876 chr10 445410 N chr10 445625 N DEL 5
SRR1766469.4920453 chr10 445325 N chr10 445451 N DUP 2
SRR1766442.24729068 chr10 445506 N chr10 445892 N DEL 1
SRR1766452.2415506 chr10 445340 N chr10 445552 N DUP 5
SRR1766447.10087363 chr10 445590 N chr10 445677 N DEL 5
SRR1766450.4982186 chr10 445399 N chr10 445612 N DUP 6
SRR1766475.1850424 chr10 445445 N chr10 445616 N DUP 4
SRR1766486.5963052 chr10 445325 N chr10 445623 N DUP 5
SRR1766444.3552471 chr10 445462 N chr10 445677 N DEL 4
SRR1766474.11730663 chr10 445363 N chr10 445789 N DUP 5
SRR1766451.7553624 chr10 445702 N chr10 445871 N DUP 4
SRR1766463.415130 chr10 445746 N chr10 446513 N DUP 6
SRR1766484.7854327 chr10 445337 N chr10 445849 N DEL 2
SRR1766479.1672678 chr10 445318 N chr10 446000 N DUP 5
SRR1766481.9498920 chr10 445341 N chr10 445983 N DEL 5
SRR1766481.4941671 chr10 446044 N chr10 446470 N DUP 5
SRR1766481.3847918 chr10 445338 N chr10 446106 N DEL 3
SRR1766481.2189223 chr10 446258 N chr10 446430 N DEL 8
SRR1766446.5387252 chr10 445895 N chr10 446152 N DEL 10
SRR1766453.7989282 chr10 445372 N chr10 446183 N DEL 8
SRR1766462.6090865 chr10 445323 N chr10 446304 N DUP 5
SRR1766485.9694072 chr10 445664 N chr10 446304 N DUP 7
SRR1766468.5257295 chr10 445349 N chr10 446328 N DUP 7
SRR1766442.5185506 chr10 445349 N chr10 446328 N DUP 7
SRR1766457.4744247 chr10 445349 N chr10 446328 N DUP 7
SRR1766463.8155675 chr10 445340 N chr10 446280 N DEL 2
SRR1766467.8666729 chr10 445335 N chr10 446318 N DEL 7
SRR1766477.2867550 chr10 445336 N chr10 446319 N DEL 6
SRR1766475.7051580 chr10 445971 N chr10 446441 N DEL 6
SRR1766444.3877225 chr10 445542 N chr10 446440 N DEL 2
SRR1766478.2911725 chr10 446232 N chr10 446532 N DEL 5
SRR1766474.7762182 chr22 10628986 N chr22 10629091 N DEL 7
SRR1766472.4128835 chr22 10629003 N chr22 10629082 N DEL 15
SRR1766452.2375989 chr22 10629003 N chr22 10629082 N DEL 15
SRR1766481.3867815 chr22 10629003 N chr22 10629082 N DEL 7
SRR1766461.5487043 chr17 8052859 N chr17 8053469 N DEL 5
SRR1766455.8976567 chr17 8052874 N chr17 8053468 N DEL 1
SRR1766484.7792505 chr17 8052874 N chr17 8053468 N DEL 4
SRR1766467.3051340 chr17 8052954 N chr17 8053049 N DEL 4
SRR1766455.8706832 chr17 8052954 N chr17 8053049 N DEL 11
SRR1766485.6518993 chr17 8052954 N chr17 8053049 N DEL 12
SRR1766484.9768915 chr17 8052954 N chr17 8053049 N DEL 13
SRR1766465.1484519 chr17 8052954 N chr17 8053049 N DEL 13
SRR1766485.11491048 chr17 8052954 N chr17 8053049 N DEL 8
SRR1766454.10234852 chr17 8052954 N chr17 8053049 N DEL 13
SRR1766456.1296154 chr17 8052954 N chr17 8053049 N DEL 13
SRR1766477.10216605 chr17 8052839 N chr17 8052901 N DEL 1
SRR1766445.5835371 chr17 8052838 N chr17 8052900 N DEL 2
SRR1766467.10438200 chr17 8052838 N chr17 8052900 N DEL 2
SRR1766476.5707643 chr17 8052839 N chr17 8052959 N DEL 3
SRR1766452.10404207 chr17 8053023 N chr17 8053112 N DEL 13
SRR1766484.3957709 chr17 8053007 N chr17 8053114 N DEL 13
SRR1766461.1212597 chr17 8052989 N chr17 8053124 N DEL 1
SRR1766486.4365436 chr17 8053010 N chr17 8053117 N DEL 10
SRR1766467.7067754 chr17 8052829 N chr17 8053240 N DUP 5
SRR1766448.8630962 chr17 8052848 N chr17 8053257 N DEL 15
SRR1766442.32287039 chr17 8053212 N chr17 8053459 N DUP 2
SRR1766465.10171917 chr17 8052830 N chr17 8053477 N DEL 9
SRR1766484.10493353 chr17 8052831 N chr17 8053478 N DEL 9
SRR1766460.9927759 chr17 8052832 N chr17 8053479 N DEL 8
SRR1766442.40272481 chr8 35305711 N chr8 35305885 N DEL 7
SRR1766451.6944760 chr8 35305719 N chr8 35305931 N DEL 13
SRR1766470.7577762 chr8 35305750 N chr8 35305809 N DUP 2
SRR1766450.5749504 chr8 35305751 N chr8 35305810 N DUP 2
SRR1766447.5749196 chr8 35305752 N chr8 35305811 N DUP 1
SRR1766449.9118938 chr19 3988963 N chr19 3989266 N DEL 10
SRR1766450.4700379 chr19 3988752 N chr19 3989056 N DEL 18
SRR1766485.9498363 chr19 3988750 N chr19 3989054 N DEL 8
SRR1766483.11999385 chr19 3988888 N chr19 3989189 N DUP 5
SRR1766452.3959367 chr19 3989011 N chr19 3989312 N DUP 3
SRR1766473.2561787 chr19 3989015 N chr19 3989317 N DUP 4
SRR1766442.41839893 chr19 3989030 N chr19 3989336 N DEL 5
SRR1766481.8708133 chr19 3989084 N chr19 3989384 N DEL 10
SRR1766442.15552778 chr19 34534847 N chr19 34534916 N DUP 21
SRR1766470.5214552 chr19 34534869 N chr19 34534942 N DUP 31
SRR1766472.2362149 chr19 34534867 N chr19 34534928 N DUP 32
SRR1766463.9286562 chr6 132349571 N chr6 132349634 N DEL 7
SRR1766473.10628115 chr6 132349571 N chr6 132349634 N DEL 7
SRR1766471.3184750 chr6 132349571 N chr6 132349634 N DEL 7
SRR1766450.8242399 chr6 132349571 N chr6 132349634 N DEL 7
SRR1766467.6821127 chr6 132349571 N chr6 132349634 N DEL 7
SRR1766468.6140808 chr6 132349560 N chr6 132349639 N DEL 7
SRR1766457.2210040 chr6 132349561 N chr6 132349640 N DEL 7
SRR1766462.6011819 chr6 132349563 N chr6 132349642 N DEL 7
SRR1766472.7887842 chr6 132349563 N chr6 132349642 N DEL 7
SRR1766483.12324950 chr6 132349563 N chr6 132349642 N DEL 7
SRR1766454.3426803 chr6 132349564 N chr6 132349643 N DEL 6
SRR1766458.6598586 chr3 159680679 N chr3 159680788 N DUP 5
SRR1766470.8166299 chr3 159680679 N chr3 159680788 N DUP 5
SRR1766485.4147163 chr3 159680679 N chr3 159680788 N DUP 5
SRR1766486.4425722 chr3 159680679 N chr3 159680823 N DUP 1
SRR1766449.10330924 chr3 159680789 N chr3 159680851 N DUP 11
SRR1766442.21337461 chr3 159680771 N chr3 159680878 N DEL 12
SRR1766482.3744270 chr3 159680752 N chr3 159680887 N DUP 10
SRR1766466.3400024 chr3 159680684 N chr3 159680891 N DUP 8
SRR1766455.9153626 chr3 159680839 N chr3 159680899 N DUP 21
SRR1766476.7357564 chr3 159680839 N chr3 159680899 N DUP 21
SRR1766484.3109046 chr3 159680738 N chr3 159680865 N DEL 14
SRR1766482.5195377 chr3 159680689 N chr3 159680880 N DEL 2
SRR1766473.1131139 chr3 159680798 N chr3 159680884 N DEL 5
SRR1766459.863560 chr3 159680799 N chr3 159680885 N DEL 4
SRR1766471.8220520 chr14 27552285 N chr14 27552427 N DEL 1
SRR1766451.4879747 chr14 27552285 N chr14 27552427 N DEL 2
SRR1766482.2716203 chr14 27552285 N chr14 27552427 N DEL 4
SRR1766461.3468532 chr14 27552285 N chr14 27552427 N DEL 4
SRR1766460.5375918 chr14 27552264 N chr14 27552412 N DUP 1
SRR1766446.2359333 chr14 27552264 N chr14 27552412 N DUP 5
SRR1766448.8389810 chr14 27552264 N chr14 27552412 N DUP 6
SRR1766474.10196249 chr14 27552264 N chr14 27552412 N DUP 6
SRR1766448.10566826 chr11 112324043 N chr11 112325032 N DEL 29
SRR1766473.3617786 chr11 112324162 N chr11 112325149 N DUP 2
SRR1766444.2614570 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766481.7287039 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766477.8427562 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766444.5666643 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766470.9780305 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766474.1238218 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766463.142400 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766470.8409529 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766457.5925607 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766459.2401871 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766453.5746792 chr5 47101365 N chr5 47101567 N DEL 5
SRR1766485.5090024 chr5 47101381 N chr5 47101581 N DUP 3
SRR1766485.1649344 chr5 47101246 N chr5 47101418 N DEL 4
SRR1766455.9467542 chr7 1009084 N chr7 1009169 N DUP 8
SRR1766465.8793087 chrX 72179191 N chrX 72179359 N DEL 15
SRR1766474.3696003 chrX 72179191 N chrX 72179359 N DEL 15
SRR1766473.523687 chrX 72179191 N chrX 72179359 N DEL 20
SRR1766465.10238656 chrX 72179169 N chrX 72179295 N DUP 5
SRR1766461.8066145 chrX 72179282 N chrX 72179448 N DUP 3
SRR1766452.440472 chrX 72179281 N chrX 72179447 N DUP 4
SRR1766450.3422374 chrX 72179206 N chrX 72179334 N DEL 5
SRR1766472.452723 chrX 72179207 N chrX 72179374 N DUP 7
SRR1766453.2661435 chrX 72179226 N chrX 72179392 N DUP 5
SRR1766469.11020599 chr20 14771807 N chr20 14771895 N DEL 7
SRR1766465.980054 chr10 25241305 N chr10 25241421 N DEL 1
SRR1766477.11008970 chr10 25241326 N chr10 25241398 N DUP 13
SRR1766483.6279612 chr10 25241326 N chr10 25241407 N DUP 3
SRR1766444.6785179 chr10 25241326 N chr10 25241407 N DUP 5
SRR1766467.7692096 chr10 25241351 N chr10 25241429 N DEL 13
SRR1766460.3490834 chr10 25241352 N chr10 25241430 N DEL 12
SRR1766476.9861398 chr10 25241351 N chr10 25241429 N DEL 14
SRR1766465.5937100 chr10 25241374 N chr10 25241443 N DEL 1
SRR1766462.4679468 chr10 25241374 N chr10 25241458 N DEL 1
SRR1766463.1550588 chr10 25241374 N chr10 25241458 N DEL 1
SRR1766475.2784346 chr10 25241374 N chr10 25241458 N DEL 1
SRR1766449.7912842 chr10 25241473 N chr10 25241529 N DEL 6
SRR1766445.6555185 chr1 248754525 N chr1 248754644 N DUP 5
SRR1766442.39598688 chr6 115855883 N chr6 115856003 N DEL 5
SRR1766468.1198636 chr1 151601112 N chr1 151601283 N DEL 5
SRR1766476.1574992 chr11 68861420 N chr11 68861577 N DEL 10
SRR1766445.1506283 chrX 40236888 N chrX 40237189 N DEL 3
SRR1766448.3072456 chrX 40236844 N chrX 40237012 N DEL 11
SRR1766471.8463675 chrX 40236845 N chrX 40237146 N DEL 2
SRR1766471.3707342 chr11 68389759 N chr11 68389870 N DUP 5
SRR1766459.3891938 chr3 143449009 N chr3 143449278 N DEL 2
SRR1766479.8543740 chr3 143449009 N chr3 143449278 N DEL 2
SRR1766446.7241564 chr3 143449009 N chr3 143449278 N DEL 2
SRR1766458.7899287 chr3 143449009 N chr3 143449278 N DEL 2
SRR1766483.4632720 chr3 143449009 N chr3 143449278 N DEL 2
SRR1766485.6598329 chr3 143449252 N chr3 143449760 N DEL 28
SRR1766445.9416049 chr3 143449252 N chr3 143449760 N DEL 19
SRR1766464.5327466 chr3 143449252 N chr3 143449760 N DEL 19
SRR1766447.6856747 chr3 143449252 N chr3 143449760 N DEL 16
SRR1766455.391530 chr3 143449252 N chr3 143449760 N DEL 16
SRR1766461.9614609 chr3 143449198 N chr3 143449763 N DEL 18
SRR1766460.2179095 chr3 143449252 N chr3 143449760 N DEL 19
SRR1766473.7367585 chr3 143449196 N chr3 143449760 N DEL 17
SRR1766452.939341 chr3 143449536 N chr3 143449697 N DUP 26
SRR1766486.2874702 chr3 143449617 N chr3 143449670 N DEL 22
SRR1766479.8359576 chr3 143449794 N chr3 143449872 N DUP 34
SRR1766479.5543580 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766469.10897100 chr3 143449198 N chr3 143449763 N DEL 18
SRR1766461.682331 chr3 143449198 N chr3 143449763 N DEL 18
SRR1766481.7765743 chr3 143449760 N chr3 143449866 N DUP 33
SRR1766484.691538 chr3 143449201 N chr3 143449794 N DEL 22
SRR1766475.8273833 chr3 143449133 N chr3 143449810 N DUP 14
SRR1766473.5147936 chr3 143449234 N chr3 143449799 N DEL 15
SRR1766462.3324729 chr3 143449198 N chr3 143449763 N DEL 19
SRR1766472.441327 chr3 143449763 N chr3 143449874 N DUP 23
SRR1766462.1510450 chr3 143449763 N chr3 143449874 N DUP 12
SRR1766464.6039803 chr3 143449133 N chr3 143449810 N DUP 14
SRR1766447.9621093 chr3 143449763 N chr3 143449874 N DUP 23
SRR1766475.10552202 chr3 143449763 N chr3 143449874 N DUP 12
SRR1766477.4764861 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766462.3480851 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766465.11120355 chr3 143449763 N chr3 143449846 N DUP 22
SRR1766475.2600938 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766484.2298927 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766473.5033895 chr3 143449493 N chr3 143449632 N DUP 19
SRR1766460.1120946 chr3 143449806 N chr3 143449860 N DUP 24
SRR1766465.928632 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766475.6857724 chr3 143449750 N chr3 143449847 N DEL 19
SRR1766442.22868292 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766446.3454657 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766482.12637828 chr3 143449763 N chr3 143449846 N DUP 24
SRR1766470.2228423 chr3 143449056 N chr3 143449826 N DEL 10
SRR1766460.10366069 chr3 143449170 N chr3 143449847 N DEL 7
SRR1766447.3401251 chr3 143450052 N chr3 143450294 N DEL 10
SRR1766465.10431200 chr3 143450052 N chr3 143450294 N DEL 11
SRR1766475.8623921 chr3 143449024 N chr3 143450073 N DEL 7
SRR1766447.3052968 chr7 49549937 N chr7 49550053 N DUP 1
SRR1766469.1639010 chr7 49549937 N chr7 49550053 N DUP 1
SRR1766457.2050852 chr11 104791456 N chr11 104791564 N DUP 5
SRR1766442.22311336 chr11 104791455 N chr11 104791563 N DUP 6
SRR1766481.10440938 chr11 104791539 N chr11 104791655 N DUP 12
SRR1766469.6294988 chr6 53305377 N chr6 53305456 N DEL 5
SRR1766458.5708386 chr6 53305267 N chr6 53305538 N DUP 5
SRR1766442.5134074 chr6 53305480 N chr6 53305531 N DEL 5
SRR1766484.7602924 chr6 53305275 N chr6 53305373 N DEL 1
SRR1766473.11544000 chr6 53305249 N chr6 53305520 N DUP 4
SRR1766477.5647143 chr6 53305306 N chr6 53305483 N DEL 6
SRR1766442.17257380 chr11 97618072 N chr11 97618155 N DUP 1
SRR1766443.10490666 chr11 97618072 N chr11 97618155 N DUP 1
SRR1766475.9821077 chr11 97618107 N chr11 97618192 N DEL 5
SRR1766477.1661476 chr11 97618107 N chr11 97618192 N DEL 5
SRR1766482.7612192 chr11 97618107 N chr11 97618192 N DEL 5
SRR1766484.826956 chr11 97618107 N chr11 97618192 N DEL 5
SRR1766479.6536326 chr11 97618107 N chr11 97618192 N DEL 5
SRR1766471.10141258 chr11 97618107 N chr11 97618192 N DEL 5
SRR1766467.7048783 chr2 98004792 N chr2 98004907 N DUP 5
SRR1766442.42910138 chr2 241628894 N chr2 241629075 N DEL 10
SRR1766464.2059090 chr18 54780343 N chr18 54780565 N DUP 1
SRR1766484.4295285 chr18 54780415 N chr18 54780468 N DUP 6
SRR1766479.6971516 chr18 54780415 N chr18 54780468 N DUP 7
SRR1766445.5066877 chr18 54780415 N chr18 54780468 N DUP 7
SRR1766456.6187668 chr18 54780415 N chr18 54780468 N DUP 7
SRR1766459.9353751 chr18 54780415 N chr18 54780468 N DUP 7
SRR1766476.7605267 chr18 54780415 N chr18 54780468 N DUP 7
SRR1766471.3750461 chr18 54780320 N chr18 54780475 N DUP 7
SRR1766449.9045870 chr18 54780320 N chr18 54780475 N DUP 7
SRR1766449.8666212 chr18 54780375 N chr18 54780531 N DEL 32
SRR1766453.4893866 chr18 54780375 N chr18 54780531 N DEL 32
SRR1766469.10985631 chr18 54780375 N chr18 54780531 N DEL 32
SRR1766460.4061683 chr18 54780375 N chr18 54780531 N DEL 25
SRR1766465.7690096 chr18 54780355 N chr18 54780511 N DEL 5
SRR1766467.4495956 chr18 54780358 N chr18 54780548 N DEL 4
SRR1766464.10089509 chr18 54780373 N chr18 54780597 N DEL 5
SRR1766452.10635577 chr18 54780361 N chr18 54780619 N DEL 10
SRR1766485.123234 chr4 118792199 N chr4 118792354 N DUP 1
SRR1766462.627304 chr4 118792244 N chr4 118792360 N DUP 2
SRR1766448.9002135 chr4 118792319 N chr4 118792478 N DUP 3
SRR1766453.10984088 chr12 39712580 N chr12 39712641 N DEL 5
SRR1766452.6416423 chr12 39712944 N chr12 39713207 N DEL 4
SRR1766475.4798919 chr12 39712944 N chr12 39713207 N DEL 4
SRR1766447.10675052 chr12 39712764 N chr12 39712865 N DEL 5
SRR1766473.7469161 chr12 39713050 N chr12 39713147 N DEL 6
SRR1766457.181046 chr12 39713053 N chr12 39713150 N DEL 3
SRR1766477.5521377 chr12 39713054 N chr12 39713151 N DEL 2
SRR1766475.2950261 chr12 39713044 N chr12 39713141 N DEL 12
SRR1766452.5669320 chr12 39713048 N chr12 39713145 N DEL 8
SRR1766477.5568562 chr12 39713045 N chr12 39713142 N DEL 11
SRR1766474.10390654 chr12 39712718 N chr12 39713275 N DUP 1
SRR1766456.680911 chr12 39712718 N chr12 39713275 N DUP 2
SRR1766474.5119959 chr12 39712718 N chr12 39713275 N DUP 2
SRR1766443.10757029 chr12 39712718 N chr12 39713275 N DUP 4
SRR1766471.1403433 chr12 39712718 N chr12 39713275 N DUP 4
SRR1766468.2239782 chr12 39712937 N chr12 39713284 N DUP 5
SRR1766474.3725297 chr12 39712968 N chr12 39713175 N DEL 14
SRR1766443.1171953 chr12 39713207 N chr12 39713385 N DUP 5
SRR1766464.4222708 chr17 47666647 N chr17 47666705 N DEL 10
SRR1766483.719063 chr17 47666598 N chr17 47666712 N DEL 3
SRR1766442.11506670 chr17 47666598 N chr17 47666712 N DEL 3
SRR1766485.6315508 chr17 47666598 N chr17 47666712 N DEL 3
SRR1766471.5538539 chr6 169957126 N chr6 169957298 N DEL 32
SRR1766455.6471980 chr6 169957128 N chr6 169957470 N DUP 8
SRR1766485.3558276 chr6 169957191 N chr6 169957500 N DUP 5
SRR1766485.9785545 chr6 169957309 N chr6 169957483 N DEL 22
SRR1766442.27253793 chr17 77245705 N chr17 77245937 N DUP 2
SRR1766450.7135947 chr17 77245705 N chr17 77245937 N DUP 2
SRR1766465.9291878 chr1 54561847 N chr1 54561899 N DEL 1
SRR1766481.8488102 chr1 54561847 N chr1 54561899 N DEL 1
SRR1766446.6391202 chr1 54561802 N chr1 54561979 N DUP 1
SRR1766448.8229826 chr1 54561795 N chr1 54561872 N DUP 8
SRR1766465.3894749 chr1 54561848 N chr1 54561947 N DUP 1
SRR1766485.8042020 chr1 54561860 N chr1 54561910 N DUP 3
SRR1766476.4480691 chr1 54561876 N chr1 54561926 N DUP 5
SRR1766442.18831192 chr11 47657874 N chr11 47658177 N DUP 12
SRR1766450.10776393 chr6 72549379 N chr6 72549449 N DEL 7
SRR1766452.5608229 chr6 72549379 N chr6 72549449 N DEL 7
SRR1766457.7630323 chr6 72549351 N chr6 72549452 N DEL 7
SRR1766458.2129122 chr7 100994660 N chr7 100995414 N DEL 4
SRR1766484.9679993 chr7 100994891 N chr7 100995645 N DEL 1
SRR1766454.3516641 chr7 100995098 N chr7 100995846 N DEL 20
SRR1766463.8817437 chr7 100995441 N chr7 100996112 N DEL 12
SRR1766479.7732507 chr7 100994654 N chr7 100995408 N DEL 25
SRR1766484.9679993 chr7 100994880 N chr7 100995634 N DEL 5
SRR1766448.10527086 chr7 100995159 N chr7 100995905 N DUP 5
SRR1766442.2648770 chr7 100995188 N chr7 100995936 N DEL 15
SRR1766483.11632997 chr10 126947762 N chr10 126948129 N DUP 8
SRR1766467.8370489 chr10 126947606 N chr10 126948140 N DUP 16
SRR1766458.555154 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766461.5131769 chr10 126947530 N chr10 126947597 N DUP 5
SRR1766470.10721999 chr10 126947572 N chr10 126947673 N DUP 8
SRR1766477.10149820 chr10 126947472 N chr10 126947538 N DEL 5
SRR1766451.354427 chr10 126947687 N chr10 126948090 N DEL 8
SRR1766442.9147252 chr10 126947990 N chr10 126948158 N DEL 5
SRR1766474.10666715 chr10 126947492 N chr10 126948056 N DEL 8
SRR1766442.45877426 chr10 126947469 N chr10 126948130 N DUP 8
SRR1766462.3225095 chr10 126947499 N chr10 126947633 N DEL 10
SRR1766485.8842533 chr10 126947994 N chr10 126948128 N DEL 5
SRR1766477.8399702 chr10 126947543 N chr10 126947612 N DEL 5
SRR1766478.1945089 chr10 126947489 N chr10 126947855 N DEL 5
SRR1766476.4085486 chr10 126947496 N chr10 126947792 N DUP 6
SRR1766455.9689092 chr10 126947496 N chr10 126948194 N DUP 11
SRR1766467.395444 chr10 126947520 N chr10 126947626 N DEL 9
SRR1766457.3935298 chr10 126947455 N chr10 126947855 N DEL 5
SRR1766445.4136760 chr10 126947597 N chr10 126947861 N DEL 6
SRR1766470.1317365 chr10 126947489 N chr10 126948090 N DEL 10
SRR1766483.11886053 chr10 126948175 N chr10 126948579 N DUP 5
SRR1766444.6514218 chr10 126947529 N chr10 126947598 N DEL 13
SRR1766452.10600804 chr10 126947693 N chr10 126947895 N DEL 11
SRR1766457.1930471 chr10 126947489 N chr10 126947855 N DEL 5
SRR1766457.610347 chr10 126947509 N chr10 126948244 N DUP 2
SRR1766466.3611394 chr10 126947499 N chr10 126947928 N DUP 5
SRR1766480.8125341 chr10 126947464 N chr10 126947663 N DEL 8
SRR1766482.4257835 chr10 126947490 N chr10 126948157 N DUP 5
SRR1766479.4026998 chr10 126947448 N chr10 126947548 N DEL 5
SRR1766451.5432020 chr10 126947458 N chr10 126948161 N DEL 5
SRR1766473.5220858 chr10 126947490 N chr10 126947888 N DUP 5
SRR1766472.8565400 chr10 126947730 N chr10 126948093 N DEL 6
SRR1766442.35767887 chr10 126947499 N chr10 126947928 N DUP 5
SRR1766452.10369077 chr10 126947463 N chr10 126947529 N DEL 4
SRR1766480.4291980 chr10 126947473 N chr10 126947673 N DUP 8
SRR1766456.5088505 chr10 126947625 N chr10 126948056 N DEL 10
SRR1766456.3914509 chr10 126947492 N chr10 126948056 N DEL 5
SRR1766458.1373923 chr10 126947464 N chr10 126948096 N DEL 10
SRR1766473.4331467 chr10 126947439 N chr10 126948341 N DUP 13
SRR1766449.2965602 chr10 126947761 N chr10 126948130 N DEL 11
SRR1766456.2051834 chr10 126947663 N chr10 126947894 N DUP 3
SRR1766452.10414938 chr10 126947663 N chr10 126947996 N DUP 10
SRR1766481.10877174 chr10 126947668 N chr10 126948569 N DEL 16
SRR1766457.3731415 chr10 126947472 N chr10 126947538 N DEL 5
SRR1766468.7456308 chr10 126947597 N chr10 126948266 N DEL 5
SRR1766472.11832695 chr10 126947950 N chr10 126948087 N DEL 15
SRR1766466.8834071 chr10 126947673 N chr10 126948172 N DEL 5
SRR1766483.12098475 chr10 126947507 N chr10 126948579 N DUP 5
SRR1766482.1453658 chr10 126947653 N chr10 126948087 N DEL 10
SRR1766455.3007093 chr10 126947429 N chr10 126947495 N DEL 1
SRR1766461.2602655 chr10 126947460 N chr10 126948197 N DEL 8
SRR1766448.2098654 chr10 126947956 N chr10 126948087 N DEL 6
SRR1766478.949831 chr10 126947599 N chr10 126948135 N DEL 4
SRR1766455.5821830 chr10 126947524 N chr10 126947953 N DUP 13
SRR1766483.11956179 chr10 126947464 N chr10 126948096 N DEL 9
SRR1766457.2896017 chr10 126948070 N chr10 126948140 N DUP 16
SRR1766462.7337065 chr10 126947495 N chr10 126948164 N DEL 8
SRR1766453.4111581 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766477.4962088 chr10 126947990 N chr10 126948192 N DEL 5
SRR1766442.21048004 chr10 126947576 N chr10 126948072 N DEL 16
SRR1766477.9586863 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766442.27314618 chr10 126947416 N chr10 126947483 N DUP 8
SRR1766473.1955765 chr10 126947544 N chr10 126947611 N DUP 2
SRR1766453.1082407 chr10 126947426 N chr10 126948257 N DUP 8
SRR1766445.1052700 chr10 126947490 N chr10 126947823 N DUP 8
SRR1766442.16115804 chr10 126947409 N chr10 126948379 N DUP 7
SRR1766464.9036473 chr10 126947430 N chr10 126948062 N DEL 9
SRR1766442.10638994 chr10 126947433 N chr10 126947830 N DEL 1
SRR1766479.13749124 chr10 126947530 N chr10 126947597 N DUP 5
SRR1766442.31900206 chr10 126948056 N chr10 126948358 N DUP 10
SRR1766484.11182107 chr10 126947537 N chr10 126947835 N DEL 5
SRR1766442.42176567 chr10 126947566 N chr10 126948199 N DUP 1
SRR1766449.649800 chr10 126947543 N chr10 126947841 N DEL 6
SRR1766464.7980941 chr10 126947820 N chr10 126948158 N DEL 5
SRR1766464.2222563 chr10 126947490 N chr10 126947922 N DUP 5
SRR1766486.10124266 chr10 126947622 N chr10 126948124 N DEL 8
SRR1766456.6130326 chr10 126947478 N chr10 126947547 N DEL 8
SRR1766483.10016097 chr10 126947461 N chr10 126948130 N DEL 2
SRR1766473.252871 chr10 126947524 N chr10 126948355 N DUP 10
SRR1766481.8098107 chr10 126947416 N chr10 126947650 N DUP 3
SRR1766468.1270051 chr10 126947979 N chr10 126948244 N DUP 13
SRR1766442.24868651 chr10 126947545 N chr10 126947843 N DEL 4
SRR1766484.3945647 chr10 126947791 N chr10 126948189 N DUP 10
SRR1766480.1000689 chr10 126947492 N chr10 126948056 N DEL 5
SRR1766442.42623292 chr10 126947538 N chr10 126947605 N DUP 5
SRR1766470.7343366 chr10 126947426 N chr10 126948189 N DUP 8
SRR1766453.3517703 chr10 126947567 N chr10 126948231 N DUP 4
SRR1766455.7700498 chr10 126947462 N chr10 126948060 N DEL 10
SRR1766479.2768839 chr10 126947605 N chr10 126948141 N DEL 8
SRR1766442.43338461 chr10 126947854 N chr10 126948056 N DEL 10
SRR1766484.1019600 chr10 126947589 N chr10 126948295 N DEL 8
SRR1766471.5691776 chr10 126947597 N chr10 126947861 N DEL 10
SRR1766442.24107140 chr10 126947589 N chr10 126947984 N DUP 11
SRR1766448.10407175 chr10 126947492 N chr10 126947657 N DEL 4
SRR1766457.2066579 chr10 126948129 N chr10 126948266 N DEL 8
SRR1766475.2606893 chr10 126947659 N chr10 126948056 N DEL 9
SRR1766465.2860578 chr10 126947524 N chr10 126947919 N DUP 13
SRR1766472.3276333 chr10 126947538 N chr10 126947605 N DUP 1
SRR1766473.6500454 chr10 126947496 N chr10 126948160 N DUP 11
SRR1766467.2230867 chr10 126947523 N chr10 126948056 N DEL 5
SRR1766479.11123758 chr10 126947415 N chr10 126948183 N DEL 5
SRR1766469.9360861 chr10 126947640 N chr10 126948174 N DUP 19
SRR1766472.8074599 chr10 126948001 N chr10 126948135 N DEL 5
SRR1766457.3990525 chr10 126947557 N chr10 126948121 N DEL 7
SRR1766479.13198733 chr10 126947855 N chr10 126947990 N DUP 5
SRR1766458.8509787 chr10 126947600 N chr10 126947830 N DEL 2
SRR1766450.3366031 chr10 126947408 N chr10 126947839 N DEL 5
SRR1766478.9289682 chr10 126948065 N chr10 126948129 N DUP 10
SRR1766442.24567591 chr10 126947654 N chr10 126948021 N DUP 7
SRR1766484.3775872 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766463.5343559 chr10 126947422 N chr10 126947591 N DUP 11
SRR1766475.1142021 chr10 126947557 N chr10 126948056 N DEL 4
SRR1766448.5193566 chr10 126947397 N chr10 126948194 N DUP 5
SRR1766450.4248701 chr10 126947557 N chr10 126948087 N DEL 6
SRR1766442.46552120 chr10 126947416 N chr10 126947483 N DUP 5
SRR1766450.661936 chr10 126947538 N chr10 126947837 N DUP 5
SRR1766464.8723702 chr10 126947456 N chr10 126948191 N DUP 19
SRR1766443.3456646 chr10 126947595 N chr10 126948299 N DUP 3
SRR1766462.816657 chr10 126947792 N chr10 126948162 N DUP 10
SRR1766457.1872434 chr10 126947623 N chr10 126948159 N DEL 5
SRR1766442.2725432 chr10 126947423 N chr10 126947623 N DUP 5
SRR1766458.6555825 chr10 126947554 N chr10 126947855 N DEL 13
SRR1766468.7633593 chr10 126947538 N chr10 126947639 N DUP 5
SRR1766443.5778745 chr10 126947496 N chr10 126947665 N DUP 5
SRR1766471.3984614 chr10 126947538 N chr10 126947605 N DUP 5
SRR1766479.2470933 chr10 126947598 N chr10 126947894 N DUP 5
SRR1766465.11046082 chr10 126947589 N chr10 126947653 N DUP 5
SRR1766473.9671552 chr10 126947467 N chr10 126947762 N DEL 16
SRR1766474.1531488 chr10 126947619 N chr10 126948155 N DEL 8
SRR1766458.5078900 chr10 126947983 N chr10 126948568 N DEL 10
SRR1766442.22480633 chr10 126947529 N chr10 126947599 N DUP 7
SRR1766452.6390281 chr10 126947855 N chr10 126948154 N DUP 8
SRR1766479.5754455 chr10 126947540 N chr10 126947601 N DUP 3
SRR1766447.9458120 chr10 126947438 N chr10 126947835 N DEL 5
SRR1766464.2863251 chr10 126947894 N chr10 126947963 N DEL 5
SRR1766446.4487313 chr10 126947497 N chr10 126947796 N DUP 11
SRR1766466.9820928 chr10 126947464 N chr10 126947598 N DEL 5
SRR1766478.5901306 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766470.1295928 chr10 126947415 N chr10 126947682 N DEL 5
SRR1766443.10323761 chr10 126947458 N chr10 126948155 N DEL 11
SRR1766462.8095013 chr10 126947602 N chr10 126948064 N DEL 9
SRR1766442.18391058 chr10 126947600 N chr10 126948569 N DEL 16
SRR1766466.5575506 chr10 126947538 N chr10 126947605 N DUP 9
SRR1766444.308462 chr10 126947588 N chr10 126947652 N DUP 8
SRR1766472.1730732 chr10 126947498 N chr10 126948164 N DEL 5
SRR1766470.1057442 chr10 126947538 N chr10 126947602 N DUP 10
SRR1766456.2981003 chr10 126947492 N chr10 126947589 N DEL 14
SRR1766460.3588091 chr10 126947597 N chr10 126947861 N DEL 6
SRR1766451.8791147 chr10 126948056 N chr10 126948358 N DUP 10
SRR1766484.5083173 chr10 126947431 N chr10 126948163 N DUP 8
SRR1766456.3242720 chr10 126947472 N chr10 126948073 N DEL 15
SRR1766467.403934 chr10 126947489 N chr10 126947889 N DEL 5
SRR1766443.9825540 chr10 126947586 N chr10 126947981 N DUP 13
SRR1766468.5746192 chr10 126947492 N chr10 126948087 N DEL 14
SRR1766481.12493910 chr10 126947422 N chr10 126947758 N DUP 11
SRR1766486.3310028 chr10 126947438 N chr10 126947538 N DEL 5
SRR1766463.4334193 chr10 126947612 N chr10 126948074 N DEL 15
SRR1766447.3414984 chr10 126947656 N chr10 126947855 N DEL 7
SRR1766464.10586500 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766467.5545917 chr10 126947394 N chr10 126947628 N DUP 5
SRR1766442.9760612 chr10 126947472 N chr10 126947538 N DEL 5
SRR1766464.10354857 chr10 126947560 N chr10 126948062 N DEL 10
SRR1766465.6816635 chr10 126947529 N chr10 126947700 N DEL 13
SRR1766476.7715033 chr10 126947490 N chr10 126948058 N DUP 10
SRR1766458.8980439 chr10 126947557 N chr10 126948056 N DEL 5
SRR1766479.6760768 chr10 126947555 N chr10 126948259 N DUP 16
SRR1766442.881293 chr10 126947627 N chr10 126948092 N DEL 5
SRR1766452.1086251 chr10 126947829 N chr10 126947998 N DUP 10
SRR1766464.1255277 chr10 126947499 N chr10 126947894 N DUP 5
SRR1766478.8754035 chr10 126947838 N chr10 126948579 N DUP 5
SRR1766457.708608 chr10 126947432 N chr10 126948064 N DEL 7
SRR1766463.5717642 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766476.9192109 chr10 126947690 N chr10 126948056 N DEL 10
SRR1766447.10618584 chr10 126947567 N chr10 126948197 N DUP 13
SRR1766448.6429749 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766476.6964575 chr10 126947490 N chr10 126947690 N DUP 10
SRR1766466.3200020 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766458.336152 chr10 126947492 N chr10 126947657 N DEL 8
SRR1766452.944221 chr10 126947458 N chr10 126948056 N DEL 9
SRR1766486.10354766 chr10 126947654 N chr10 126947919 N DUP 5
SRR1766483.8768564 chr10 126947490 N chr10 126947724 N DUP 10
SRR1766442.46766163 chr10 126947455 N chr10 126948192 N DEL 8
SRR1766480.7506955 chr10 126947439 N chr10 126948105 N DEL 5
SRR1766463.10781725 chr10 126947458 N chr10 126947688 N DEL 11
SRR1766464.9185707 chr10 126947461 N chr10 126947530 N DEL 10
SRR1766486.3159852 chr10 126947496 N chr10 126947665 N DUP 10
SRR1766442.35767887 chr10 126947529 N chr10 126948130 N DEL 2
SRR1766474.11220296 chr10 126947462 N chr10 126947565 N DEL 6
SRR1766466.10076539 chr10 126947455 N chr10 126948192 N DEL 8
SRR1766442.46106457 chr10 126947416 N chr10 126947483 N DUP 3
SRR1766476.5666329 chr10 126947524 N chr10 126947953 N DUP 13
SRR1766477.7448786 chr10 126947464 N chr10 126948099 N DEL 10
SRR1766449.1373511 chr10 126947472 N chr10 126947538 N DEL 5
SRR1766443.4519148 chr10 126947458 N chr10 126948056 N DEL 5
SRR1766483.8061414 chr10 126947687 N chr10 126947957 N DEL 11
SRR1766454.3067439 chr10 126947605 N chr10 126948098 N DEL 4
SRR1766464.10110510 chr10 126947490 N chr10 126947922 N DUP 5
SRR1766443.5137469 chr10 126947435 N chr10 126948101 N DEL 5
SRR1766455.7694475 chr10 126947523 N chr10 126948056 N DEL 5
SRR1766476.8762156 chr10 126947453 N chr10 126947553 N DEL 10
SRR1766468.2416860 chr10 126947436 N chr10 126947502 N DEL 3
SRR1766480.4180718 chr10 126947928 N chr10 126948065 N DEL 10
SRR1766467.3799356 chr10 126947854 N chr10 126948056 N DEL 10
SRR1766467.395444 chr10 126947439 N chr10 126948139 N DEL 5
SRR1766445.8895111 chr10 126948069 N chr10 126948133 N DUP 6
SRR1766443.4270624 chr10 126947631 N chr10 126948130 N DEL 5
SRR1766485.2246586 chr10 126947631 N chr10 126948133 N DEL 5
SRR1766481.7412743 chr10 126947417 N chr10 126948149 N DUP 7
SRR1766442.8092381 chr10 126947622 N chr10 126948158 N DEL 5
SRR1766479.12841830 chr10 126947597 N chr10 126947762 N DEL 8
SRR1766482.9325736 chr10 126947588 N chr10 126948090 N DEL 8
SRR1766459.7324251 chr10 126947409 N chr10 126947840 N DEL 5
SRR1766455.9053641 chr10 126947600 N chr10 126948569 N DEL 16
SRR1766460.4444383 chr10 126947492 N chr10 126948056 N DEL 6
SRR1766486.7105853 chr10 126948154 N chr10 126948294 N DEL 11
SRR1766454.6079038 chr10 126947492 N chr10 126948056 N DEL 5
SRR1766463.7227385 chr10 126947885 N chr10 126948090 N DEL 13
SRR1766484.5083173 chr10 126947854 N chr10 126948056 N DEL 10
SRR1766442.26434261 chr10 126947600 N chr10 126947697 N DEL 21
SRR1766477.10130098 chr10 126947473 N chr10 126947673 N DUP 14
SRR1766473.3618414 chr10 126947538 N chr10 126948137 N DUP 5
SRR1766461.9334837 chr10 126947553 N chr10 126948188 N DEL 3
SRR1766465.992590 chr10 126947455 N chr10 126948158 N DEL 5
SRR1766456.667337 chr10 126947659 N chr10 126948056 N DEL 6
SRR1766446.2763432 chr10 126947458 N chr10 126948056 N DEL 8
SRR1766481.8711825 chr10 126947542 N chr10 126947840 N DEL 7
SRR1766479.2834000 chr10 126947440 N chr10 126947837 N DEL 4
SRR1766458.6555825 chr10 126947554 N chr10 126948192 N DEL 13
SRR1766476.7878364 chr10 126947458 N chr10 126948087 N DEL 11
SRR1766480.7017878 chr10 126947436 N chr10 126947833 N DEL 4
SRR1766482.1413227 chr10 126947913 N chr10 126948081 N DEL 6
SRR1766473.5082680 chr10 126947619 N chr10 126948087 N DEL 10
SRR1766477.8680668 chr10 126947422 N chr10 126947984 N DUP 6
SRR1766474.6464341 chr10 126947467 N chr10 126947762 N DEL 11
SRR1766445.8873658 chr10 126947487 N chr10 126947687 N DUP 10
SRR1766447.3414984 chr10 126947537 N chr10 126948070 N DEL 10
SRR1766479.3811633 chr10 126947492 N chr10 126948056 N DEL 8
SRR1766466.6446607 chr10 126947464 N chr10 126947598 N DEL 5
SRR1766486.10086493 chr10 126947410 N chr10 126948144 N DEL 1
SRR1766486.703255 chr10 126947437 N chr10 126947834 N DEL 5
SRR1766464.1518048 chr10 126947437 N chr10 126948137 N DEL 5
SRR1766465.7527784 chr10 126947464 N chr10 126948065 N DEL 10
SRR1766479.2610269 chr10 126947601 N chr10 126947696 N DUP 13
SRR1766442.26515337 chr10 126947690 N chr10 126948056 N DEL 10
SRR1766467.4314972 chr10 126947489 N chr10 126947558 N DEL 5
SRR1766466.5228074 chr10 126947557 N chr10 126948022 N DEL 13
SRR1766475.5006454 chr10 126947551 N chr10 126948186 N DEL 1
SRR1766484.7170907 chr10 126947458 N chr10 126948056 N DEL 9
SRR1766447.9463604 chr10 126948030 N chr10 126948130 N DEL 10
SRR1766481.4694938 chr10 126947588 N chr10 126948294 N DEL 13
SRR1766442.20448537 chr10 126947499 N chr10 126947928 N DUP 5
SRR1766463.8960878 chr10 126947500 N chr10 126947637 N DEL 8
SRR1766476.3797964 chr10 126947526 N chr10 126947632 N DEL 13
SRR1766480.5125150 chr10 126947538 N chr10 126947868 N DUP 5
SRR1766474.8064010 chr10 126947762 N chr10 126947897 N DUP 11
SRR1766483.11217878 chr10 126947472 N chr10 126947538 N DEL 5
SRR1766444.4487769 chr10 126947464 N chr10 126948096 N DEL 5
SRR1766460.6774972 chr10 126947665 N chr10 126947929 N DEL 5
SRR1766478.6182520 chr10 126947632 N chr10 126947693 N DUP 15
SRR1766455.5952960 chr10 126947544 N chr10 126948247 N DEL 5
SRR1766453.4514866 chr10 126947567 N chr10 126948265 N DUP 7
SRR1766454.739332 chr10 126947996 N chr10 126948164 N DEL 4
SRR1766479.6988366 chr10 126947472 N chr10 126947538 N DEL 5
SRR1766442.8139622 chr10 126947490 N chr10 126947856 N DEL 5
SRR1766442.27847155 chr10 126947490 N chr10 126947659 N DUP 5
SRR1766482.5512073 chr10 126947442 N chr10 126948108 N DEL 5
SRR1766442.11016442 chr10 126947520 N chr10 126948090 N DEL 8
SRR1766463.10450632 chr10 126947589 N chr10 126947659 N DUP 16
SRR1766481.7736104 chr10 126947480 N chr10 126948348 N DUP 5
SRR1766463.172660 chr10 126947589 N chr10 126948321 N DUP 10
SRR1766453.9252034 chr10 126947623 N chr10 126947890 N DEL 10
SRR1766472.11290418 chr10 126947499 N chr10 126948197 N DUP 13
SRR1766482.1000987 chr10 126947625 N chr10 126948155 N DEL 11
SRR1766475.5089322 chr10 126947492 N chr10 126947756 N DEL 5
SRR1766457.2011452 chr10 126948087 N chr10 126948185 N DUP 15
SRR1766442.9696251 chr10 126947489 N chr10 126947855 N DEL 5
SRR1766461.6115088 chr10 126947489 N chr10 126948593 N DEL 22
SRR1766473.1787874 chr10 126947574 N chr10 126948176 N DUP 12
SRR1766454.5842197 chr10 126947608 N chr10 126948070 N DEL 16
SRR1766483.3461090 chr10 126947557 N chr10 126948056 N DEL 6
SRR1766450.7225942 chr10 126947523 N chr10 126948056 N DEL 5
SRR1766442.42354949 chr10 126947434 N chr10 126948234 N DUP 7
SRR1766475.5226263 chr10 126947464 N chr10 126948133 N DEL 5
SRR1766479.12517576 chr10 126947537 N chr10 126948070 N DEL 10
SRR1766482.6077681 chr10 126947461 N chr10 126947564 N DEL 5
SRR1766442.743146 chr10 126947479 N chr10 126948080 N DEL 15
SRR1766445.1530850 chr10 126947631 N chr10 126948133 N DEL 5
SRR1766459.7799527 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766447.4034789 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766466.8330554 chr10 126947928 N chr10 126948065 N DEL 10
SRR1766476.8738587 chr10 126947472 N chr10 126947538 N DEL 5
SRR1766486.3310028 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766460.1682100 chr10 126947416 N chr10 126948049 N DUP 10
SRR1766468.7633593 chr10 126947990 N chr10 126948124 N DEL 5
SRR1766466.3607113 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766485.11887715 chr10 126947492 N chr10 126947589 N DEL 6
SRR1766460.24420 chr10 126947990 N chr10 126948594 N DUP 8
SRR1766460.2510294 chr10 126947472 N chr10 126947538 N DEL 5
SRR1766479.7839205 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766465.3944793 chr10 126947461 N chr10 126948056 N DEL 13
SRR1766459.10666098 chr10 126947504 N chr10 126948341 N DUP 7
SRR1766467.3840542 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766469.7597183 chr10 126947998 N chr10 126948132 N DEL 10
SRR1766442.26250424 chr10 126947509 N chr10 126948043 N DUP 1
SRR1766468.3568200 chr10 126947625 N chr10 126948056 N DEL 10
SRR1766473.4539366 chr10 126947424 N chr10 126948056 N DEL 10
SRR1766474.10666715 chr10 126947461 N chr10 126948062 N DEL 5
SRR1766471.6935264 chr10 126947684 N chr10 126947988 N DEL 13
SRR1766442.35813991 chr10 126947458 N chr10 126948056 N DEL 10
SRR1766445.6817241 chr10 126947475 N chr10 126947774 N DUP 13
SRR1766456.2763124 chr10 126947408 N chr10 126947839 N DEL 5
SRR1766442.41498703 chr10 126947529 N chr10 126947666 N DEL 8
SRR1766452.5933781 chr10 126947692 N chr10 126948129 N DEL 12
SRR1766451.3133203 chr10 126947990 N chr10 126948158 N DEL 5
SRR1766470.6100919 chr10 126948073 N chr10 126948174 N DUP 10
SRR1766481.9683000 chr10 126947451 N chr10 126948120 N DEL 8
SRR1766470.2993009 chr10 126947499 N chr10 126947999 N DUP 3
SRR1766468.5746192 chr10 126947490 N chr10 126948157 N DUP 5
SRR1766483.800063 chr10 126947521 N chr10 126947659 N DUP 16
SRR1766449.8384614 chr10 126948090 N chr10 126948188 N DUP 10
SRR1766480.1095781 chr10 126947597 N chr10 126948062 N DEL 5
SRR1766483.6681557 chr10 126947697 N chr10 126948129 N DUP 8
SRR1766484.6915975 chr10 126947597 N chr10 126947762 N DEL 8
SRR1766479.1654671 chr10 126947434 N chr10 126947831 N DEL 2
SRR1766460.3588091 chr10 126947611 N chr10 126947841 N DEL 4
SRR1766463.10450632 chr10 126947467 N chr10 126948062 N DEL 13
SRR1766457.5185976 chr10 126947597 N chr10 126947861 N DEL 5
SRR1766478.6823772 chr10 126947830 N chr10 126948129 N DUP 5
SRR1766443.6461950 chr10 126947430 N chr10 126948130 N DEL 5
SRR1766485.8136446 chr10 126947436 N chr10 126948136 N DEL 5
SRR1766459.5707317 chr10 126947455 N chr10 126947855 N DEL 5
SRR1766445.8616746 chr10 126947458 N chr10 126947722 N DEL 6
SRR1766442.20389188 chr10 126947426 N chr10 126947954 N DUP 8
SRR1766446.54148 chr10 126947600 N chr10 126948569 N DEL 16
SRR1766473.332021 chr10 126947965 N chr10 126948569 N DEL 16
SRR1766449.10330771 chr10 126947489 N chr10 126947855 N DEL 5
SRR1766455.9583299 chr10 126947464 N chr10 126948130 N DEL 5
SRR1766470.8762546 chr10 126947422 N chr10 126947916 N DUP 8
SRR1766442.33223973 chr10 126947483 N chr10 126948118 N DEL 10
SRR1766484.2498783 chr10 126947490 N chr10 126947659 N DUP 5
SRR1766446.32319 chr10 126947929 N chr10 126948129 N DUP 5
SRR1766481.7736104 chr10 126947626 N chr10 126947990 N DUP 5
SRR1766469.7094554 chr10 126947557 N chr10 126948121 N DEL 16
SRR1766455.4480818 chr10 126947538 N chr10 126948585 N DUP 5
SRR1766473.9135770 chr10 126947560 N chr10 126947756 N DEL 19
SRR1766459.8682439 chr10 126947501 N chr10 126947599 N DUP 4
SRR1766447.9641406 chr10 126947966 N chr10 126948299 N DUP 1
SRR1766443.4926066 chr10 126947600 N chr10 126948569 N DEL 16
SRR1766460.8112376 chr10 126947520 N chr10 126947626 N DEL 9
SRR1766442.7834194 chr4 146008342 N chr4 146008432 N DEL 10
SRR1766445.10374695 chr4 146008376 N chr4 146008588 N DUP 8
SRR1766451.4265697 chr14 94591581 N chr14 94591647 N DEL 2
SRR1766455.6878962 chr9 95083489 N chr9 95083585 N DUP 10
SRR1766474.1715210 chr9 95083554 N chr9 95083677 N DUP 4
SRR1766473.11796588 chr15 29950339 N chr15 29950442 N DEL 6
SRR1766445.10202271 chr1 153261418 N chr1 153261509 N DEL 5
SRR1766442.1874461 chr1 153261450 N chr1 153261595 N DEL 3
SRR1766479.11752573 chr1 153261307 N chr1 153261633 N DUP 1
SRR1766442.33664634 chr11 59585617 N chr11 59585783 N DUP 1
SRR1766459.4254733 chr22 12571521 N chr22 12571575 N DEL 16
SRR1766484.8340491 chr19 31051650 N chr19 31051829 N DEL 3
SRR1766450.5235893 chr19 31051651 N chr19 31051830 N DEL 2
SRR1766456.6467327 chr2 187868327 N chr2 187868570 N DUP 5
SRR1766482.511069 chr2 187868470 N chr2 187868519 N DUP 5
SRR1766482.461356 chr14 65692405 N chr14 65692531 N DUP 5
SRR1766442.19355189 chr14 65692480 N chr14 65692579 N DEL 5
SRR1766453.9243517 chr14 65692378 N chr14 65692549 N DUP 9
SRR1766445.1669995 chr14 65692366 N chr14 65692494 N DEL 5
SRR1766481.4585224 chr14 65692481 N chr14 65692578 N DUP 2
SRR1766476.3763825 chr14 65692608 N chr14 65692659 N DEL 9
SRR1766451.2501926 chr14 65692608 N chr14 65692659 N DEL 11
SRR1766442.20100569 chr14 65692371 N chr14 65692595 N DUP 5
SRR1766442.11004184 chr14 65692530 N chr14 65692627 N DUP 5
SRR1766478.8939399 chr14 65692627 N chr14 65692680 N DEL 1
SRR1766476.8496447 chr14 65692388 N chr14 65692515 N DEL 7
SRR1766447.6442183 chr14 65692354 N chr14 65692627 N DUP 4
SRR1766473.5567176 chr14 65692608 N chr14 65692659 N DEL 11
SRR1766471.1461452 chr14 65692474 N chr14 65692620 N DUP 3
SRR1766447.4355277 chr14 65692474 N chr14 65692620 N DUP 2
SRR1766473.10421972 chr14 65692568 N chr14 65692665 N DUP 5
SRR1766460.4039312 chr14 65692475 N chr14 65692572 N DUP 8
SRR1766451.9326935 chr14 65692608 N chr14 65692659 N DEL 11
SRR1766477.3899820 chr14 65692692 N chr14 65692909 N DEL 9
SRR1766450.9586330 chr14 65692608 N chr14 65692659 N DEL 11
SRR1766486.1974416 chr14 65692559 N chr14 65692659 N DEL 11
SRR1766477.11545340 chr14 65692560 N chr14 65692660 N DEL 11
SRR1766460.1278588 chr14 65692558 N chr14 65692658 N DEL 11
SRR1766484.4796887 chr14 65692510 N chr14 65692659 N DEL 6
SRR1766446.2126669 chr14 65692510 N chr14 65692659 N DEL 6
SRR1766442.21052918 chr14 65692510 N chr14 65692659 N DEL 6
SRR1766449.1170484 chr14 65692388 N chr14 65692664 N DEL 6
SRR1766486.6223801 chr14 65692385 N chr14 65692712 N DEL 3
SRR1766458.8486522 chr14 65692424 N chr14 65692876 N DUP 3
SRR1766468.4303449 chr22 44264987 N chr22 44265047 N DEL 5
SRR1766486.11290209 chr10 52834578 N chr10 52834717 N DEL 12
SRR1766445.7941808 chr10 52834911 N chr10 52835518 N DEL 5
SRR1766446.10614688 chr10 52834357 N chr10 52835506 N DUP 16
SRR1766482.2724377 chr10 52834294 N chr10 52834592 N DEL 5
SRR1766475.5677341 chr10 52834289 N chr10 52834484 N DEL 23
SRR1766486.11375031 chr10 52835133 N chr10 52835344 N DEL 5
SRR1766482.3501267 chr10 52834343 N chr10 52834494 N DUP 16
SRR1766468.3609739 chr10 52834246 N chr10 52834302 N DUP 25
SRR1766446.9239849 chr10 52834546 N chr10 52835178 N DEL 3
SRR1766473.1894817 chr10 52834617 N chr10 52834964 N DEL 26
SRR1766449.8174668 chr10 52835303 N chr10 52835477 N DEL 10
SRR1766457.8165387 chr10 52834976 N chr10 52835039 N DUP 18
SRR1766475.6106743 chr10 52835035 N chr10 52835450 N DEL 16
SRR1766483.11905056 chr10 52834294 N chr10 52834592 N DEL 5
SRR1766467.1847330 chr10 52834351 N chr10 52834437 N DUP 7
SRR1766471.3025623 chr10 52834265 N chr10 52834466 N DUP 27
SRR1766449.968100 chr10 52834920 N chr10 52835443 N DEL 18
SRR1766445.998017 chr10 52835051 N chr10 52835188 N DEL 4
SRR1766475.897889 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766472.3257059 chr10 52835053 N chr10 52835190 N DEL 2
SRR1766469.4864618 chr10 52834137 N chr10 52834343 N DEL 12
SRR1766467.10368151 chr10 52835238 N chr10 52835344 N DEL 5
SRR1766461.2464575 chr10 52834217 N chr10 52834597 N DEL 5
SRR1766463.6887868 chr10 52834204 N chr10 52834306 N DEL 2
SRR1766456.1725809 chr10 52835133 N chr10 52835344 N DEL 5
SRR1766465.4275800 chr10 52834306 N chr10 52834544 N DEL 22
SRR1766443.10336536 chr10 52834262 N chr10 52834925 N DUP 17
SRR1766450.2855943 chr10 52834663 N chr10 52834923 N DUP 7
SRR1766459.3416325 chr10 52834566 N chr10 52834751 N DEL 11
SRR1766445.3085099 chr10 52834568 N chr10 52834753 N DEL 9
SRR1766473.1894817 chr10 52835273 N chr10 52835344 N DEL 5
SRR1766445.998017 chr10 52834902 N chr10 52834959 N DEL 12
SRR1766461.8929824 chr10 52834328 N chr10 52834861 N DUP 10
SRR1766484.4009 chr10 52835393 N chr10 52835520 N DUP 23
SRR1766469.5343569 chr10 52834295 N chr10 52834602 N DEL 5
SRR1766481.9970168 chr10 52835344 N chr10 52835516 N DUP 10
SRR1766468.5156569 chr10 52834486 N chr10 52834698 N DUP 21
SRR1766446.2610479 chr10 52834119 N chr10 52834895 N DUP 3
SRR1766450.5499935 chr10 52834845 N chr10 52834903 N DEL 10
SRR1766485.1300459 chr10 52834218 N chr10 52835181 N DEL 5
SRR1766446.8358406 chr10 52834297 N chr10 52834906 N DEL 5
SRR1766463.3027132 chr10 52835106 N chr10 52835177 N DEL 1
SRR1766467.824677 chr10 52834481 N chr10 52834553 N DUP 24
SRR1766442.1991002 chr10 52835233 N chr10 52835477 N DEL 14
SRR1766470.10552302 chr10 52834192 N chr10 52834339 N DUP 21
SRR1766486.4689209 chr10 52834961 N chr10 52835471 N DUP 27
SRR1766466.10643060 chr10 52834584 N chr10 52834705 N DEL 27
SRR1766478.11851232 chr10 52834216 N chr10 52834548 N DEL 2
SRR1766477.6829744 chr10 52834231 N chr10 52834896 N DEL 24
SRR1766447.4203927 chr10 52834218 N chr10 52834967 N DEL 9
SRR1766482.7296177 chr10 52834722 N chr10 52834832 N DUP 5
SRR1766481.7605879 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766481.11586842 chr10 52834312 N chr10 52834564 N DEL 6
SRR1766458.64645 chr10 52834295 N chr10 52834593 N DEL 5
SRR1766457.538449 chr10 52834215 N chr10 52834348 N DEL 22
SRR1766470.4965910 chr10 52834920 N chr10 52835443 N DEL 11
SRR1766483.4245322 chr10 52834329 N chr10 52834501 N DEL 22
SRR1766473.4486536 chr10 52834377 N chr10 52834998 N DUP 20
SRR1766469.7981130 chr10 52834159 N chr10 52834344 N DEL 10
SRR1766477.6236954 chr10 52834513 N chr10 52834668 N DUP 16
SRR1766472.4290255 chr10 52834546 N chr10 52835491 N DEL 1
SRR1766461.5280901 chr10 52835100 N chr10 52835484 N DEL 5
SRR1766471.11790596 chr10 52834246 N chr10 52834302 N DUP 25
SRR1766483.8037494 chr10 52834271 N chr10 52834472 N DUP 18
SRR1766476.7922702 chr10 52834262 N chr10 52834452 N DUP 24
SRR1766484.12078672 chr10 52834348 N chr10 52834996 N DUP 21
SRR1766476.4215052 chr10 52835303 N chr10 52835477 N DEL 5
SRR1766451.4203021 chr10 52834348 N chr10 52834444 N DUP 7
SRR1766447.5677813 chr10 52834663 N chr10 52834932 N DUP 17
SRR1766477.9734454 chr10 52834602 N chr10 52835010 N DEL 9
SRR1766447.5252054 chr10 52835303 N chr10 52835477 N DEL 5
SRR1766450.7046305 chr10 52834882 N chr10 52835011 N DUP 25
SRR1766482.2492207 chr10 52834312 N chr10 52834564 N DEL 6
SRR1766470.4965910 chr10 52834546 N chr10 52835011 N DEL 9
SRR1766443.1483430 chr10 52834262 N chr10 52834925 N DUP 14
SRR1766451.4111021 chr10 52834352 N chr10 52834901 N DUP 11
SRR1766482.2991508 chr10 52834307 N chr10 52834538 N DEL 11
SRR1766472.3641776 chr10 52834201 N chr10 52835022 N DUP 8
SRR1766477.45011 chr10 52834568 N chr10 52834753 N DEL 9
SRR1766452.5302509 chr10 52834377 N chr10 52834998 N DUP 20
SRR1766447.9597022 chr10 52834351 N chr10 52834408 N DUP 2
SRR1766459.10529944 chr10 52834299 N chr10 52834675 N DEL 13
SRR1766483.8857063 chr10 52834340 N chr10 52834916 N DEL 2
SRR1766442.34281151 chr10 52835050 N chr10 52835187 N DEL 5
SRR1766460.7474422 chr10 52834265 N chr10 52834466 N DUP 22
SRR1766484.1379780 chr10 52834190 N chr10 52834464 N DUP 12
SRR1766476.9776208 chr10 52834578 N chr10 52834717 N DEL 13
SRR1766472.2495678 chr10 52835012 N chr10 52835442 N DEL 20
SRR1766470.6280216 chr10 52834352 N chr10 52834409 N DUP 9
SRR1766486.8024372 chr10 52834357 N chr10 52834419 N DUP 16
SRR1766451.4429732 chr10 52834165 N chr10 52834302 N DEL 6
SRR1766486.5568017 chr10 52834468 N chr10 52835479 N DEL 14
SRR1766482.7760437 chr10 52834451 N chr10 52835482 N DEL 11
SRR1766473.7015063 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766471.1547623 chr10 52835063 N chr10 52835478 N DEL 5
SRR1766463.10093305 chr10 52834294 N chr10 52834592 N DEL 5
SRR1766455.8223662 chr10 52834663 N chr10 52834932 N DUP 17
SRR1766482.7630141 chr10 52834348 N chr10 52834444 N DUP 7
SRR1766461.4776924 chr10 52834904 N chr10 52834961 N DEL 12
SRR1766449.9944294 chr10 52835238 N chr10 52835344 N DEL 5
SRR1766476.10022101 chr10 52834262 N chr10 52834452 N DUP 23
SRR1766444.6733059 chr10 52835062 N chr10 52835477 N DEL 11
SRR1766475.11081218 chr10 52834282 N chr10 52834479 N DEL 23
SRR1766468.5156569 chr10 52834265 N chr10 52834320 N DUP 8
SRR1766442.37160149 chr10 52835133 N chr10 52835344 N DEL 5
SRR1766471.9964514 chr10 52834138 N chr10 52834205 N DEL 7
SRR1766460.11045787 chr10 52834161 N chr10 52834298 N DEL 7
SRR1766448.6669711 chr10 52834180 N chr10 52834262 N DUP 19
SRR1766476.3496000 chr10 52834228 N chr10 52834360 N DEL 12
SRR1766471.430497 chr10 52834281 N chr10 52834641 N DUP 9
SRR1766475.3720762 chr10 52834217 N chr10 52834899 N DEL 12
SRR1766478.4140472 chr10 52834285 N chr10 52835479 N DEL 3
SRR1766460.37586 chr10 52834606 N chr10 52834886 N DUP 19
SRR1766462.8407781 chr10 52835233 N chr10 52835477 N DEL 14
SRR1766482.7296177 chr10 52834344 N chr10 52834401 N DUP 9
SRR1766470.7228887 chr10 52835238 N chr10 52835344 N DEL 5
SRR1766466.9421547 chr10 52835051 N chr10 52835188 N DEL 4
SRR1766452.1154619 chr10 52834548 N chr10 52834731 N DEL 1
SRR1766452.5180251 chr10 52834527 N chr10 52834878 N DUP 11
SRR1766442.24974403 chr10 52834548 N chr10 52834731 N DEL 1
SRR1766485.2973743 chr10 52834212 N chr10 52834357 N DEL 25
SRR1766482.6922359 chr10 52834547 N chr10 52835354 N DEL 5
SRR1766442.41431891 chr10 52834333 N chr10 52834392 N DUP 15
SRR1766459.4892629 chr10 52834527 N chr10 52834878 N DUP 11
SRR1766471.430497 chr10 52834845 N chr10 52834903 N DEL 24
SRR1766454.3397677 chr10 52834348 N chr10 52834444 N DUP 10
SRR1766465.887054 chr10 52834584 N chr10 52834705 N DEL 27
SRR1766478.6423002 chr10 52834265 N chr10 52834466 N DUP 22
SRR1766457.451781 chr10 52834513 N chr10 52834668 N DUP 15
SRR1766485.2831073 chr10 52834180 N chr10 52834262 N DUP 19
SRR1766442.14654078 chr10 52834159 N chr10 52834344 N DEL 9
SRR1766454.4973854 chr10 52834189 N chr10 52834434 N DUP 7
SRR1766453.3232373 chr10 52835238 N chr10 52835344 N DEL 5
SRR1766450.9493129 chr10 52834213 N chr10 52834296 N DUP 15
SRR1766472.7631750 chr10 52834219 N chr10 52834352 N DEL 11
SRR1766447.7849046 chr10 52834348 N chr10 52834996 N DUP 22
SRR1766467.9335405 chr10 52834963 N chr10 52835230 N DUP 23
SRR1766475.5829802 chr10 52834282 N chr10 52834479 N DEL 18
SRR1766479.744178 chr10 52834299 N chr10 52834675 N DEL 14
SRR1766484.4661740 chr10 52835133 N chr10 52835344 N DEL 5
SRR1766442.14019273 chr10 52834527 N chr10 52834878 N DUP 11
SRR1766484.4009 chr10 52835303 N chr10 52835477 N DEL 5
SRR1766454.4786326 chr10 52834468 N chr10 52835479 N DEL 15
SRR1766452.2901713 chr10 52834349 N chr10 52834406 N DUP 8
SRR1766478.2839191 chr10 52834529 N chr10 52834587 N DEL 14
SRR1766467.11742701 chr10 52834547 N chr10 52835012 N DEL 9
SRR1766461.4203167 chr10 52834888 N chr10 52834982 N DUP 23
SRR1766484.10035188 chr10 52834333 N chr10 52834390 N DUP 5
SRR1766485.1762585 chr10 52834348 N chr10 52834444 N DUP 9
SRR1766442.42273243 chr10 52834343 N chr10 52834400 N DUP 11
SRR1766474.3510913 chr10 52834888 N chr10 52834959 N DEL 8
SRR1766479.5222674 chr10 52834248 N chr10 52834457 N DUP 18
SRR1766469.6471787 chr10 52834156 N chr10 52834623 N DEL 1
SRR1766448.2894725 chr10 52834573 N chr10 52834758 N DEL 11
SRR1766446.10614688 chr10 52834180 N chr10 52834262 N DUP 16
SRR1766450.9493129 chr10 52834136 N chr10 52834342 N DEL 6
SRR1766449.5184961 chr10 52834462 N chr10 52834649 N DEL 17
SRR1766471.10560647 chr10 52835133 N chr10 52835344 N DEL 5
SRR1766477.8918353 chr10 52835062 N chr10 52835477 N DEL 14
SRR1766471.5208502 chr10 52834309 N chr10 52834385 N DUP 14
SRR1766486.11290209 chr10 52834218 N chr10 52835014 N DEL 9
SRR1766472.9945022 chr10 52835133 N chr10 52835344 N DEL 5
SRR1766479.12101956 chr10 52834344 N chr10 52834401 N DUP 7
SRR1766481.10193444 chr10 52835128 N chr10 52835477 N DEL 14
SRR1766453.3279804 chr10 52834663 N chr10 52834932 N DUP 12
SRR1766475.9590094 chr10 52834171 N chr10 52834445 N DUP 16
SRR1766464.9075706 chr10 52834888 N chr10 52834959 N DEL 8
SRR1766483.12347230 chr10 52834548 N chr10 52834999 N DEL 1
SRR1766448.1365620 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766482.5479155 chr10 52834959 N chr10 52835506 N DUP 17
SRR1766468.4270493 chr10 52834196 N chr10 52834313 N DUP 16
SRR1766442.32287062 chr10 52834348 N chr10 52834444 N DUP 5
SRR1766449.3394212 chr10 52834329 N chr10 52834501 N DEL 10
SRR1766454.8238494 chr10 52834214 N chr10 52834333 N DEL 14
SRR1766452.7871041 chr10 52834592 N chr10 52834953 N DUP 22
SRR1766478.2839191 chr10 52834223 N chr10 52834988 N DEL 5
SRR1766447.9225541 chr10 52834348 N chr10 52834444 N DUP 20
SRR1766464.10330159 chr10 52834600 N chr10 52834917 N DEL 1
SRR1766465.5664335 chr10 52835303 N chr10 52835477 N DEL 5
SRR1766442.28290693 chr10 52834974 N chr10 52835037 N DUP 20
SRR1766466.7311472 chr10 52834191 N chr10 52834386 N DUP 7
SRR1766458.2707345 chr10 52834309 N chr10 52834433 N DUP 10
SRR1766464.9075706 chr10 52834162 N chr10 52834347 N DEL 6
SRR1766453.10178649 chr10 52835303 N chr10 52835477 N DEL 8
SRR1766483.3848811 chr10 52834959 N chr10 52835506 N DUP 15
SRR1766452.2697857 chr10 52834348 N chr10 52834444 N DUP 8
SRR1766443.2792696 chr10 52834212 N chr10 52834357 N DEL 24
SRR1766442.32442699 chr10 52835099 N chr10 52835483 N DEL 5
SRR1766443.817493 chr10 52835063 N chr10 52835478 N DEL 5
SRR1766452.7240253 chr10 52834573 N chr10 52834758 N DEL 9
SRR1766465.4606849 chr10 52834312 N chr10 52834564 N DEL 6
SRR1766458.2193736 chr10 52835303 N chr10 52835477 N DEL 7
SRR1766448.5502724 chr10 52834468 N chr10 52835479 N DEL 14
SRR1766483.4662958 chr10 52834235 N chr10 52834755 N DEL 13
SRR1766448.6012014 chr10 52835316 N chr10 52835500 N DEL 14
SRR1766464.6711284 chr10 52834300 N chr10 52834541 N DEL 20
SRR1766457.6722196 chr10 52834215 N chr10 52834348 N DEL 15
SRR1766467.961717 chr10 52834208 N chr10 52834341 N DEL 17
SRR1766473.3750949 chr10 52834246 N chr10 52834302 N DUP 15
SRR1766470.2999087 chr10 52834262 N chr10 52834423 N DUP 13
SRR1766460.6127982 chr10 52834132 N chr10 52834492 N DEL 3
SRR1766444.3871796 chr10 52835062 N chr10 52835477 N DEL 6
SRR1766468.4012834 chr10 52834584 N chr10 52834705 N DEL 22
SRR1766448.10886233 chr10 52835128 N chr10 52835477 N DEL 14
SRR1766453.10706545 chr10 52834571 N chr10 52835182 N DEL 5
SRR1766462.8407781 chr10 52834272 N chr10 52835317 N DUP 12
SRR1766464.1752034 chr10 52835238 N chr10 52835344 N DEL 5
SRR1766459.4380243 chr10 52834526 N chr10 52834663 N DUP 17
SRR1766456.1725809 chr10 52834966 N chr10 52835029 N DUP 29
SRR1766464.6430532 chr10 52834343 N chr10 52834494 N DUP 12
SRR1766482.12101491 chr10 52835303 N chr10 52835477 N DEL 5
SRR1766446.2319339 chr10 52834845 N chr10 52834903 N DEL 23
SRR1766442.14654078 chr10 52834343 N chr10 52834494 N DUP 15
SRR1766459.11359956 chr10 52834348 N chr10 52834444 N DUP 15
SRR1766444.2642762 chr10 52834234 N chr10 52834348 N DEL 7
SRR1766459.141569 chr10 52834985 N chr10 52835480 N DEL 11
SRR1766442.27176991 chr10 52834399 N chr10 52834662 N DEL 19
SRR1766483.2483593 chr10 52834171 N chr10 52834689 N DUP 29
SRR1766442.14728366 chr10 52834344 N chr10 52834401 N DUP 9
SRR1766447.10406924 chr10 52834348 N chr10 52834444 N DUP 8
SRR1766442.18310656 chr10 52834374 N chr10 52834538 N DEL 16
SRR1766461.2464575 chr10 52834192 N chr10 52834318 N DUP 26
SRR1766442.39697121 chr10 52835103 N chr10 52835487 N DEL 5
SRR1766480.2943060 chr10 52835273 N chr10 52835344 N DEL 5
SRR1766482.5595008 chr10 52835103 N chr10 52835349 N DEL 5
SRR1766461.2952880 chr10 52834592 N chr10 52834669 N DUP 14
SRR1766458.5578702 chr10 52834215 N chr10 52834348 N DEL 15
SRR1766455.5570219 chr10 52834294 N chr10 52834592 N DEL 5
SRR1766469.4913358 chr10 52834302 N chr10 52834512 N DEL 15
SRR1766482.3501267 chr10 52834364 N chr10 52834435 N DEL 16
SRR1766469.4130133 chr10 52834606 N chr10 52834886 N DUP 18
SRR1766467.7400907 chr10 52834239 N chr10 52834290 N DEL 8
SRR1766465.9287042 chr10 52834283 N chr10 52834643 N DUP 9
SRR1766469.8460650 chr10 52835047 N chr10 52835184 N DEL 5
SRR1766474.10669696 chr10 52834546 N chr10 52835178 N DEL 3
SRR1766476.5757096 chr10 52835268 N chr10 52835477 N DEL 14
SRR1766459.4207964 chr10 52835133 N chr10 52835344 N DEL 5
SRR1766454.11115193 chr10 52835238 N chr10 52835344 N DEL 5
SRR1766465.8571054 chr10 52834287 N chr10 52834636 N DUP 16
SRR1766484.3548182 chr10 52834592 N chr10 52834953 N DUP 22
SRR1766442.6349846 chr10 52834211 N chr10 52834528 N DUP 11
SRR1766453.2168285 chr10 52834882 N chr10 52835011 N DUP 27
SRR1766459.4207964 chr10 52834222 N chr10 52834896 N DEL 15
SRR1766464.46233 chr10 52834566 N chr10 52834751 N DEL 11
SRR1766448.5519213 chr10 52834307 N chr10 52834538 N DEL 10
SRR1766454.1715984 chr7 152487421 N chr7 152487490 N DEL 11
SRR1766475.10384997 chr11 1914629 N chr11 1914739 N DUP 3
SRR1766479.6186913 chr11 1914747 N chr11 1914874 N DEL 5
SRR1766466.4098909 chr11 1914644 N chr11 1914700 N DEL 2
SRR1766475.10981755 chr11 1914585 N chr11 1914871 N DUP 5
SRR1766482.4827801 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766480.2623144 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766480.818389 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766454.7846305 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766446.7630853 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766483.4936861 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766442.2172999 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766464.2079031 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766479.12690752 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766443.4502369 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766479.9858863 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766454.9243505 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766449.7264974 chr18 1747175 N chr18 1747232 N DEL 5
SRR1766461.8160401 chr18 1747179 N chr18 1747240 N DUP 20
SRR1766455.7967884 chr18 1747201 N chr18 1747262 N DUP 15
SRR1766482.5069586 chr18 1747189 N chr18 1747282 N DUP 19
SRR1766470.774084 chr18 1747179 N chr18 1747252 N DUP 18
SRR1766464.8511475 chr18 1747181 N chr18 1747280 N DUP 17
SRR1766485.11357864 chr18 1747179 N chr18 1747270 N DUP 14
SRR1766445.673797 chr18 1747233 N chr18 1747296 N DUP 4
SRR1766464.8756450 chr18 1747223 N chr18 1747310 N DUP 12
SRR1766453.1027038 chr18 1747206 N chr18 1747323 N DEL 13
SRR1766453.7278841 chr18 1747210 N chr18 1747327 N DEL 9
SRR1766452.2782993 chr18 1747219 N chr18 1747402 N DEL 18
SRR1766467.9813751 chr7 20278120 N chr7 20278203 N DEL 6
SRR1766467.2550308 chr5 38832207 N chr5 38832338 N DEL 12
SRR1766470.4484859 chr5 38832209 N chr5 38832338 N DEL 13
SRR1766481.9098975 chr5 38832231 N chr5 38832326 N DUP 1
SRR1766474.7799439 chr5 38832255 N chr5 38832348 N DUP 12
SRR1766456.508299 chr5 38832212 N chr5 38832289 N DEL 10
SRR1766451.1863865 chr5 38832210 N chr5 38832313 N DEL 6
SRR1766459.5551605 chr5 38832251 N chr5 38832338 N DEL 20
SRR1766457.5919399 chr5 38832251 N chr5 38832338 N DEL 12
SRR1766475.6073013 chr5 38832210 N chr5 38832347 N DEL 6
SRR1766464.10940282 chr5 38832210 N chr5 38832347 N DEL 6
SRR1766472.6618929 chr17 83120066 N chr17 83120165 N DEL 12
SRR1766452.9628770 chr17 83120204 N chr17 83120258 N DEL 25
SRR1766451.6950533 chr17 83120081 N chr17 83120266 N DEL 6
SRR1766449.3155568 chr3 50076518 N chr3 50076824 N DEL 26
SRR1766477.8242704 chr5 174982971 N chr5 174983086 N DUP 4
SRR1766480.2808339 chr10 6413623 N chr10 6413738 N DEL 22
SRR1766442.12402026 chr10 6413688 N chr10 6413832 N DEL 14
SRR1766469.7269358 chr10 6413688 N chr10 6413832 N DEL 15
SRR1766481.6314684 chr10 6413628 N chr10 6413686 N DUP 21
SRR1766471.10342797 chr10 6413627 N chr10 6413787 N DEL 33
SRR1766485.5284021 chr10 6413627 N chr10 6413787 N DEL 35
SRR1766477.3440084 chr10 6413686 N chr10 6413883 N DEL 12
SRR1766486.2323722 chr10 6413700 N chr10 6413787 N DEL 30
SRR1766452.10099801 chr10 6413796 N chr10 6413889 N DUP 5
SRR1766442.36883666 chr10 6413631 N chr10 6413791 N DEL 11
SRR1766456.1229338 chr10 6413633 N chr10 6413793 N DEL 9
SRR1766471.9762153 chr10 6413634 N chr10 6413794 N DEL 8
SRR1766442.44511183 chr10 6413635 N chr10 6413795 N DEL 1
SRR1766479.7530171 chr10 6413786 N chr10 6413838 N DUP 13
SRR1766474.9353504 chr10 6413686 N chr10 6413883 N DEL 12
SRR1766484.4952826 chr10 6413786 N chr10 6413881 N DUP 13
SRR1766446.8155806 chr10 6413789 N chr10 6413925 N DUP 13
SRR1766462.7981236 chr10 6413786 N chr10 6413881 N DUP 14
SRR1766447.3135905 chr10 6413687 N chr10 6413884 N DEL 13
SRR1766451.6067218 chr10 6413688 N chr10 6413885 N DEL 13
SRR1766442.20028075 chr10 6413693 N chr10 6413890 N DEL 8
SRR1766482.8213441 chr10 6413690 N chr10 6413887 N DEL 11
SRR1766469.8753172 chr6 164021962 N chr6 164022033 N DEL 1
SRR1766461.604290 chr6 160855432 N chr6 160855523 N DUP 5
SRR1766466.4873651 chr7 118266726 N chr7 118266920 N DUP 5
SRR1766475.4991623 chr7 118266685 N chr7 118266851 N DUP 7
SRR1766471.11386848 chr7 118266685 N chr7 118266851 N DUP 7
SRR1766442.24365806 chr7 118266685 N chr7 118266851 N DUP 7
SRR1766473.3152290 chr7 118266685 N chr7 118266851 N DUP 7
SRR1766473.2814108 chr7 118266685 N chr7 118266851 N DUP 7
SRR1766453.10492959 chr7 118266685 N chr7 118266851 N DUP 7
SRR1766484.1433841 chr7 118266685 N chr7 118266851 N DUP 7
SRR1766460.2331825 chr7 118266708 N chr7 118266852 N DEL 5
SRR1766472.3474390 chr7 118266708 N chr7 118266852 N DEL 9
SRR1766479.11587849 chr7 112391504 N chr7 112391791 N DEL 3
SRR1766486.1490529 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766474.8047790 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766462.8765076 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766452.4460274 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766479.6029697 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766455.8401804 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766476.9245016 chr7 112391550 N chr7 112391785 N DEL 10
SRR1766442.43306086 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766453.6178582 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766454.5842177 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766464.4237874 chr7 112391497 N chr7 112391574 N DUP 7
SRR1766467.10254535 chr7 112391530 N chr7 112391739 N DEL 5
SRR1766467.5651111 chr7 112391504 N chr7 112391791 N DEL 5
SRR1766442.24644621 chr7 112391530 N chr7 112392025 N DEL 10
SRR1766453.2580210 chr7 112391508 N chr7 112391795 N DEL 5
SRR1766477.5170727 chr7 112391509 N chr7 112391796 N DEL 5
SRR1766478.8757906 chr7 112391514 N chr7 112391801 N DEL 5
SRR1766448.9221969 chr7 112391497 N chr7 112391626 N DUP 3
SRR1766442.20469549 chr7 112391702 N chr7 112391989 N DEL 5
SRR1766483.8993707 chr7 112391702 N chr7 112391989 N DEL 5
SRR1766458.409043 chr7 112391517 N chr7 112391804 N DEL 2
SRR1766475.9956056 chr7 112391518 N chr7 112391805 N DEL 1
SRR1766447.1853055 chr7 112391495 N chr7 112391808 N DEL 2
SRR1766476.6868882 chr7 112391619 N chr7 112391802 N DEL 5
SRR1766475.5599785 chr7 112391805 N chr7 112391908 N DUP 5
SRR1766442.36512405 chr7 112391805 N chr7 112391908 N DUP 5
SRR1766458.5069920 chr7 112391805 N chr7 112391908 N DUP 5
SRR1766483.12466808 chr7 112391805 N chr7 112391908 N DUP 5
SRR1766478.4536212 chr7 112391805 N chr7 112391908 N DUP 5
SRR1766483.5940038 chr7 112391805 N chr7 112391908 N DUP 5
SRR1766467.7658214 chr7 112391805 N chr7 112391908 N DUP 5
SRR1766451.6861621 chr7 112391805 N chr7 112391908 N DUP 5
SRR1766442.36191933 chr7 112391622 N chr7 112391805 N DEL 5
SRR1766458.6181297 chr7 112391622 N chr7 112391805 N DEL 5
SRR1766464.1976 chr7 112391622 N chr7 112391805 N DEL 5
SRR1766479.13049005 chr7 112391622 N chr7 112391805 N DEL 5
SRR1766474.1414707 chr7 112391668 N chr7 112392059 N DEL 10
SRR1766450.5205204 chr7 112391690 N chr7 112392107 N DEL 5
SRR1766451.1415670 chr7 112391622 N chr7 112391805 N DEL 5
SRR1766455.6918568 chr7 112391622 N chr7 112391805 N DEL 5
SRR1766486.2296179 chr7 112392027 N chr7 112392106 N DEL 7
SRR1766449.9305565 chr7 112391626 N chr7 112392017 N DEL 5
SRR1766486.5617474 chr7 112391702 N chr7 112391989 N DEL 5
SRR1766477.3642909 chr7 112391612 N chr7 112391819 N DUP 15
SRR1766461.8546996 chr7 112391708 N chr7 112391995 N DEL 5
SRR1766463.1863768 chr7 112391715 N chr7 112392002 N DEL 2
SRR1766462.3231539 chr7 112391509 N chr7 112392106 N DUP 2
SRR1766479.10868894 chr7 112391819 N chr7 112392106 N DEL 5
SRR1766442.2713876 chr7 112391473 N chr7 112392096 N DUP 8
SRR1766485.11629303 chr7 112391509 N chr7 112392106 N DUP 5
SRR1766480.4986645 chr7 112391795 N chr7 112392106 N DUP 5
SRR1766447.4304736 chr7 112391795 N chr7 112392106 N DUP 5
SRR1766478.4207645 chr7 112391795 N chr7 112392106 N DUP 5
SRR1766480.3140755 chr7 112391795 N chr7 112391898 N DUP 5
SRR1766446.498063 chr7 112391795 N chr7 112391898 N DUP 5
SRR1766468.5296447 chr7 112391795 N chr7 112391898 N DUP 5
SRR1766458.9197167 chr7 112391795 N chr7 112391898 N DUP 5
SRR1766458.2803713 chr7 112391795 N chr7 112391898 N DUP 5
SRR1766466.10706763 chr7 112391795 N chr7 112391898 N DUP 5
SRR1766457.6661971 chr7 112391499 N chr7 112392174 N DUP 1
SRR1766464.6474469 chr7 112391802 N chr7 112391905 N DUP 5
SRR1766465.9231362 chr7 112391482 N chr7 112392183 N DUP 8
SRR1766445.2534350 chr7 112391612 N chr7 112391795 N DEL 5
SRR1766474.5711040 chr7 112391612 N chr7 112391795 N DEL 5
SRR1766471.11482953 chr7 112391612 N chr7 112391795 N DEL 5
SRR1766475.8434690 chr7 112391617 N chr7 112391800 N DEL 5
SRR1766476.61887 chr7 112391617 N chr7 112391800 N DEL 5
SRR1766472.5536930 chr7 112391659 N chr7 112392258 N DEL 15
SRR1766475.8434690 chr7 112392116 N chr7 112392221 N DEL 5
SRR1766443.9825298 chr7 112391885 N chr7 112392302 N DEL 65
SRR1766454.6572817 chr7 43247894 N chr7 43248057 N DEL 7
SRR1766443.9655547 chr7 43247894 N chr7 43248057 N DEL 7
SRR1766474.11235264 chr7 43247841 N chr7 43248226 N DEL 1
SRR1766443.8510253 chrX 2446459 N chrX 2446947 N DEL 15
SRR1766474.2665763 chrX 2446500 N chrX 2446700 N DUP 5
SRR1766442.1086178 chrX 2446616 N chrX 2446715 N DUP 5
SRR1766484.4524200 chrX 2446432 N chrX 2446672 N DEL 11
SRR1766474.10561355 chrX 2446520 N chrX 2446819 N DUP 1
SRR1766446.284581 chrX 2446630 N chrX 2446828 N DUP 5
SRR1766458.4128312 chrX 2446430 N chrX 2446819 N DEL 5
SRR1766453.4164470 chrX 2446750 N chrX 2446947 N DUP 5
SRR1766456.4498277 chr2 1679234 N chr2 1679428 N DUP 1
SRR1766467.69689 chr16 3062313 N chr16 3063042 N DEL 4
SRR1766482.11538486 chr16 3062313 N chr16 3063042 N DEL 5
SRR1766482.9235664 chr16 3062346 N chr16 3063073 N DUP 5
SRR1766457.4766476 chr16 3062346 N chr16 3063073 N DUP 5
SRR1766472.262120 chr16 3062346 N chr16 3063073 N DUP 5
SRR1766484.3885919 chr16 3062350 N chr16 3063077 N DUP 5
SRR1766472.3644320 chr16 3062519 N chr16 3063241 N DUP 5
SRR1766474.5856253 chr16 3062628 N chr16 3063352 N DEL 10
SRR1766449.148659 chr16 3062774 N chr16 3063498 N DEL 17
SRR1766460.9155194 chr8 7107227 N chr8 7107284 N DEL 1
SRR1766445.4839265 chr5 62514053 N chr5 62514326 N DEL 5
SRR1766484.5375214 chr5 62514078 N chr5 62514272 N DEL 5
SRR1766442.32707040 chr5 62513951 N chr5 62514185 N DEL 2
SRR1766450.10657166 chr13 41102760 N chr13 41103076 N DUP 2
SRR1766481.11161675 chr13 41102939 N chr13 41102997 N DEL 5
SRR1766453.2487347 chr9 64773276 N chr9 64773393 N DEL 10
SRR1766463.6339014 chr9 64773482 N chr9 64773754 N DUP 11
SRR1766443.3992319 chr17 41051507 N chr17 41051560 N DUP 7
SRR1766481.3218934 chr2 70149051 N chr2 70149171 N DEL 12
SRR1766470.1387572 chr2 70148977 N chr2 70149214 N DUP 5
SRR1766482.6596411 chr17 46227294 N chr17 46227430 N DUP 3
SRR1766453.7920040 chr17 46227294 N chr17 46227430 N DUP 4
SRR1766443.10182651 chr3 195710912 N chr3 195711138 N DEL 10
SRR1766442.41509030 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766445.9976419 chr3 195710745 N chr3 195710881 N DEL 23
SRR1766455.5079765 chr3 195710833 N chr3 195711237 N DUP 10
SRR1766474.8942288 chr3 195710873 N chr3 195710962 N DUP 1
SRR1766473.3015078 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766460.3349304 chr3 195710639 N chr3 195711178 N DUP 5
SRR1766442.44332938 chr3 195710427 N chr3 195711191 N DUP 1
SRR1766486.10732033 chr3 195710880 N chr3 195710971 N DEL 10
SRR1766476.6415116 chr3 195710507 N chr3 195711453 N DEL 5
SRR1766483.1831430 chr3 195710663 N chr3 195711159 N DEL 4
SRR1766473.9842351 chr3 195710658 N chr3 195710884 N DEL 5
SRR1766446.5311731 chr3 195710507 N chr3 195711453 N DEL 5
SRR1766450.10621828 chr3 195710594 N chr3 195710773 N DUP 10
SRR1766476.639670 chr3 195710926 N chr3 195711195 N DUP 5
SRR1766479.8268678 chr3 195710782 N chr3 195711413 N DEL 7
SRR1766457.3462539 chr3 195710507 N chr3 195711574 N DEL 15
SRR1766474.8942288 chr3 195710672 N chr3 195711168 N DEL 18
SRR1766445.5508784 chr3 195710655 N chr3 195710926 N DEL 5
SRR1766445.7215442 chr3 195710475 N chr3 195711106 N DEL 5
SRR1766442.30048324 chr3 195710777 N chr3 195711138 N DEL 20
SRR1766475.5597405 chr3 195710910 N chr3 195711572 N DEL 15
SRR1766448.9376852 chr3 195711152 N chr3 195711376 N DUP 10
SRR1766442.21389072 chr3 195710647 N chr3 195711098 N DEL 9
SRR1766460.6671650 chr3 195710687 N chr3 195710913 N DEL 5
SRR1766448.5636186 chr3 195710517 N chr3 195710878 N DEL 5
SRR1766485.1377181 chr3 195710507 N chr3 195711453 N DEL 5
SRR1766455.9004478 chr3 195710727 N chr3 195711133 N DEL 10
SRR1766474.1491531 chr3 195710912 N chr3 195711138 N DEL 10
SRR1766442.19902109 chr3 195710637 N chr3 195711221 N DUP 20
SRR1766460.4964616 chr3 195710427 N chr3 195710516 N DUP 10
SRR1766474.4518123 chr3 195711087 N chr3 195711268 N DEL 5
SRR1766474.9856445 chr3 195711182 N chr3 195711453 N DEL 22
SRR1766451.2486518 chr3 195710672 N chr3 195711123 N DEL 5
SRR1766460.8032200 chr3 195710855 N chr3 195711034 N DUP 8
SRR1766468.3988988 chr3 195710457 N chr3 195711133 N DEL 5
SRR1766484.9848909 chr3 195711168 N chr3 195711347 N DUP 10
SRR1766449.5724436 chr3 195710912 N chr3 195711273 N DEL 15
SRR1766483.4753288 chr3 195710745 N chr3 195710881 N DEL 10
SRR1766442.29532329 chr3 195710465 N chr3 195711141 N DEL 4
SRR1766454.7061863 chr3 195710857 N chr3 195711351 N DUP 6
SRR1766442.19981783 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766476.5840858 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766467.4323641 chr3 195710427 N chr3 195710921 N DUP 9
SRR1766477.10566214 chr3 195710833 N chr3 195711327 N DUP 10
SRR1766465.5826697 chr3 195710594 N chr3 195711223 N DUP 10
SRR1766469.3467702 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766478.4854940 chr3 195710547 N chr3 195711614 N DEL 5
SRR1766447.7067491 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766453.2806591 chr3 195710745 N chr3 195710836 N DEL 20
SRR1766442.36643126 chr3 195710521 N chr3 195711152 N DEL 1
SRR1766455.5079765 chr3 195710475 N chr3 195711286 N DEL 10
SRR1766479.754355 chr3 195710645 N chr3 195711096 N DEL 7
SRR1766467.10289914 chr3 195710700 N chr3 195710836 N DEL 18
SRR1766464.3323994 chr3 195710655 N chr3 195710926 N DEL 5
SRR1766452.6045983 chr3 195710745 N chr3 195711106 N DEL 15
SRR1766476.6169700 chr3 195710837 N chr3 195711151 N DUP 5
SRR1766442.20460302 chr3 195710746 N chr3 195711330 N DUP 10
SRR1766459.1023357 chr3 195710428 N chr3 195710652 N DUP 5
SRR1766478.6919910 chr3 195710704 N chr3 195710840 N DEL 10
SRR1766481.12050387 chr3 195710833 N chr3 195711237 N DUP 8
SRR1766476.5840858 chr3 195711103 N chr3 195711372 N DUP 15
SRR1766442.16760103 chr3 195710653 N chr3 195710967 N DUP 10
SRR1766459.2602484 chr3 195710475 N chr3 195711151 N DEL 5
SRR1766486.4866519 chr3 195711242 N chr3 195711333 N DEL 5
SRR1766473.1854743 chr3 195711012 N chr3 195711148 N DEL 15
SRR1766473.10023160 chr3 195711012 N chr3 195711148 N DEL 5
SRR1766457.9207961 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766481.401328 chr3 195710880 N chr3 195710971 N DEL 10
SRR1766460.5415474 chr3 195710745 N chr3 195710836 N DEL 25
SRR1766469.3986800 chr3 195710925 N chr3 195711331 N DEL 10
SRR1766450.9305504 chr3 195710913 N chr3 195711227 N DUP 10
SRR1766442.15852406 chr3 195710745 N chr3 195711061 N DEL 5
SRR1766460.1511398 chr3 195710789 N chr3 195711373 N DUP 20
SRR1766474.8532251 chr3 195710970 N chr3 195711151 N DEL 15
SRR1766451.5868940 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766472.4780329 chr3 195710912 N chr3 195711093 N DEL 10
SRR1766484.6714236 chr3 195711182 N chr3 195711273 N DEL 1
SRR1766476.11238745 chr3 195710676 N chr3 195711217 N DEL 5
SRR1766442.12486994 chr3 195710672 N chr3 195711213 N DEL 10
SRR1766476.6082131 chr3 195710732 N chr3 195711273 N DEL 10
SRR1766442.11963976 chr3 195710509 N chr3 195711050 N DEL 1
SRR1766459.9666726 chr3 195710732 N chr3 195711273 N DEL 10
SRR1766448.6660259 chr3 195710464 N chr3 195711140 N DEL 5
SRR1766442.17853161 chr3 195710512 N chr3 195711233 N DEL 5
SRR1766470.8672911 chr3 195710656 N chr3 195710745 N DUP 13
SRR1766442.29153075 chr3 195710826 N chr3 195711412 N DEL 5
SRR1766478.8736120 chr3 195710633 N chr3 195711262 N DUP 12
SRR1766474.7567723 chr3 195711103 N chr3 195711372 N DUP 15
SRR1766444.3503240 chr3 195710722 N chr3 195711308 N DEL 19
SRR1766442.293454 chr3 195710732 N chr3 195711228 N DEL 5
SRR1766471.9995658 chr3 195710830 N chr3 195711146 N DEL 5
SRR1766468.6713900 chr3 195710686 N chr3 195711092 N DEL 1
SRR1766454.2024097 chr3 195710836 N chr3 195710925 N DUP 12
SRR1766465.553161 chr3 195710970 N chr3 195711106 N DEL 10
SRR1766448.8109133 chr3 195710618 N chr3 195710979 N DEL 5
SRR1766450.394408 chr3 195710638 N chr3 195711177 N DUP 10
SRR1766453.5877578 chr3 195710573 N chr3 195710799 N DEL 23
SRR1766473.10829557 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766470.1634696 chr3 195711143 N chr3 195711232 N DUP 9
SRR1766477.7248460 chr3 195710426 N chr3 195711057 N DEL 10
SRR1766451.5719409 chr3 195710507 N chr3 195711453 N DEL 5
SRR1766454.8857819 chr3 195710426 N chr3 195711057 N DEL 5
SRR1766484.6714236 chr3 195710547 N chr3 195711614 N DEL 5
SRR1766466.6654618 chr3 195711013 N chr3 195711192 N DUP 11
SRR1766479.12475779 chr3 195711088 N chr3 195711357 N DUP 10
SRR1766447.5846248 chr3 195710833 N chr3 195710967 N DUP 11
SRR1766443.4776958 chr3 195710881 N chr3 195711541 N DUP 3
SRR1766485.5620443 chr3 195710745 N chr3 195710836 N DEL 12
SRR1766477.2032102 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766462.7946574 chr3 195711182 N chr3 195711273 N DEL 10
SRR1766474.7022316 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766485.5033270 chr3 195710970 N chr3 195711331 N DEL 5
SRR1766445.4460209 chr3 195711182 N chr3 195711273 N DEL 2
SRR1766443.4603466 chr3 195710970 N chr3 195711061 N DEL 10
SRR1766455.9004478 chr3 195710427 N chr3 195710741 N DUP 10
SRR1766466.1081679 chr3 195710745 N chr3 195711286 N DEL 19
SRR1766470.8820644 chr3 195710913 N chr3 195711227 N DUP 5
SRR1766449.8071792 chr3 195710812 N chr3 195711083 N DEL 4
SRR1766477.8888269 chr3 195710547 N chr3 195711614 N DEL 5
SRR1766454.10630146 chr3 195710778 N chr3 195711409 N DEL 21
SRR1766485.7085306 chr3 195710514 N chr3 195711100 N DEL 5
SRR1766477.10568729 chr3 195710550 N chr3 195711091 N DEL 5
SRR1766442.31880571 chr3 195710871 N chr3 195711185 N DUP 2
SRR1766463.7189814 chr3 195710777 N chr3 195711093 N DEL 10
SRR1766474.532605 chr3 195710913 N chr3 195711227 N DUP 10
SRR1766466.9588803 chr3 195710853 N chr3 195711212 N DUP 5
SRR1766477.5874484 chr3 195710660 N chr3 195710974 N DUP 4
SRR1766479.8854023 chr3 195710878 N chr3 195711372 N DUP 17
SRR1766480.7071623 chr3 195710549 N chr3 195711571 N DEL 5
SRR1766463.8865853 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766477.6908917 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766476.7856287 chr3 195710639 N chr3 195711133 N DUP 10
SRR1766455.3351269 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766443.6487521 chr3 195710673 N chr3 195711032 N DUP 5
SRR1766457.8737280 chr3 195710628 N chr3 195711347 N DUP 4
SRR1766468.5751723 chr3 195710628 N chr3 195710897 N DUP 10
SRR1766481.13112492 chr3 195710970 N chr3 195711331 N DEL 5
SRR1766449.6616360 chr3 195710833 N chr3 195711192 N DUP 14
SRR1766482.12935902 chr3 195710781 N chr3 195711277 N DEL 8
SRR1766464.9617415 chr3 195710687 N chr3 195710913 N DEL 5
SRR1766450.887153 chr3 195711148 N chr3 195711372 N DUP 11
SRR1766447.408951 chr3 195710926 N chr3 195711375 N DUP 15
SRR1766449.6367427 chr3 195710732 N chr3 195711273 N DEL 10
SRR1766465.10858498 chr3 195710507 N chr3 195711093 N DEL 3
SRR1766442.1312105 chr3 195710713 N chr3 195710849 N DEL 2
SRR1766447.2783696 chr3 195710457 N chr3 195711133 N DEL 5
SRR1766467.6525917 chr3 195710976 N chr3 195711337 N DEL 5
SRR1766461.5477121 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766443.4420589 chr3 195710431 N chr3 195711105 N DUP 5
SRR1766459.7609795 chr3 195710777 N chr3 195711093 N DEL 10
SRR1766448.6428267 chr3 195710507 N chr3 195710868 N DEL 3
SRR1766466.5167720 chr3 195711452 N chr3 195711619 N DEL 7
SRR1766466.3648164 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766459.9666726 chr3 195710687 N chr3 195710913 N DEL 5
SRR1766474.606011 chr3 195711087 N chr3 195711268 N DEL 7
SRR1766483.75109 chr3 195710913 N chr3 195711227 N DUP 10
SRR1766482.9329879 chr3 195710665 N chr3 195711161 N DEL 2
SRR1766466.5914983 chr3 195710475 N chr3 195711286 N DEL 10
SRR1766457.8172859 chr3 195711229 N chr3 195711363 N DUP 10
SRR1766485.5308376 chr3 195711239 N chr3 195711330 N DEL 5
SRR1766475.336802 chr3 195710459 N chr3 195711270 N DEL 5
SRR1766486.3483938 chr3 195710913 N chr3 195711227 N DUP 10
SRR1766468.5959020 chr3 195710923 N chr3 195711104 N DEL 10
SRR1766477.1346454 chr3 195710700 N chr3 195710836 N DEL 20
SRR1766464.3221854 chr3 195711078 N chr3 195711347 N DUP 10
SRR1766479.2256567 chr3 195710652 N chr3 195711283 N DEL 15
SRR1766476.5257357 chr3 195710626 N chr3 195711345 N DUP 9
SRR1766479.12792430 chr3 195710781 N chr3 195711578 N DEL 25
SRR1766443.10088010 chr3 195711267 N chr3 195711614 N DEL 8
SRR1766480.7694544 chr3 195710745 N chr3 195710836 N DEL 10
SRR1766465.8842441 chr3 195710459 N chr3 195711405 N DEL 19
SRR1766466.7668531 chr3 195711147 N chr3 195711371 N DUP 5
SRR1766481.5904257 chr3 195710723 N chr3 195711172 N DUP 6
SRR1766467.10289914 chr3 195710862 N chr3 195711268 N DEL 15
SRR1766445.10054146 chr3 195710789 N chr3 195711283 N DUP 9
SRR1766484.8928592 chr3 195710789 N chr3 195711373 N DUP 10
SRR1766450.7082925 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766482.13286804 chr3 195711147 N chr3 195711371 N DUP 5
SRR1766476.2866907 chr3 195710656 N chr3 195710745 N DUP 11
SRR1766481.5149619 chr3 195710644 N chr3 195711005 N DEL 5
SRR1766448.837598 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766465.553161 chr3 195711140 N chr3 195711319 N DUP 10
SRR1766445.9596139 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766471.169227 chr3 195710868 N chr3 195711182 N DUP 12
SRR1766480.7559984 chr3 195710457 N chr3 195711133 N DEL 10
SRR1766458.189902 chr3 195710727 N chr3 195711133 N DEL 10
SRR1766483.10796568 chr3 195710475 N chr3 195711151 N DEL 10
SRR1766452.5175672 chr3 195710464 N chr3 195711140 N DEL 5
SRR1766486.8021375 chr3 195710441 N chr3 195710802 N DEL 2
SRR1766464.8428911 chr3 195710547 N chr3 195710863 N DEL 15
SRR1766474.4221618 chr3 195710428 N chr3 195710652 N DUP 5
SRR1766464.8428911 chr3 195710745 N chr3 195710836 N DEL 23
SRR1766460.8663933 chr3 195710911 N chr3 195711137 N DEL 15
SRR1766468.6262396 chr3 195710475 N chr3 195711061 N DEL 14
SRR1766445.6058925 chr3 195710574 N chr3 195711293 N DUP 2
SRR1766460.6925891 chr3 195711078 N chr3 195711347 N DUP 10
SRR1766452.10612767 chr3 195710877 N chr3 195711011 N DUP 1
SRR1766459.2913378 chr3 195710661 N chr3 195711067 N DEL 5
SRR1766463.8588399 chr3 195710898 N chr3 195711032 N DUP 10
SRR1766442.14751536 chr3 195710547 N chr3 195710863 N DEL 15
SRR1766460.10106805 chr3 195710789 N chr3 195711148 N DUP 17
SRR1766476.2578643 chr3 195710511 N chr3 195710872 N DEL 5
SRR1766455.8059299 chr3 195710478 N chr3 195711154 N DEL 5
SRR1766445.4101327 chr3 195710672 N chr3 195711123 N DEL 5
SRR1766478.3047540 chr3 195710992 N chr3 195711128 N DEL 4
SRR1766442.37821852 chr3 195710673 N chr3 195711032 N DUP 5
SRR1766449.2039271 chr3 195710833 N chr3 195710922 N DUP 20
SRR1766459.6172648 chr3 195710656 N chr3 195710745 N DUP 20
SRR1766473.3028541 chr3 195711012 N chr3 195711148 N DEL 5
SRR1766450.1336038 chr3 195710745 N chr3 195711286 N DEL 10
SRR1766482.10001994 chr3 195710878 N chr3 195711372 N DUP 10
SRR1766455.2201857 chr3 195711012 N chr3 195711148 N DEL 15
SRR1766485.984262 chr3 195710732 N chr3 195711138 N DEL 10
SRR1766463.7304346 chr3 195710633 N chr3 195711217 N DUP 10
SRR1766449.8188394 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766465.10858498 chr3 195710712 N chr3 195711073 N DEL 6
SRR1766444.2574313 chr3 195711012 N chr3 195711283 N DEL 10
SRR1766466.2910937 chr3 195710788 N chr3 195710879 N DEL 20
SRR1766472.6476867 chr3 195710687 N chr3 195710913 N DEL 5
SRR1766465.5399817 chr3 195710789 N chr3 195711373 N DUP 16
SRR1766482.4252815 chr3 195710652 N chr3 195711103 N DEL 10
SRR1766445.5415585 chr3 195711047 N chr3 195711574 N DEL 25
SRR1766483.8839114 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766447.11284297 chr3 195710574 N chr3 195710888 N DUP 25
SRR1766467.3594565 chr3 195710457 N chr3 195711133 N DEL 5
SRR1766455.781242 chr3 195710833 N chr3 195711237 N DUP 10
SRR1766465.2899998 chr3 195710399 N chr3 195711120 N DEL 4
SRR1766442.40652704 chr3 195711093 N chr3 195711182 N DUP 5
SRR1766464.9019755 chr3 195710907 N chr3 195711268 N DEL 9
SRR1766453.258496 chr3 195710732 N chr3 195710868 N DEL 10
SRR1766451.7640748 chr3 195710745 N chr3 195711286 N DEL 20
SRR1766479.10121880 chr3 195710970 N chr3 195711331 N DEL 5
SRR1766442.5212229 chr3 195710447 N chr3 195710673 N DEL 5
SRR1766447.11282149 chr3 195710926 N chr3 195711105 N DUP 15
SRR1766442.33584866 chr3 195710912 N chr3 195711138 N DEL 15
SRR1766471.11641451 chr3 195710833 N chr3 195711192 N DUP 17
SRR1766485.6423844 chr3 195710598 N chr3 195711272 N DUP 2
SRR1766478.7676866 chr3 195710897 N chr3 195711123 N DEL 10
SRR1766452.1746923 chr3 195710507 N chr3 195711273 N DEL 10
SRR1766450.887153 chr3 195710912 N chr3 195711273 N DEL 15
SRR1766451.7640748 chr3 195710469 N chr3 195711055 N DEL 5
SRR1766466.8126136 chr3 195710912 N chr3 195711273 N DEL 5
SRR1766458.2233427 chr3 195710590 N chr3 195710949 N DUP 17
SRR1766471.11429162 chr3 195711058 N chr3 195711372 N DUP 10
SRR1766479.12295867 chr3 195710873 N chr3 195711277 N DUP 6
SRR1766485.135474 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766469.3824058 chr3 195710574 N chr3 195711338 N DUP 7
SRR1766442.12466425 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766468.3137871 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766455.1921365 chr3 195710594 N chr3 195711223 N DUP 2
SRR1766442.19765338 chr3 195710426 N chr3 195711057 N DEL 5
SRR1766470.10029457 chr3 195710779 N chr3 195711363 N DUP 15
SRR1766442.14027655 chr3 195710427 N chr3 195711191 N DUP 5
SRR1766455.2498048 chr3 195710475 N chr3 195710836 N DEL 10
SRR1766443.9803251 chr3 195710457 N chr3 195711133 N DEL 5
SRR1766457.9375446 chr3 195710970 N chr3 195711331 N DEL 5
SRR1766467.2743063 chr3 195710777 N chr3 195711093 N DEL 15
SRR1766469.3750314 chr3 195710745 N chr3 195710881 N DEL 12
SRR1766461.655496 chr3 195710789 N chr3 195711013 N DUP 15
SRR1766442.40725359 chr3 195710907 N chr3 195711133 N DEL 10
SRR1766469.1880462 chr3 195710506 N chr3 195710955 N DUP 6
SRR1766448.6550910 chr3 195710789 N chr3 195711283 N DUP 5
SRR1766467.3570635 chr3 195710420 N chr3 195711622 N DEL 5
SRR1766451.7364049 chr3 195710833 N chr3 195710967 N DUP 23
SRR1766477.5150813 chr3 195710511 N chr3 195711097 N DEL 5
SRR1766479.12986549 chr3 195711012 N chr3 195711148 N DEL 5
SRR1766472.4723707 chr3 195710542 N chr3 195710633 N DEL 15
SRR1766473.2465703 chr3 195710518 N chr3 195711149 N DEL 4
SRR1766462.10039965 chr3 195710701 N chr3 195711240 N DUP 13
SRR1766446.3317050 chr3 195711089 N chr3 195711405 N DEL 26
SRR1766482.8002010 chr3 195710777 N chr3 195711138 N DEL 21
SRR1766460.9110915 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766485.7394197 chr3 195711008 N chr3 195711232 N DUP 10
SRR1766475.1528665 chr3 195710604 N chr3 195711491 N DEL 8
SRR1766443.4940134 chr3 195710628 N chr3 195710897 N DUP 12
SRR1766465.5487908 chr3 195710549 N chr3 195711571 N DEL 2
SRR1766484.9848909 chr3 195710832 N chr3 195711238 N DEL 15
SRR1766483.7588933 chr3 195711023 N chr3 195711159 N DEL 5
SRR1766481.10232930 chr3 195710826 N chr3 195711142 N DEL 10
SRR1766477.11193780 chr3 195710475 N chr3 195711061 N DEL 10
SRR1766467.3593080 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766476.6082131 chr3 195711140 N chr3 195711319 N DUP 10
SRR1766442.14525844 chr3 195710454 N chr3 195710590 N DEL 7
SRR1766475.11050212 chr3 195710912 N chr3 195711228 N DEL 14
SRR1766461.8740540 chr3 195711133 N chr3 195711222 N DUP 9
SRR1766474.7596352 chr3 195710735 N chr3 195711141 N DEL 10
SRR1766482.10001994 chr3 195710789 N chr3 195711148 N DUP 5
SRR1766451.1034834 chr3 195710511 N chr3 195711142 N DEL 10
SRR1766480.8347394 chr3 195710912 N chr3 195711138 N DEL 15
SRR1766482.5996566 chr3 195710912 N chr3 195711273 N DEL 15
SRR1766474.3914400 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766468.5127411 chr3 195710746 N chr3 195711240 N DUP 14
SRR1766442.29999421 chr3 195710475 N chr3 195711061 N DEL 10
SRR1766478.8736120 chr3 195710652 N chr3 195711148 N DEL 10
SRR1766442.22842530 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766460.7485758 chr3 195711023 N chr3 195711247 N DUP 5
SRR1766479.10878674 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766442.20797997 chr3 195710479 N chr3 195711065 N DEL 5
SRR1766442.21743469 chr3 195711012 N chr3 195711148 N DEL 5
SRR1766481.808784 chr3 195710626 N chr3 195711165 N DUP 10
SRR1766442.44460459 chr3 195710745 N chr3 195711286 N DEL 15
SRR1766442.7377992 chr3 195711052 N chr3 195711278 N DEL 5
SRR1766477.10498053 chr3 195711182 N chr3 195711453 N DEL 5
SRR1766442.44343984 chr3 195710998 N chr3 195711087 N DUP 10
SRR1766475.6189519 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766482.8002010 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766453.8621984 chr3 195710664 N chr3 195711115 N DEL 3
SRR1766483.6659795 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766467.8598360 chr3 195711078 N chr3 195711347 N DUP 10
SRR1766460.10906873 chr3 195710897 N chr3 195711123 N DEL 8
SRR1766447.11284297 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766477.2482102 chr3 195710833 N chr3 195711192 N DUP 12
SRR1766474.9856445 chr3 195711103 N chr3 195711372 N DUP 15
SRR1766457.7812382 chr3 195711023 N chr3 195711202 N DUP 11
SRR1766443.3206408 chr3 195710557 N chr3 195711276 N DUP 5
SRR1766481.7925783 chr3 195710520 N chr3 195711466 N DEL 2
SRR1766485.12053858 chr3 195710642 N chr3 195710821 N DUP 5
SRR1766477.7248460 chr3 195710673 N chr3 195711167 N DUP 14
SRR1766449.9957371 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766457.6375563 chr3 195710745 N chr3 195711061 N DEL 10
SRR1766483.4905663 chr3 195710507 N chr3 195711453 N DEL 5
SRR1766459.6172648 chr3 195710656 N chr3 195710745 N DUP 10
SRR1766481.12111596 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766452.8068716 chr3 195710819 N chr3 195711223 N DUP 9
SRR1766470.2259799 chr3 195710732 N chr3 195711093 N DEL 5
SRR1766458.6590782 chr3 195710728 N chr3 195710819 N DEL 19
SRR1766463.8429951 chr3 195710633 N chr3 195711262 N DUP 14
SRR1766479.4039026 chr3 195710431 N chr3 195711150 N DUP 10
SRR1766478.9067448 chr3 195710878 N chr3 195711012 N DUP 9
SRR1766477.937789 chr3 195710701 N chr3 195711195 N DUP 10
SRR1766457.1670099 chr3 195711023 N chr3 195711202 N DUP 11
SRR1766444.2574313 chr3 195711177 N chr3 195711268 N DEL 7
SRR1766453.7617469 chr3 195711013 N chr3 195711192 N DUP 10
SRR1766472.9410030 chr3 195710626 N chr3 195711300 N DUP 5
SRR1766477.5150813 chr3 195710537 N chr3 195710853 N DEL 10
SRR1766467.7695697 chr3 195710754 N chr3 195711070 N DEL 8
SRR1766450.9241373 chr3 195710897 N chr3 195711258 N DEL 5
SRR1766471.5020912 chr3 195710789 N chr3 195711373 N DUP 10
SRR1766457.8733614 chr3 195710878 N chr3 195711372 N DUP 20
SRR1766468.6262396 chr3 195710907 N chr3 195711133 N DEL 12
SRR1766443.6423575 chr3 195710547 N chr3 195710863 N DEL 15
SRR1766457.7812382 chr3 195710921 N chr3 195711147 N DEL 5
SRR1766461.214453 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766470.635997 chr3 195710925 N chr3 195711061 N DEL 10
SRR1766473.6701931 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766451.7364049 chr3 195710897 N chr3 195711213 N DEL 10
SRR1766472.6537572 chr3 195710925 N chr3 195711331 N DEL 10
SRR1766451.5868940 chr3 195711123 N chr3 195711347 N DUP 3
SRR1766486.8021375 chr3 195710428 N chr3 195710652 N DUP 5
SRR1766453.1984628 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766467.2489668 chr3 195711058 N chr3 195711372 N DUP 10
SRR1766467.6409670 chr3 195710907 N chr3 195711133 N DEL 15
SRR1766471.169227 chr3 195710548 N chr3 195711089 N DEL 12
SRR1766463.3808006 chr3 195710833 N chr3 195711237 N DUP 11
SRR1766475.10734632 chr3 195710853 N chr3 195711212 N DUP 10
SRR1766460.8958663 chr3 195710558 N chr3 195711277 N DUP 5
SRR1766478.5474506 chr3 195710853 N chr3 195711212 N DUP 5
SRR1766467.11909659 chr3 195710459 N chr3 195711405 N DEL 19
SRR1766447.408951 chr3 195710878 N chr3 195711012 N DUP 10
SRR1766485.3535942 chr3 195710836 N chr3 195710970 N DUP 17
SRR1766469.10349295 chr3 195711123 N chr3 195711347 N DUP 8
SRR1766472.2927865 chr3 195710656 N chr3 195710745 N DUP 11
SRR1766457.8733614 chr3 195710547 N chr3 195711223 N DEL 5
SRR1766453.1131910 chr3 195710510 N chr3 195710644 N DUP 5
SRR1766455.8921189 chr3 195710745 N chr3 195711331 N DEL 10
SRR1766475.11201508 chr3 195710732 N chr3 195711093 N DEL 10
SRR1766462.1423334 chr3 195710547 N chr3 195711614 N DEL 5
SRR1766465.6527679 chr3 195710712 N chr3 195711073 N DEL 3
SRR1766482.1767085 chr3 195710997 N chr3 195711223 N DEL 6
SRR1766466.6347383 chr3 195710626 N chr3 195711210 N DUP 13
SRR1766458.3852551 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766453.934597 chr3 195710907 N chr3 195711133 N DEL 11
SRR1766442.18697877 chr3 195710869 N chr3 195711183 N DUP 2
SRR1766472.7658271 chr3 195710672 N chr3 195711168 N DEL 11
SRR1766469.2776848 chr3 195710898 N chr3 195711032 N DUP 7
SRR1766445.6863892 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766459.5970256 chr3 195710475 N chr3 195711061 N DEL 10
SRR1766485.568774 chr3 195710477 N chr3 195711198 N DEL 5
SRR1766485.4252295 chr3 195710475 N chr3 195711151 N DEL 10
SRR1766475.336802 chr3 195710470 N chr3 195711056 N DEL 7
SRR1766473.5114181 chr3 195711001 N chr3 195711618 N DEL 5
SRR1766477.4833033 chr3 195710833 N chr3 195710922 N DUP 17
SRR1766482.7511894 chr3 195710595 N chr3 195711406 N DEL 10
SRR1766442.42200322 chr3 195711000 N chr3 195711572 N DEL 5
SRR1766448.5164000 chr3 195710823 N chr3 195711362 N DUP 5
SRR1766467.7695697 chr3 195711048 N chr3 195711362 N DUP 10
SRR1766450.9959800 chr3 195710467 N chr3 195711143 N DEL 5
SRR1766443.6423575 chr3 195711179 N chr3 195711403 N DUP 7
SRR1766470.1238586 chr3 195710457 N chr3 195711133 N DEL 10
SRR1766469.3249156 chr3 195711182 N chr3 195711273 N DEL 7
SRR1766442.44460459 chr3 195710788 N chr3 195710879 N DEL 15
SRR1766453.6263591 chr3 195710590 N chr3 195710814 N DUP 15
SRR1766456.6505169 chr3 195710886 N chr3 195711020 N DUP 10
SRR1766481.401328 chr3 195711048 N chr3 195711362 N DUP 10
SRR1766467.3593080 chr3 195710475 N chr3 195711106 N DEL 5
SRR1766442.36079111 chr3 195710454 N chr3 195710590 N DEL 10
SRR1766444.2118210 chr3 195710427 N chr3 195711236 N DUP 10
SRR1766443.4031060 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766463.1797560 chr3 195710574 N chr3 195711248 N DUP 1
SRR1766484.2346909 chr3 195710652 N chr3 195711058 N DEL 10
SRR1766454.4427009 chr3 195711023 N chr3 195711202 N DUP 10
SRR1766465.4223871 chr3 195710574 N chr3 195711203 N DUP 3
SRR1766485.8375728 chr3 195710970 N chr3 195711331 N DEL 5
SRR1766475.1528665 chr3 195710912 N chr3 195711273 N DEL 5
SRR1766484.2182020 chr3 195710898 N chr3 195710987 N DUP 14
SRR1766442.29532329 chr3 195711452 N chr3 195711619 N DEL 10
SRR1766447.4999222 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766478.7315258 chr3 195710687 N chr3 195710913 N DEL 5
SRR1766477.4976749 chr3 195710462 N chr3 195711048 N DEL 5
SRR1766460.9197482 chr3 195711016 N chr3 195711152 N DEL 5
SRR1766442.24904724 chr3 195711140 N chr3 195711319 N DUP 10
SRR1766463.9254572 chr3 195710475 N chr3 195711061 N DEL 10
SRR1766442.25239751 chr3 195711002 N chr3 195711619 N DEL 5
SRR1766467.6409670 chr3 195710665 N chr3 195711339 N DUP 5
SRR1766478.9067448 chr3 195710679 N chr3 195711085 N DEL 5
SRR1766481.3123362 chr3 195710459 N chr3 195711405 N DEL 19
SRR1766469.10933803 chr3 195710897 N chr3 195711123 N DEL 10
SRR1766445.10054146 chr3 195710868 N chr3 195711227 N DUP 2
SRR1766479.9477024 chr3 195711033 N chr3 195711347 N DUP 5
SRR1766442.28754406 chr3 195710514 N chr3 195711145 N DEL 8
SRR1766449.8071792 chr3 195710507 N chr3 195711273 N DEL 9
SRR1766454.5799610 chr3 195710701 N chr3 195711150 N DUP 15
SRR1766468.3988988 chr3 195711143 N chr3 195711232 N DUP 6
SRR1766477.6908917 chr3 195711012 N chr3 195711148 N DEL 10
SRR1766442.31055253 chr3 195710864 N chr3 195711268 N DUP 6
SRR1766447.4999222 chr3 195710514 N chr3 195711415 N DEL 9
SRR1766446.4027275 chr3 195710897 N chr3 195711258 N DEL 10
SRR1766449.9872863 chr3 195710745 N chr3 195711106 N DEL 10
SRR1766451.1444838 chr3 195710833 N chr3 195711327 N DUP 10
SRR1766479.9603242 chr3 195710925 N chr3 195711151 N DEL 20
SRR1766474.3832772 chr3 195711355 N chr3 195711477 N DEL 11
SRR1766467.1984014 chr3 195710732 N chr3 195711273 N DEL 10
SRR1766477.10566214 chr3 195710598 N chr3 195711227 N DUP 4
SRR1766467.3277409 chr3 195710457 N chr3 195711133 N DEL 13
SRR1766466.2795537 chr3 195711047 N chr3 195711574 N DEL 28
SRR1766451.8266069 chr3 195710475 N chr3 195711061 N DEL 5
SRR1766464.3221854 chr3 195710574 N chr3 195711203 N DUP 2
SRR1766485.10768266 chr3 195710912 N chr3 195711273 N DEL 13
SRR1766465.5903205 chr3 195710659 N chr3 195711200 N DEL 5
SRR1766478.4595593 chr3 195710618 N chr3 195710799 N DEL 5
SRR1766442.17749054 chr3 195710853 N chr3 195711212 N DUP 5
SRR1766442.46715952 chr3 195710789 N chr3 195711013 N DUP 11
SRR1766471.4813397 chr3 195710789 N chr3 195711373 N DUP 22
SRR1766454.618683 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766474.10077014 chr3 195711452 N chr3 195711619 N DEL 10
SRR1766456.3324189 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766459.7117162 chr3 195710745 N chr3 195710881 N DEL 11
SRR1766467.9044595 chr3 195710788 N chr3 195710879 N DEL 20
SRR1766455.3351269 chr3 195710907 N chr3 195711133 N DEL 15
SRR1766480.2665669 chr3 195711123 N chr3 195711347 N DUP 5
SRR1766479.12986549 chr3 195710475 N chr3 195711061 N DEL 5
SRR1766480.5745705 chr3 195710624 N chr3 195711030 N DEL 10
SRR1766460.2495660 chr3 195710789 N chr3 195711148 N DUP 5
SRR1766474.11674016 chr3 195710396 N chr3 195711207 N DEL 5
SRR1766464.4828612 chr3 195710833 N chr3 195711192 N DUP 16
SRR1766484.2346909 chr3 195710508 N chr3 195711274 N DEL 7
SRR1766471.10686592 chr3 195710472 N chr3 195710833 N DEL 20
SRR1766479.12475779 chr3 195710477 N chr3 195711063 N DEL 5
SRR1766473.1750188 chr3 195710493 N chr3 195710897 N DUP 1
SRR1766446.3366022 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766462.493625 chr3 195710475 N chr3 195710656 N DEL 10
SRR1766454.63412 chr3 195710788 N chr3 195710879 N DEL 20
SRR1766475.6189519 chr3 195710580 N chr3 195711031 N DEL 4
SRR1766472.6838449 chr3 195710878 N chr3 195711012 N DUP 10
SRR1766442.16760103 chr3 195710686 N chr3 195711092 N DEL 1
SRR1766470.3593366 chr3 195710916 N chr3 195711097 N DEL 10
SRR1766450.7953199 chr3 195710672 N chr3 195711168 N DEL 10
SRR1766471.11163655 chr3 195710653 N chr3 195711192 N DUP 10
SRR1766478.10257051 chr3 195710476 N chr3 195711195 N DUP 1
SRR1766449.8359246 chr3 195710925 N chr3 195711286 N DEL 10
SRR1766454.8857819 chr3 195710867 N chr3 195711048 N DEL 15
SRR1766470.5933755 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766442.43840210 chr3 195711078 N chr3 195711347 N DUP 10
SRR1766448.9248612 chr3 195710672 N chr3 195711168 N DEL 10
SRR1766474.3832772 chr3 195711360 N chr3 195711572 N DEL 13
SRR1766448.8568638 chr3 195711182 N chr3 195711273 N DEL 1
SRR1766455.5643578 chr3 195710742 N chr3 195711013 N DEL 10
SRR1766446.7445980 chr3 195711183 N chr3 195711409 N DEL 15
SRR1766464.1659129 chr3 195710700 N chr3 195710836 N DEL 15
SRR1766473.2465703 chr3 195710878 N chr3 195711012 N DUP 10
SRR1766458.3098634 chr3 195710897 N chr3 195711123 N DEL 5
SRR1766485.12053858 chr3 195710633 N chr3 195711217 N DUP 15
SRR1766478.5473077 chr3 195710682 N chr3 195711133 N DEL 10
SRR1766479.2058122 chr3 195710656 N chr3 195710925 N DUP 1
SRR1766472.9674977 chr3 195710643 N chr3 195711272 N DUP 10
SRR1766466.6514721 chr3 195710703 N chr3 195711242 N DUP 8
SRR1766454.535141 chr3 195710925 N chr3 195711151 N DEL 10
SRR1766442.21983193 chr3 195710619 N chr3 195711158 N DUP 10
SRR1766473.10023160 chr3 195711012 N chr3 195711148 N DEL 16
SRR1766452.3317975 chr3 195710422 N chr3 195711624 N DEL 5
SRR1766464.416862 chr3 195710833 N chr3 195710922 N DUP 20
SRR1766476.6046694 chr3 195710868 N chr3 195711182 N DUP 5
SRR1766467.9978162 chr3 195710517 N chr3 195710833 N DEL 15
SRR1766472.3839632 chr3 195710628 N chr3 195711347 N DUP 15
SRR1766461.2698733 chr3 195710456 N chr3 195710862 N DEL 5
SRR1766454.4427009 chr3 195710831 N chr3 195711147 N DEL 5
SRR1766442.12466967 chr3 195710507 N chr3 195711408 N DEL 12
SRR1766450.9241373 chr3 195710818 N chr3 195711613 N DUP 20
SRR1766469.3711865 chr3 195710542 N chr3 195710633 N DEL 10
SRR1766465.1693275 chr3 195710700 N chr3 195710836 N DEL 10
SRR1766442.44332938 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766486.7315157 chr3 195711148 N chr3 195711372 N DUP 10
SRR1766457.8737280 chr3 195710897 N chr3 195711258 N DEL 10
SRR1766462.9596106 chr3 195710833 N chr3 195711237 N DUP 10
SRR1766448.4758028 chr3 195711058 N chr3 195711372 N DUP 10
SRR1766448.8109133 chr3 195710659 N chr3 195711245 N DEL 5
SRR1766465.8004613 chr3 195710480 N chr3 195710661 N DEL 10
SRR1766483.12014076 chr18 71578741 N chr18 71578842 N DEL 2
SRR1766461.519050 chr18 71578741 N chr18 71578842 N DEL 5
SRR1766447.11043875 chr18 71578741 N chr18 71578842 N DEL 5
SRR1766469.9280579 chr18 71578741 N chr18 71578842 N DEL 5
SRR1766447.1168348 chr18 71578660 N chr18 71578815 N DUP 5
SRR1766462.6508956 chr18 71578775 N chr18 71578874 N DUP 5
SRR1766475.855396 chr18 71578775 N chr18 71578874 N DUP 5
SRR1766452.8108916 chr18 71578775 N chr18 71578874 N DUP 5
SRR1766443.9152429 chr18 71578775 N chr18 71578874 N DUP 5
SRR1766459.9523322 chr18 71578775 N chr18 71578874 N DUP 5
SRR1766442.10687144 chr18 71578689 N chr18 71578775 N DEL 5
SRR1766462.7730105 chr18 71578689 N chr18 71578775 N DEL 5
SRR1766453.7944194 chr1 204047301 N chr1 204047602 N DEL 3
SRR1766444.4464954 chr14 64895053 N chr14 64895178 N DUP 12
SRR1766474.1360317 chr14 64895068 N chr14 64895243 N DUP 1
SRR1766463.5530793 chr14 64895056 N chr14 64895232 N DUP 7
SRR1766469.3268333 chr9 95568252 N chr9 95568346 N DUP 5
SRR1766464.1152254 chr1 79571551 N chr1 79571707 N DEL 1
SRR1766454.5589754 chr1 79571551 N chr1 79571707 N DEL 2
SRR1766443.4974883 chr1 79571551 N chr1 79571707 N DEL 4
SRR1766459.4665147 chr1 79571551 N chr1 79571707 N DEL 5
SRR1766451.8157929 chr1 79571551 N chr1 79571707 N DEL 9
SRR1766470.3710924 chr1 79571577 N chr1 79571638 N DEL 11
SRR1766483.9491342 chr1 79571577 N chr1 79571638 N DEL 12
SRR1766462.2485562 chr1 79571577 N chr1 79571638 N DEL 18
SRR1766447.9312595 chr1 79571577 N chr1 79571638 N DEL 18
SRR1766468.2163352 chr1 79571577 N chr1 79571638 N DEL 11
SRR1766445.6834832 chr1 79571577 N chr1 79571638 N DEL 9
SRR1766479.2136570 chr1 79571577 N chr1 79571638 N DEL 9
SRR1766464.1152254 chr1 79571577 N chr1 79571638 N DEL 9
SRR1766442.46978073 chr1 79571577 N chr1 79571638 N DEL 9
SRR1766464.1584583 chr1 79571577 N chr1 79571638 N DEL 9
SRR1766470.6782266 chr1 79571577 N chr1 79571638 N DEL 9
SRR1766445.835143 chr1 79571577 N chr1 79571638 N DEL 9
SRR1766458.5205069 chr1 79571542 N chr1 79571640 N DEL 9
SRR1766464.7680293 chr1 79571543 N chr1 79571641 N DEL 9
SRR1766480.3857006 chr1 79571544 N chr1 79571642 N DEL 9
SRR1766442.6934538 chr1 79571637 N chr1 79571733 N DEL 5
SRR1766476.4456532 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766476.3195710 chr1 79571577 N chr1 79571638 N DEL 9
SRR1766472.3299137 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766469.377743 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766442.7662026 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766443.8232803 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766463.4150678 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766448.7277387 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766451.3351771 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766460.8778761 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766480.3442912 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766442.9810081 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766483.5211576 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766442.7521562 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766475.10799737 chr1 79571606 N chr1 79571733 N DEL 5
SRR1766442.34987791 chr1 79571575 N chr1 79571733 N DEL 5
SRR1766464.7210430 chr1 79571575 N chr1 79571733 N DEL 5
SRR1766485.6941882 chr1 79571576 N chr1 79571734 N DEL 5
SRR1766485.6088331 chr1 79571578 N chr1 79571736 N DEL 5
SRR1766471.3873562 chr1 79571584 N chr1 79571742 N DEL 5
SRR1766462.7687431 chr1 79571589 N chr1 79571747 N DEL 1
SRR1766453.193853 chr1 79571589 N chr1 79571747 N DEL 1
SRR1766466.2422678 chr1 79571527 N chr1 79571916 N DUP 5
SRR1766486.245566 chr1 79571742 N chr1 79572213 N DEL 5
SRR1766479.3944827 chr1 79571809 N chr1 79572039 N DUP 5
SRR1766484.4134481 chr1 79571591 N chr1 79571914 N DEL 5
SRR1766459.186126 chr1 79571595 N chr1 79571918 N DEL 5
SRR1766463.3463369 chr1 79571467 N chr1 79571920 N DEL 5
SRR1766444.2960860 chr1 79571471 N chr1 79571957 N DEL 3
SRR1766445.4988124 chr1 79571837 N chr1 79572271 N DEL 3
SRR1766473.1100049 chr1 79571837 N chr1 79572271 N DEL 4
SRR1766484.5726957 chr1 79571837 N chr1 79572271 N DEL 4
SRR1766482.11845042 chr1 79571837 N chr1 79572271 N DEL 6
SRR1766450.351323 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766451.60802 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766443.2923144 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766464.2812842 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766481.11316416 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766483.3428038 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766442.8520686 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766474.7616984 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766483.1754277 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766486.7423014 chr1 79571840 N chr1 79572274 N DEL 7
SRR1766468.1487330 chr1 79571837 N chr1 79572271 N DEL 7
SRR1766460.1984075 chr1 79571837 N chr1 79572271 N DEL 8
SRR1766456.4088034 chr1 79571738 N chr1 79572271 N DEL 9
SRR1766471.5590163 chr1 79571738 N chr1 79572271 N DEL 11
SRR1766451.6894104 chr1 79571738 N chr1 79572271 N DEL 11
SRR1766451.377465 chr1 79571593 N chr1 79571916 N DEL 5
SRR1766450.5211909 chr1 79571468 N chr1 79571921 N DEL 5
SRR1766482.2941539 chr1 79571469 N chr1 79571922 N DEL 5
SRR1766465.5167239 chr1 79571470 N chr1 79571923 N DEL 4
SRR1766473.435674 chr1 79571702 N chr1 79571870 N DUP 5
SRR1766478.2432253 chr1 79571583 N chr1 79572174 N DEL 2
SRR1766470.3219154 chr1 79572283 N chr1 79572412 N DEL 2
SRR1766442.43099332 chr1 79572249 N chr1 79572316 N DEL 9
SRR1766442.34987791 chr1 79571818 N chr1 79572324 N DEL 12
SRR1766454.981903 chr1 79571738 N chr1 79572271 N DEL 9
SRR1766465.4421590 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766442.34633864 chr1 79571738 N chr1 79572271 N DEL 13
SRR1766471.11304270 chr1 79571546 N chr1 79572271 N DEL 13
SRR1766468.4178449 chr1 79571546 N chr1 79572271 N DEL 13
SRR1766483.765213 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766475.3118020 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766459.9780871 chr1 79571546 N chr1 79572271 N DEL 13
SRR1766454.3186304 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766460.8432457 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766474.9231037 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766475.1183310 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766443.7852331 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766460.5991061 chr1 79572047 N chr1 79572283 N DEL 3
SRR1766451.3131881 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766484.4196086 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766461.3837126 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766482.201463 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766443.10484431 chr1 79572044 N chr1 79572280 N DEL 6
SRR1766451.8157929 chr1 79571849 N chr1 79572322 N DEL 7
SRR1766459.4278511 chr1 79572045 N chr1 79572281 N DEL 5
SRR1766471.3873562 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766472.4628388 chr1 79572046 N chr1 79572282 N DEL 4
SRR1766472.8949561 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766459.157507 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766479.10784 chr1 79571884 N chr1 79572324 N DEL 5
SRR1766468.1030876 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766447.9312595 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766468.7833859 chr1 79571851 N chr1 79572324 N DEL 7
SRR1766471.8827931 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766462.6763755 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766471.8768431 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766449.7778003 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766483.5698462 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766450.9872343 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766452.6853322 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766464.1126126 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766448.2060148 chr1 79571818 N chr1 79572324 N DEL 7
SRR1766453.140967 chr1 79571821 N chr1 79572327 N DEL 7
SRR1766470.8936373 chr1 79571823 N chr1 79572329 N DEL 7
SRR1766479.9098947 chr1 79571824 N chr1 79572330 N DEL 7
SRR1766459.2702298 chr1 79572375 N chr1 79572438 N DUP 3
SRR1766442.23727577 chr15 64283737 N chr15 64283877 N DUP 5
SRR1766482.10679612 chr20 62468131 N chr20 62468280 N DEL 5
SRR1766462.10832966 chr20 62468162 N chr20 62468237 N DUP 5
SRR1766485.9742900 chr20 62468304 N chr20 62468453 N DEL 5
SRR1766466.6472936 chr20 62468134 N chr20 62468359 N DEL 3
SRR1766450.6767124 chr20 62468022 N chr20 62468401 N DEL 5
SRR1766478.11854794 chr9 90694383 N chr9 90694506 N DUP 5
SRR1766450.8992540 chr9 90694451 N chr9 90694564 N DUP 5
SRR1766484.2311303 chr9 90694476 N chr9 90694591 N DUP 3
SRR1766443.11159798 chr9 90694480 N chr9 90694838 N DUP 9
SRR1766458.6322359 chr9 90694423 N chr9 90694534 N DEL 8
SRR1766448.10726856 chr9 90694423 N chr9 90694568 N DEL 10
SRR1766474.3124810 chr9 90694495 N chr9 90694568 N DEL 7
SRR1766446.7121008 chr9 90694423 N chr9 90694576 N DEL 7
SRR1766456.3782054 chr9 90694423 N chr9 90694596 N DEL 9
SRR1766468.472974 chr9 90694423 N chr9 90694596 N DEL 9
SRR1766444.4532583 chr9 90694419 N chr9 90694712 N DUP 5
SRR1766484.11213057 chr9 90694623 N chr9 90694744 N DUP 10
SRR1766474.4940835 chr9 90694646 N chr9 90694824 N DUP 11
SRR1766449.10917059 chr9 90694475 N chr9 90694648 N DEL 6
SRR1766474.2813747 chr9 90694600 N chr9 90694685 N DEL 1
SRR1766448.4220388 chr9 90694609 N chr9 90694720 N DEL 3
SRR1766442.20801769 chr9 90694367 N chr9 90694720 N DEL 3
SRR1766479.11860620 chr9 90694564 N chr9 90694745 N DEL 5
SRR1766464.4947309 chr9 90694601 N chr9 90694849 N DEL 5
SRR1766479.13054677 chr9 90694440 N chr9 90694848 N DEL 12
SRR1766449.1601969 chr9 90694430 N chr9 90694836 N DEL 9
SRR1766473.4176554 chr9 90694422 N chr9 90694840 N DEL 3
SRR1766460.9711307 chr3 194352335 N chr3 194352487 N DEL 6
SRR1766480.7379172 chr3 194352311 N chr3 194352574 N DEL 4
SRR1766477.2010859 chr3 194352327 N chr3 194352590 N DEL 5
SRR1766457.3464068 chr3 194352328 N chr3 194352726 N DEL 5
SRR1766456.2591922 chr7 1384768 N chr7 1384842 N DEL 28
SRR1766453.6868035 chr8 138805065 N chr8 138806007 N DEL 30
SRR1766468.6491039 chr8 138805094 N chr8 138805217 N DEL 2
SRR1766444.6219366 chr8 138804912 N chr8 138805343 N DEL 3
SRR1766449.4929856 chr8 138804955 N chr8 138805481 N DEL 2
SRR1766480.2776149 chr8 138805595 N chr8 138806291 N DEL 1
SRR1766485.961294 chr8 138805184 N chr8 138805561 N DEL 1
SRR1766442.9147543 chr8 138804943 N chr8 138805771 N DUP 4
SRR1766454.76778 chr8 138805414 N chr8 138805682 N DEL 13
SRR1766478.1613639 chr8 138805744 N chr8 138805837 N DUP 5
SRR1766468.6437353 chr8 138805111 N chr8 138805740 N DEL 7
SRR1766480.1881716 chr8 138805448 N chr8 138805740 N DEL 12
SRR1766455.2623661 chr8 138804938 N chr8 138805891 N DUP 5
SRR1766486.7169460 chr8 138805175 N chr8 138805798 N DEL 10
SRR1766446.9095398 chr8 138805054 N chr8 138805994 N DUP 10
SRR1766461.3031397 chr8 138805434 N chr8 138806025 N DUP 5
SRR1766460.9763 chr8 138804873 N chr8 138805942 N DEL 7
SRR1766478.4750141 chr8 138805196 N chr8 138805972 N DEL 1
SRR1766480.4933065 chr8 138805462 N chr8 138805968 N DEL 12
SRR1766442.11117306 chr8 138804958 N chr8 138806005 N DEL 5
SRR1766471.5669650 chr8 138804915 N chr8 138806006 N DEL 5
SRR1766453.6868035 chr8 138805066 N chr8 138806008 N DEL 8
SRR1766485.10107641 chr8 138805433 N chr8 138806146 N DUP 4
SRR1766443.1574743 chr8 138804941 N chr8 138806182 N DUP 3
SRR1766449.6096411 chr8 138805315 N chr8 138806197 N DUP 14
SRR1766452.10003270 chr8 138805198 N chr8 138806198 N DUP 5
SRR1766472.11727144 chr8 138805198 N chr8 138806198 N DUP 5
SRR1766459.2573484 chr8 138805198 N chr8 138806198 N DUP 5
SRR1766466.2450056 chr8 138805199 N chr8 138806199 N DUP 5
SRR1766475.4687866 chr8 138806181 N chr8 138806256 N DEL 9
SRR1766476.6070649 chr8 138806181 N chr8 138806256 N DEL 9
SRR1766477.2720172 chr8 138806218 N chr8 138806279 N DEL 21
SRR1766483.5259067 chr8 138806218 N chr8 138806279 N DEL 24
SRR1766453.10004252 chr8 138806218 N chr8 138806279 N DEL 24
SRR1766482.4581115 chr8 138805094 N chr8 138806180 N DEL 19
SRR1766442.6216434 chr8 138805147 N chr8 138806181 N DEL 10
SRR1766461.361097 chr8 138806218 N chr8 138806279 N DEL 17
SRR1766478.10005766 chr8 138806005 N chr8 138806287 N DUP 11
SRR1766480.4873748 chr8 138804955 N chr8 138806182 N DEL 8
SRR1766468.6535455 chr8 138804861 N chr8 138806298 N DUP 7
SRR1766480.679171 chr8 138806199 N chr8 138806308 N DUP 14
SRR1766459.2573484 chr8 138805779 N chr8 138806287 N DEL 9
SRR1766468.4190891 chr8 138805441 N chr8 138806328 N DEL 15
SRR1766479.7239807 chr8 138806070 N chr8 138806329 N DEL 10
SRR1766482.7592090 chr8 138805225 N chr8 138806353 N DEL 5
SRR1766459.5658021 chr8 138805088 N chr8 138806366 N DEL 10
SRR1766483.272223 chr8 138805780 N chr8 138806364 N DEL 15
SRR1766481.7277607 chr8 138805146 N chr8 138806392 N DEL 8
SRR1766449.6096411 chr8 138805669 N chr8 138806401 N DEL 2
SRR1766442.40920424 chr8 138805700 N chr8 138806396 N DEL 5
SRR1766448.1300589 chr8 138805195 N chr8 138806417 N DEL 5
SRR1766483.10336421 chr14 70612030 N chr14 70612165 N DEL 7
SRR1766478.3745896 chr14 70612030 N chr14 70612165 N DEL 9
SRR1766442.32097664 chr16 9676239 N chr16 9676324 N DEL 10
SRR1766477.5740264 chr16 9676241 N chr16 9676326 N DEL 10
SRR1766473.8526256 chr16 9676256 N chr16 9676339 N DEL 4
SRR1766476.6595284 chr16 9676256 N chr16 9676339 N DEL 1
SRR1766484.2759844 chr8 94590769 N chr8 94590850 N DEL 5
SRR1766461.362780 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766446.8673535 chr22 18387819 N chr22 18389317 N DEL 9
SRR1766442.37291015 chr22 18387819 N chr22 18389317 N DEL 14
SRR1766446.10195195 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766478.1374096 chr22 18387819 N chr22 18389317 N DEL 13
SRR1766474.8038828 chr22 18387819 N chr22 18389317 N DEL 8
SRR1766451.5862318 chr22 18387815 N chr22 18389190 N DEL 12
SRR1766442.25580045 chr22 18387815 N chr22 18389190 N DEL 9
SRR1766473.1550864 chr22 18387819 N chr22 18389317 N DEL 9
SRR1766480.3894290 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766461.10893418 chr22 18387821 N chr22 18389216 N DEL 16
SRR1766467.4451300 chr22 18387819 N chr22 18389317 N DEL 8
SRR1766466.253232 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766483.5166676 chr22 18387817 N chr22 18389259 N DEL 9
SRR1766460.1696267 chr22 18387819 N chr22 18389317 N DEL 8
SRR1766475.533854 chr22 18387819 N chr22 18389317 N DEL 8
SRR1766449.6324853 chr22 18387753 N chr22 18388498 N DUP 11
SRR1766463.10308022 chr22 18387821 N chr22 18389216 N DEL 16
SRR1766465.11277751 chr22 18387819 N chr22 18389317 N DEL 8
SRR1766448.10593927 chr22 18387819 N chr22 18389317 N DEL 8
SRR1766483.4408848 chr22 18387817 N chr22 18389259 N DEL 7
SRR1766454.5110384 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766445.10494697 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766470.2806549 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766449.6787736 chr22 18387819 N chr22 18389317 N DEL 9
SRR1766453.120350 chr22 18387820 N chr22 18389262 N DEL 8
SRR1766449.6285817 chr22 18387821 N chr22 18389216 N DEL 16
SRR1766466.2877894 chr22 18387988 N chr22 18388042 N DEL 6
SRR1766485.9767809 chr22 18387960 N chr22 18388065 N DUP 8
SRR1766442.14194275 chr22 18387817 N chr22 18389259 N DEL 7
SRR1766442.6786160 chr22 18387819 N chr22 18389317 N DEL 13
SRR1766486.2857285 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766459.3491401 chr22 18387819 N chr22 18389317 N DEL 13
SRR1766460.7443124 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766472.6563883 chr22 18387819 N chr22 18389317 N DEL 9
SRR1766459.6350600 chr22 18387817 N chr22 18389259 N DEL 9
SRR1766442.25590207 chr22 18387815 N chr22 18389159 N DEL 4
SRR1766486.5100544 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766471.3409642 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766477.2435337 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766464.10167303 chr22 18387819 N chr22 18389317 N DEL 13
SRR1766442.627522 chr22 18387819 N chr22 18389317 N DEL 12
SRR1766463.6239642 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766453.2973441 chr22 18387819 N chr22 18389317 N DEL 9
SRR1766459.8404462 chr22 18388339 N chr22 18389057 N DUP 12
SRR1766485.9898568 chr22 18387821 N chr22 18389216 N DEL 16
SRR1766462.295527 chr22 18387821 N chr22 18389216 N DEL 17
SRR1766466.9704657 chr22 18387815 N chr22 18389190 N DEL 12
SRR1766446.9368363 chr22 18387819 N chr22 18389317 N DEL 7
SRR1766445.9778081 chr12 58598039 N chr12 58598102 N DUP 5
SRR1766467.4444426 chr12 58598054 N chr12 58598123 N DEL 11
SRR1766442.34493468 chr12 58598052 N chr12 58598123 N DEL 9
SRR1766458.7469939 chr12 58598052 N chr12 58598123 N DEL 9
SRR1766483.2597789 chr12 58598058 N chr12 58598127 N DEL 11
SRR1766461.8872403 chr12 58598034 N chr12 58598129 N DEL 9
SRR1766475.2757423 chr12 58598036 N chr12 58598131 N DEL 7
SRR1766462.1882871 chr12 58598037 N chr12 58598132 N DEL 6
SRR1766452.1089578 chr12 58598035 N chr12 58598130 N DEL 8
SRR1766458.7430657 chr12 58598036 N chr12 58598131 N DEL 7
SRR1766446.7563359 chr12 58598037 N chr12 58598134 N DEL 6
SRR1766449.339505 chr8 502785 N chr8 502837 N DUP 5
SRR1766474.3177292 chr8 502811 N chr8 503024 N DEL 3
SRR1766463.2623028 chr8 502863 N chr8 502970 N DEL 4
SRR1766471.9749542 chr8 502871 N chr8 503915 N DEL 10
SRR1766468.1894795 chr8 502904 N chr8 503700 N DEL 1
SRR1766484.2977765 chr8 502923 N chr8 503667 N DEL 4
SRR1766448.7695397 chr8 502758 N chr8 502916 N DUP 5
SRR1766469.6440352 chr8 502890 N chr8 503881 N DEL 15
SRR1766476.9458167 chr8 502747 N chr8 502905 N DUP 10
SRR1766466.2680788 chr8 502760 N chr8 502918 N DUP 5
SRR1766484.1851163 chr8 502898 N chr8 503889 N DEL 15
SRR1766446.2760902 chr8 502944 N chr8 503316 N DEL 5
SRR1766484.2613476 chr8 502758 N chr8 502916 N DUP 5
SRR1766442.5406160 chr8 502766 N chr8 502977 N DUP 1
SRR1766459.10877371 chr8 502819 N chr8 502873 N DEL 5
SRR1766462.3741656 chr8 503004 N chr8 503589 N DEL 5
SRR1766468.411684 chr8 502914 N chr8 503956 N DUP 10
SRR1766451.7719733 chr8 502860 N chr8 502914 N DEL 10
SRR1766452.1336127 chr8 502854 N chr8 502908 N DEL 5
SRR1766478.6657668 chr8 502754 N chr8 502914 N DEL 13
SRR1766477.9232687 chr8 502831 N chr8 502938 N DEL 1
SRR1766461.3768528 chr8 503056 N chr8 503588 N DEL 1
SRR1766452.3233212 chr8 502868 N chr8 503079 N DUP 10
SRR1766453.3917157 chr8 502745 N chr8 503062 N DUP 15
SRR1766450.6298960 chr8 503089 N chr8 504134 N DEL 1
SRR1766447.5116629 chr8 502845 N chr8 503109 N DUP 5
SRR1766474.9940333 chr8 503021 N chr8 503073 N DUP 5
SRR1766486.5016702 chr8 503094 N chr8 503467 N DEL 5
SRR1766458.6835877 chr8 502786 N chr8 503156 N DUP 1
SRR1766450.1299375 chr8 503163 N chr8 503589 N DEL 4
SRR1766464.770196 chr8 502851 N chr8 503064 N DEL 2
SRR1766483.11971083 chr8 502851 N chr8 503064 N DEL 2
SRR1766442.35191377 chr8 503183 N chr8 503556 N DEL 3
SRR1766474.7220807 chr8 502983 N chr8 503141 N DUP 5
SRR1766474.7086772 chr8 503083 N chr8 503913 N DUP 15
SRR1766459.4770579 chr8 503201 N chr8 503874 N DEL 3
SRR1766474.8472392 chr8 503209 N chr8 503582 N DEL 11
SRR1766474.3177292 chr8 502799 N chr8 503118 N DEL 5
SRR1766460.2584201 chr8 503216 N chr8 503483 N DEL 5
SRR1766469.3854778 chr8 503201 N chr8 503874 N DEL 10
SRR1766447.228955 chr8 502978 N chr8 503189 N DUP 9
SRR1766454.4203599 chr8 503201 N chr8 503874 N DEL 10
SRR1766483.7222789 chr8 502840 N chr8 503159 N DEL 10
SRR1766455.7355902 chr8 503183 N chr8 503607 N DUP 10
SRR1766456.3322045 chr8 503108 N chr8 503268 N DEL 15
SRR1766475.2914781 chr8 502842 N chr8 503214 N DEL 10
SRR1766449.439714 chr8 503072 N chr8 503232 N DEL 5
SRR1766447.7788760 chr8 502774 N chr8 503356 N DUP 2
SRR1766446.1508973 chr8 502785 N chr8 503263 N DEL 5
SRR1766471.9749542 chr8 502778 N chr8 503256 N DEL 5
SRR1766478.2408549 chr8 503356 N chr8 504136 N DEL 5
SRR1766469.1389377 chr8 503356 N chr8 504136 N DEL 5
SRR1766467.2669623 chr8 503356 N chr8 504136 N DEL 5
SRR1766445.6372168 chr8 503372 N chr8 504152 N DEL 2
SRR1766470.7093941 chr8 503361 N chr8 504141 N DEL 7
SRR1766462.7980233 chr8 503372 N chr8 504152 N DEL 4
SRR1766443.8211845 chr8 503292 N chr8 503504 N DUP 5
SRR1766470.8872816 chr8 502764 N chr8 503295 N DEL 14
SRR1766471.4867034 chr8 503372 N chr8 504152 N DEL 5
SRR1766445.2484560 chr8 503386 N chr8 504006 N DEL 7
SRR1766483.5664643 chr8 503304 N chr8 503922 N DUP 10
SRR1766479.7689727 chr8 502771 N chr8 503460 N DUP 5
SRR1766470.274256 chr8 502771 N chr8 503460 N DUP 5
SRR1766462.3741656 chr8 502771 N chr8 503460 N DUP 5
SRR1766478.1782770 chr8 503400 N chr8 504020 N DEL 10
SRR1766464.3156060 chr8 502771 N chr8 503460 N DUP 5
SRR1766454.7023090 chr8 503405 N chr8 503670 N DUP 5
SRR1766470.274256 chr8 503401 N chr8 503666 N DUP 5
SRR1766459.3220664 chr8 503403 N chr8 503668 N DUP 5
SRR1766476.2152719 chr8 502745 N chr8 503487 N DUP 11
SRR1766473.5382196 chr8 503035 N chr8 503407 N DEL 5
SRR1766477.3519783 chr8 503036 N chr8 503408 N DEL 5
SRR1766473.5118661 chr8 502978 N chr8 503508 N DUP 10
SRR1766486.2540170 chr8 503467 N chr8 504085 N DUP 10
SRR1766463.4366073 chr8 503020 N chr8 503603 N DUP 2
SRR1766479.5732944 chr8 502843 N chr8 503481 N DEL 4
SRR1766483.9440751 chr8 503020 N chr8 503603 N DUP 5
SRR1766473.9919515 chr8 502778 N chr8 503522 N DEL 10
SRR1766450.1299375 chr8 502778 N chr8 503522 N DEL 10
SRR1766442.43144820 chr8 502844 N chr8 503639 N DUP 5
SRR1766449.7788583 chr8 502856 N chr8 503547 N DEL 6
SRR1766474.8472392 chr8 502803 N chr8 503547 N DEL 5
SRR1766474.5890640 chr8 503652 N chr8 504006 N DEL 5
SRR1766467.2669623 chr8 503554 N chr8 503959 N DUP 5
SRR1766448.4247165 chr8 502725 N chr8 503575 N DEL 19
SRR1766481.2298660 chr8 503037 N chr8 503569 N DEL 1
SRR1766475.3154532 chr8 502843 N chr8 503640 N DEL 7
SRR1766484.381490 chr8 503452 N chr8 503665 N DEL 5
SRR1766475.9926268 chr8 503311 N chr8 503876 N DUP 5
SRR1766484.255249 chr8 503037 N chr8 503781 N DEL 2
SRR1766455.8063520 chr8 503765 N chr8 503905 N DUP 10
SRR1766459.5269282 chr8 502792 N chr8 503940 N DUP 5
SRR1766467.2848120 chr8 503921 N chr8 503973 N DUP 3
SRR1766464.7799382 chr8 503940 N chr8 504101 N DEL 5
SRR1766447.7788760 chr8 502822 N chr8 503919 N DEL 1
SRR1766454.9865753 chr8 503930 N chr8 504249 N DUP 5
SRR1766478.4598638 chr8 502791 N chr8 503941 N DEL 5
SRR1766466.5474389 chr8 503644 N chr8 504050 N DUP 5
SRR1766481.1093183 chr8 502812 N chr8 504067 N DUP 5
SRR1766465.7889520 chr8 502818 N chr8 504073 N DUP 5
SRR1766445.6372168 chr8 503037 N chr8 503975 N DEL 12
SRR1766476.4373402 chr8 502763 N chr8 504124 N DUP 5
SRR1766456.2422347 chr8 503196 N chr8 504082 N DEL 6
SRR1766478.3420881 chr8 503791 N chr8 504093 N DEL 10
SRR1766483.10767576 chr8 503601 N chr8 504115 N DEL 1
SRR1766486.5961332 chr8 503957 N chr8 504118 N DEL 15
SRR1766474.5890640 chr8 503958 N chr8 504119 N DEL 17
SRR1766453.8635391 chr8 502858 N chr8 504168 N DEL 1
SRR1766469.2981189 chr8 502858 N chr8 504168 N DEL 1
SRR1766469.6888198 chr8 504055 N chr8 504216 N DEL 5
SRR1766471.8546668 chr8 503613 N chr8 504234 N DEL 5
SRR1766451.1332878 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766471.12261751 chr6 21924866 N chr6 21925158 N DEL 8
SRR1766460.3952785 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766484.8637781 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766463.5609095 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766484.5995642 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766452.7585819 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766442.46813684 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766483.8263349 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766452.2416066 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766466.8013217 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766453.3667729 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766455.855838 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766467.11708448 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766445.3825181 chr6 21924821 N chr6 21925014 N DEL 5
SRR1766452.7244451 chr6 21924821 N chr6 21925014 N DEL 6
SRR1766460.6410031 chr6 21924878 N chr6 21925069 N DUP 5
SRR1766449.4557653 chr6 21924878 N chr6 21924973 N DUP 5
SRR1766442.32937888 chr6 21924878 N chr6 21924973 N DUP 5
SRR1766460.1114102 chr6 21924884 N chr6 21924979 N DUP 5
SRR1766479.2072560 chr6 21924892 N chr6 21924987 N DUP 1
SRR1766458.1477835 chr6 21924927 N chr6 21925024 N DEL 5
SRR1766459.4479576 chr6 21924878 N chr6 21924973 N DUP 5
SRR1766454.7723045 chr6 21924884 N chr6 21924979 N DUP 5
SRR1766461.8770299 chr6 21924887 N chr6 21924982 N DUP 5
SRR1766459.9457250 chr6 21924833 N chr6 21925026 N DEL 3
SRR1766451.7523505 chr6 21924858 N chr6 21925145 N DUP 1
SRR1766486.6701759 chr6 21925070 N chr6 21925165 N DUP 5
SRR1766442.20428499 chr6 21924977 N chr6 21925077 N DEL 8
SRR1766442.8473460 chr6 21925034 N chr6 21925131 N DEL 5
SRR1766447.203849 chr6 21925034 N chr6 21925131 N DEL 5
SRR1766458.5027861 chr6 21925034 N chr6 21925131 N DEL 5
SRR1766482.8190630 chr6 21925034 N chr6 21925131 N DEL 5
SRR1766461.4946742 chr6 21925034 N chr6 21925131 N DEL 5
SRR1766469.2069644 chr6 21924842 N chr6 21925131 N DEL 5
SRR1766452.2416066 chr6 21924842 N chr6 21925131 N DEL 5
SRR1766445.2672982 chr6 21924842 N chr6 21925131 N DEL 5
SRR1766453.2852723 chr6 21924842 N chr6 21925131 N DEL 5
SRR1766442.23438213 chr6 21924853 N chr6 21925142 N DEL 5
SRR1766474.2170047 chr6 21924857 N chr6 21925146 N DEL 10
SRR1766475.145449 chr9 84409469 N chr9 84409670 N DEL 5
SRR1766468.793562 chr9 84409354 N chr9 84409555 N DEL 5
SRR1766450.1843718 chr19 55320963 N chr19 55321039 N DEL 1
SRR1766462.6434833 chr9 136570000 N chr9 136570141 N DUP 9
SRR1766442.649802 chr9 136569920 N chr9 136570027 N DEL 1
SRR1766450.10415770 chr9 136569930 N chr9 136570065 N DEL 2
SRR1766466.2231024 chr1 4946707 N chr1 4946770 N DUP 5
SRR1766446.1327524 chr1 4946681 N chr1 4946823 N DEL 1
SRR1766457.2101709 chr12 132533240 N chr12 132533435 N DEL 15
SRR1766457.3530397 chr12 132533373 N chr12 132533503 N DEL 5
SRR1766442.38902953 chr12 132533434 N chr12 132533562 N DUP 5
SRR1766477.5629072 chr12 132533434 N chr12 132533562 N DUP 5
SRR1766467.4585161 chr12 132533434 N chr12 132533519 N DUP 5
SRR1766473.1844425 chr19 14314279 N chr19 14314430 N DEL 20
SRR1766457.6497928 chr19 14314321 N chr19 14314434 N DEL 8
SRR1766447.10099578 chr19 14314284 N chr19 14314435 N DEL 10
SRR1766460.7025797 chr9 134729779 N chr9 134729880 N DUP 15
SRR1766486.8180357 chr1 26657770 N chr1 26657941 N DEL 5
SRR1766446.5208260 chrY 10806663 N chrY 10806764 N DEL 2
SRR1766455.5008121 chr13 112028178 N chr13 112028283 N DEL 1
SRR1766476.5691877 chr13 112028213 N chr13 112028511 N DUP 8
SRR1766470.2653132 chr4 110267179 N chr4 110267313 N DEL 5
SRR1766471.4714434 chr4 110267179 N chr4 110267313 N DEL 7
SRR1766451.8778622 chr4 110267179 N chr4 110267313 N DEL 10
SRR1766442.8150643 chr13 114055281 N chr13 114055381 N DUP 5
SRR1766472.992139 chr13 114055282 N chr13 114055382 N DUP 5
SRR1766457.4088739 chr8 60457643 N chr8 60457703 N DEL 1
SRR1766462.2551589 chr8 60457643 N chr8 60457703 N DEL 1
SRR1766446.1827229 chr8 60457643 N chr8 60457703 N DEL 5
SRR1766481.2644960 chr8 60457643 N chr8 60457703 N DEL 5
SRR1766455.4441729 chr16 938438 N chr16 938605 N DEL 10
SRR1766466.8554651 chr5 108387688 N chr5 108387836 N DEL 3
SRR1766458.1750505 chr5 108387690 N chr5 108387836 N DEL 5
SRR1766460.10470763 chr5 108387690 N chr5 108387836 N DEL 5
SRR1766460.3865548 chr20 51961807 N chr20 51961932 N DEL 1
SRR1766460.2212240 chr20 51961825 N chr20 51961881 N DEL 17
SRR1766481.2524873 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766442.42263299 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766448.11007892 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766463.9881219 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766462.4506747 chr20 51961825 N chr20 51961881 N DEL 20
SRR1766443.4588696 chr20 51961833 N chr20 51961884 N DUP 4
SRR1766484.8808183 chr20 51961808 N chr20 51961869 N DUP 13
SRR1766448.9185081 chr20 51961808 N chr20 51961869 N DUP 14
SRR1766478.4537233 chr20 51961808 N chr20 51961869 N DUP 11
SRR1766477.10973196 chr20 51961825 N chr20 51961908 N DUP 2
SRR1766480.701141 chr20 51961825 N chr20 51961908 N DUP 5
SRR1766442.42031432 chr20 51961825 N chr20 51961908 N DUP 7
SRR1766454.9791823 chr20 51961825 N chr20 51961908 N DUP 8
SRR1766482.5816062 chr20 51961860 N chr20 51961918 N DEL 13
SRR1766445.5371765 chr20 51961860 N chr20 51961918 N DEL 14
SRR1766442.12650950 chr20 51961827 N chr20 51961918 N DEL 12
SRR1766455.5205531 chr6 68875206 N chr6 68875313 N DEL 2
SRR1766472.5846179 chr5 139446617 N chr5 139446678 N DUP 7
SRR1766481.9655942 chr5 139446617 N chr5 139446678 N DUP 16
SRR1766473.4289833 chr5 139446634 N chr5 139446711 N DUP 7
SRR1766480.2158684 chr5 139446591 N chr5 139446644 N DEL 2
SRR1766472.1673771 chr14 97895786 N chr14 97896012 N DUP 5
SRR1766455.7374344 chr14 97895787 N chr14 97896013 N DUP 5
SRR1766449.1774319 chr14 97895814 N chr14 97895905 N DUP 5
SRR1766467.5821614 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766459.348981 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766484.5847301 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766459.1242378 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766470.4484043 chr20 30503974 N chr20 30504204 N DEL 5
SRR1766482.4850044 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766466.11192490 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766445.10358410 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766479.5788744 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766477.11652881 chr20 30503985 N chr20 30504215 N DEL 5
SRR1766459.5635024 chr20 30504032 N chr20 30504215 N DEL 5
SRR1766477.724543 chr20 30504032 N chr20 30504215 N DEL 5
SRR1766468.3461841 chr20 30503835 N chr20 30504068 N DUP 5
SRR1766447.2372633 chr20 30504003 N chr20 30504231 N DUP 5
SRR1766475.5987311 chr20 30504010 N chr20 30504238 N DUP 1
SRR1766453.9103258 chr20 30504010 N chr20 30504238 N DUP 1
SRR1766469.4138406 chr21 30210368 N chr21 30210452 N DEL 18
SRR1766442.23746175 chr21 30210368 N chr21 30210452 N DEL 18
SRR1766474.3070299 chr21 30210368 N chr21 30210452 N DEL 18
SRR1766453.2777982 chr21 30210371 N chr21 30210421 N DUP 21
SRR1766478.9624827 chr21 30210371 N chr21 30210421 N DUP 25
SRR1766460.2600477 chr21 30210328 N chr21 30210459 N DUP 11
SRR1766442.26075966 chr21 30210443 N chr21 30210505 N DEL 11
SRR1766477.5122969 chr21 30210443 N chr21 30210505 N DEL 11
SRR1766442.47170639 chr21 30210441 N chr21 30210505 N DEL 13
SRR1766446.1279658 chr21 30210368 N chr21 30210509 N DEL 9
SRR1766481.13058358 chr1 152910417 N chr1 152910808 N DEL 5
SRR1766483.2051446 chr1 152910446 N chr1 152911137 N DEL 5
SRR1766477.3189701 chr1 152910473 N chr1 152910984 N DEL 2
SRR1766477.5047197 chr1 152910459 N chr1 152910910 N DEL 35
SRR1766484.7504615 chr1 152910444 N chr1 152910715 N DEL 20
SRR1766469.4894138 chr1 152910510 N chr1 152910751 N DEL 3
SRR1766478.5480002 chr1 152910471 N chr1 152910560 N DUP 5
SRR1766481.4143107 chr1 152910584 N chr1 152910855 N DEL 5
SRR1766472.5054308 chr1 152910467 N chr1 152910676 N DUP 15
SRR1766474.2656039 chr1 152910467 N chr1 152910586 N DUP 10
SRR1766475.4591905 chr1 152910598 N chr1 152910959 N DEL 10
SRR1766473.7371420 chr1 152910605 N chr1 152910876 N DEL 7
SRR1766470.4229988 chr1 152910467 N chr1 152910676 N DUP 12
SRR1766479.6615232 chr1 152910718 N chr1 152910959 N DEL 5
SRR1766476.2082186 chr1 152910718 N chr1 152910959 N DEL 10
SRR1766442.6346928 chr1 152910725 N chr1 152910876 N DEL 10
SRR1766469.1778429 chr1 152910722 N chr1 152910963 N DEL 10
SRR1766461.10997945 chr1 152910702 N chr1 152910943 N DEL 18
SRR1766468.5389221 chr1 152910505 N chr1 152910656 N DEL 5
SRR1766442.1937426 chr1 152910562 N chr1 152910713 N DEL 20
SRR1766473.7020687 chr1 152910460 N chr1 152910579 N DUP 10
SRR1766466.8512346 chr1 152910775 N chr1 152910956 N DEL 5
SRR1766473.1929648 chr1 152910785 N chr1 152910966 N DEL 3
SRR1766477.8541968 chr1 152910808 N chr1 152910959 N DEL 6
SRR1766474.5184617 chr1 152910808 N chr1 152910959 N DEL 7
SRR1766482.10614598 chr1 152910812 N chr1 152910963 N DEL 10
SRR1766442.8667672 chr1 152910468 N chr1 152910857 N DUP 14
SRR1766479.4135798 chr1 152910751 N chr1 152910900 N DUP 5
SRR1766443.2486898 chr1 152910474 N chr1 152910833 N DUP 15
SRR1766443.1604200 chr1 152910431 N chr1 152910762 N DEL 4
SRR1766478.6407112 chr1 152910492 N chr1 152910763 N DEL 3
SRR1766457.5372066 chr1 152910864 N chr1 152910985 N DEL 5
SRR1766464.2543136 chr1 152910530 N chr1 152910801 N DEL 20
SRR1766469.4745346 chr1 152910864 N chr1 152911216 N DEL 5
SRR1766485.8810549 chr1 152910808 N chr1 152910897 N DUP 10
SRR1766468.2904263 chr1 152910904 N chr1 152911085 N DEL 12
SRR1766471.5759242 chr1 152910525 N chr1 152910856 N DEL 9
SRR1766485.4980742 chr1 152910926 N chr1 152911167 N DEL 5
SRR1766457.8542648 chr1 152910449 N chr1 152910840 N DEL 5
SRR1766444.374611 chr1 152910560 N chr1 152910891 N DEL 45
SRR1766446.190333 chr1 152910747 N chr1 152910838 N DEL 5
SRR1766486.5821747 chr1 152910460 N chr1 152910969 N DUP 3
SRR1766450.2000008 chr1 152910528 N chr1 152910859 N DEL 5
SRR1766467.9626364 chr1 152910495 N chr1 152910856 N DEL 18
SRR1766483.2051446 chr1 152910545 N chr1 152910876 N DEL 15
SRR1766456.1192869 chr1 152910860 N chr1 152911360 N DUP 5
SRR1766442.23555628 chr1 152910419 N chr1 152910870 N DEL 1
SRR1766442.34098364 chr1 152910515 N chr1 152910876 N DEL 18
SRR1766446.1888144 chr1 152910424 N chr1 152910875 N DEL 5
SRR1766461.10997945 chr1 152910915 N chr1 152911004 N DUP 5
SRR1766455.6899229 chr1 152910916 N chr1 152911005 N DUP 10
SRR1766468.2073554 chr1 152910492 N chr1 152910943 N DEL 10
SRR1766477.438229 chr1 152910474 N chr1 152911013 N DUP 15
SRR1766447.6054186 chr1 152910510 N chr1 152910961 N DEL 17
SRR1766448.115485 chr1 152910590 N chr1 152911011 N DEL 29
SRR1766475.4591905 chr1 152910492 N chr1 152910973 N DEL 1
SRR1766443.2486898 chr1 152910902 N chr1 152911023 N DEL 5
SRR1766467.5614620 chr1 152911058 N chr1 152911318 N DUP 5
SRR1766451.6599576 chr1 152910500 N chr1 152911071 N DEL 14
SRR1766481.1817538 chr1 152911091 N chr1 152911291 N DUP 3
SRR1766477.8541968 chr1 152910498 N chr1 152911099 N DEL 10
SRR1766483.3118710 chr1 152911016 N chr1 152911137 N DEL 16
SRR1766452.8789642 chr1 152910977 N chr1 152911207 N DUP 5
SRR1766485.11975511 chr1 152911017 N chr1 152911108 N DEL 4
SRR1766481.13058358 chr1 152910988 N chr1 152911139 N DEL 10
SRR1766473.1929648 chr1 152910986 N chr1 152911137 N DEL 10
SRR1766455.6368920 chr1 152911003 N chr1 152911205 N DEL 10
SRR1766466.1015030 chr1 152910934 N chr1 152911175 N DEL 5
SRR1766469.1778429 chr1 152910973 N chr1 152911184 N DEL 5
SRR1766474.2656039 chr1 152910488 N chr1 152911290 N DEL 5
SRR1766448.5359956 chr1 152910573 N chr1 152911375 N DEL 38
SRR1766468.7180568 chr1 152910873 N chr1 152911375 N DEL 22
SRR1766473.7020687 chr1 152910503 N chr1 152911365 N DEL 4
SRR1766472.5154068 chr1 152910931 N chr1 152911523 N DEL 2
SRR1766444.126691 chr1 152911161 N chr1 152911513 N DEL 12
SRR1766454.9217799 chr2 3110861 N chr2 3110982 N DUP 1
SRR1766444.6103202 chr2 3110945 N chr2 3111003 N DUP 4
SRR1766456.4777182 chr12 128469805 N chr12 128469862 N DEL 5
SRR1766453.4008033 chr12 128469805 N chr12 128469862 N DEL 5
SRR1766451.5327738 chr12 128469805 N chr12 128469862 N DEL 5
SRR1766450.2219045 chr17 79412044 N chr17 79412167 N DEL 5
SRR1766483.2376317 chr17 79412044 N chr17 79412167 N DEL 5
SRR1766483.1377171 chr17 79412044 N chr17 79412167 N DEL 5
SRR1766484.1732583 chr17 79412044 N chr17 79412167 N DEL 5
SRR1766475.10343417 chr17 79412044 N chr17 79412167 N DEL 5
SRR1766483.2055950 chr17 79412060 N chr17 79412181 N DUP 5
SRR1766466.7653531 chr17 79412061 N chr17 79412182 N DUP 5
SRR1766442.37309050 chr17 79412062 N chr17 79412183 N DUP 5
SRR1766450.10426767 chr17 79412060 N chr17 79412181 N DUP 3
SRR1766474.11587450 chr17 79412060 N chr17 79412181 N DUP 5
SRR1766467.7344065 chr17 79412071 N chr17 79412192 N DUP 4
SRR1766442.15255955 chr8 53947673 N chr8 53947742 N DEL 5
SRR1766461.10462432 chr8 53947673 N chr8 53947742 N DEL 5
SRR1766486.139652 chr8 53947673 N chr8 53947742 N DEL 5
SRR1766463.6024088 chr8 53947673 N chr8 53947742 N DEL 5
SRR1766448.7910398 chr8 53947673 N chr8 53947742 N DEL 5
SRR1766459.6085056 chr8 53947673 N chr8 53947742 N DEL 5
SRR1766485.2564690 chr8 53947673 N chr8 53947742 N DEL 5
SRR1766460.4209150 chr8 53947657 N chr8 53947829 N DEL 5
SRR1766443.7399887 chr8 53947605 N chr8 53947742 N DEL 5
SRR1766444.4043028 chr8 53947728 N chr8 53948216 N DUP 5
SRR1766474.6590917 chr8 53947793 N chr8 53947934 N DEL 5
SRR1766451.5475424 chr8 53947793 N chr8 53947934 N DEL 5
SRR1766454.4706499 chr8 53947793 N chr8 53947934 N DEL 5
SRR1766459.2719441 chr8 53947793 N chr8 53947934 N DEL 5
SRR1766474.7823885 chr8 53947793 N chr8 53947934 N DEL 5
SRR1766452.8096064 chr8 53947758 N chr8 53947934 N DEL 5
SRR1766477.6852517 chr8 53947758 N chr8 53947934 N DEL 5
SRR1766486.1706081 chr8 53947764 N chr8 53947940 N DEL 5
SRR1766466.429651 chr8 53947766 N chr8 53947942 N DEL 5
SRR1766469.4159881 chr8 53947768 N chr8 53947944 N DEL 5
SRR1766448.10025853 chr8 53947770 N chr8 53947946 N DEL 3
SRR1766477.6852517 chr8 53948535 N chr8 53949379 N DEL 5
SRR1766478.3413941 chr8 53948538 N chr8 53949132 N DEL 5
SRR1766466.5657857 chr8 53948538 N chr8 53949132 N DEL 5
SRR1766455.440908 chr8 53948538 N chr8 53949132 N DEL 5
SRR1766474.132880 chr8 53948483 N chr8 53948548 N DUP 5
SRR1766459.6193818 chr8 53948568 N chr8 53949445 N DEL 2
SRR1766480.5367214 chr8 53948069 N chr8 53948492 N DEL 10
SRR1766475.10239803 chr8 53948571 N chr8 53949132 N DEL 20
SRR1766458.4485813 chr8 53948469 N chr8 53948534 N DEL 12
SRR1766452.789325 chr8 53948564 N chr8 53949406 N DUP 5
SRR1766464.1550396 chr8 53948564 N chr8 53949156 N DUP 5
SRR1766460.8989042 chr8 53948671 N chr8 53949139 N DEL 1
SRR1766446.4554292 chr8 53948564 N chr8 53949156 N DUP 5
SRR1766475.9441953 chr8 53948564 N chr8 53949156 N DUP 5
SRR1766448.4220291 chr8 53948499 N chr8 53948566 N DEL 5
SRR1766452.10203243 chr8 53948078 N chr8 53948567 N DEL 1
SRR1766456.6386289 chr8 53948150 N chr8 53948569 N DEL 5
SRR1766442.3697057 chr8 53948546 N chr8 53948702 N DUP 19
SRR1766461.8517233 chr8 53948579 N chr8 53948640 N DUP 8
SRR1766458.2724304 chr8 53948579 N chr8 53948640 N DUP 7
SRR1766475.1319809 chr8 53948579 N chr8 53948640 N DUP 7
SRR1766457.1535324 chr8 53948546 N chr8 53948702 N DUP 15
SRR1766484.975708 chr8 53948681 N chr8 53948775 N DEL 10
SRR1766450.3178060 chr8 53948579 N chr8 53948640 N DUP 6
SRR1766451.734687 chr8 53948694 N chr8 53949379 N DEL 19
SRR1766450.5317269 chr8 53948650 N chr8 53948775 N DEL 9
SRR1766464.5791201 chr8 53948650 N chr8 53948775 N DEL 9
SRR1766474.8039837 chr8 53948546 N chr8 53948671 N DUP 14
SRR1766443.2383968 chr8 53948546 N chr8 53948671 N DUP 14
SRR1766459.10040263 chr8 53948650 N chr8 53948775 N DEL 9
SRR1766453.3326613 chr8 53948088 N chr8 53948579 N DEL 5
SRR1766456.5768170 chr8 53948717 N chr8 53948813 N DEL 1
SRR1766483.1400840 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766455.209010 chr8 53948650 N chr8 53948744 N DEL 7
SRR1766459.4283077 chr8 53948546 N chr8 53948702 N DUP 10
SRR1766459.3073024 chr8 53948088 N chr8 53948579 N DEL 5
SRR1766483.7556167 chr8 53948650 N chr8 53948744 N DEL 9
SRR1766443.3007941 chr8 53948546 N chr8 53948671 N DUP 14
SRR1766472.10061483 chr8 53948546 N chr8 53948702 N DUP 12
SRR1766480.5367214 chr8 53948546 N chr8 53948702 N DUP 12
SRR1766444.7016915 chr8 53948579 N chr8 53948640 N DUP 6
SRR1766471.3337781 chr8 53948546 N chr8 53948702 N DUP 15
SRR1766477.10730121 chr8 53948681 N chr8 53948775 N DEL 14
SRR1766451.10491113 chr8 53948579 N chr8 53948640 N DUP 10
SRR1766482.3077480 chr8 53948546 N chr8 53948702 N DUP 18
SRR1766448.6887847 chr8 53948733 N chr8 53948798 N DEL 5
SRR1766443.453978 chr8 53948461 N chr8 53948809 N DUP 5
SRR1766459.7983865 chr8 53948546 N chr8 53948671 N DUP 14
SRR1766472.6925159 chr8 53948681 N chr8 53948775 N DEL 14
SRR1766472.3520083 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766478.7083075 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766477.7993044 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766453.6186332 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766486.8335902 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766451.9742482 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766458.6096115 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766467.3611520 chr8 53948650 N chr8 53948775 N DEL 10
SRR1766466.5657857 chr8 53948619 N chr8 53948775 N DEL 7
SRR1766475.9760433 chr8 53948619 N chr8 53948775 N DEL 6
SRR1766459.235554 chr8 53948619 N chr8 53948775 N DEL 5
SRR1766461.7130029 chr8 53948619 N chr8 53948775 N DEL 5
SRR1766461.8517233 chr8 53948619 N chr8 53948775 N DEL 5
SRR1766484.1150369 chr8 53948619 N chr8 53948775 N DEL 5
SRR1766452.9734761 chr8 53948635 N chr8 53949039 N DEL 10
SRR1766479.524443 chr8 53948635 N chr8 53949039 N DEL 12
SRR1766442.43476354 chr8 53948573 N chr8 53948793 N DEL 4
SRR1766451.8329546 chr8 53948588 N chr8 53948808 N DEL 5
SRR1766453.5991941 chr8 53948588 N chr8 53948808 N DEL 5
SRR1766460.5722005 chr8 53948588 N chr8 53948808 N DEL 5
SRR1766475.2137122 chr8 53948588 N chr8 53948808 N DEL 5
SRR1766448.3359006 chr8 53948588 N chr8 53948808 N DEL 5
SRR1766456.725851 chr8 53948555 N chr8 53948808 N DEL 5
SRR1766472.554390 chr8 53948555 N chr8 53948808 N DEL 5
SRR1766461.7248765 chr8 53947491 N chr8 53949019 N DEL 4
SRR1766465.9141214 chr8 53948555 N chr8 53948808 N DEL 5
SRR1766460.1204472 chr8 53948555 N chr8 53948808 N DEL 5
SRR1766461.7911605 chr8 53948555 N chr8 53948808 N DEL 5
SRR1766442.11481844 chr8 53948813 N chr8 53949469 N DUP 10
SRR1766472.3450154 chr8 53948568 N chr8 53948790 N DEL 10
SRR1766442.17659267 chr8 53948765 N chr8 53949169 N DUP 5
SRR1766473.1960105 chr8 53948557 N chr8 53948810 N DEL 5
SRR1766454.1159425 chr8 53948079 N chr8 53948820 N DEL 3
SRR1766486.3895286 chr8 53948808 N chr8 53949148 N DUP 5
SRR1766477.6496736 chr8 53948808 N chr8 53949148 N DUP 5
SRR1766458.3558332 chr8 53948561 N chr8 53948814 N DEL 5
SRR1766457.5540177 chr8 53948555 N chr8 53948808 N DEL 5
SRR1766475.11456791 chr8 53948080 N chr8 53948790 N DEL 7
SRR1766442.42960044 chr8 53948556 N chr8 53948809 N DEL 5
SRR1766474.11750021 chr8 53948080 N chr8 53948790 N DEL 8
SRR1766443.7087286 chr8 53948555 N chr8 53948808 N DEL 5
SRR1766483.1589819 chr8 53948558 N chr8 53948811 N DEL 5
SRR1766457.8191312 chr8 53948559 N chr8 53948812 N DEL 5
SRR1766454.10800682 chr8 53948079 N chr8 53948820 N DEL 3
SRR1766446.9871823 chr8 53948808 N chr8 53949148 N DUP 5
SRR1766442.34832224 chr8 53949025 N chr8 53949148 N DUP 5
SRR1766481.6853877 chr8 53948808 N chr8 53949148 N DUP 5
SRR1766455.440908 chr8 53949056 N chr8 53949148 N DUP 5
SRR1766446.7915095 chr8 53949087 N chr8 53949148 N DUP 5
SRR1766457.8578835 chr8 53948581 N chr8 53949142 N DEL 2
SRR1766467.209832 chr8 53949193 N chr8 53949382 N DEL 2
SRR1766449.10901844 chr8 53949193 N chr8 53949382 N DEL 3
SRR1766486.901531 chr8 53949193 N chr8 53949382 N DEL 4
SRR1766448.3359006 chr8 53949358 N chr8 53949423 N DUP 23
SRR1766444.7125359 chr8 53949351 N chr8 53949416 N DUP 22
SRR1766460.6027258 chr8 53949349 N chr8 53949414 N DUP 20
SRR1766473.1960105 chr8 53949349 N chr8 53949414 N DUP 26
SRR1766442.4347839 chr8 53949349 N chr8 53949414 N DUP 25
SRR1766481.1865092 chr8 53949349 N chr8 53949414 N DUP 25
SRR1766460.5722005 chr8 53949349 N chr8 53949414 N DUP 15
SRR1766442.3386806 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766454.3170456 chr8 53949349 N chr8 53949414 N DUP 16
SRR1766461.10896229 chr8 53949349 N chr8 53949414 N DUP 21
SRR1766475.6495258 chr8 53949349 N chr8 53949414 N DUP 18
SRR1766485.4518706 chr8 53949349 N chr8 53949414 N DUP 18
SRR1766442.26590434 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766443.2522726 chr8 53949349 N chr8 53949414 N DUP 18
SRR1766451.3608378 chr8 53949349 N chr8 53949414 N DUP 22
SRR1766474.3445500 chr8 53949349 N chr8 53949414 N DUP 23
SRR1766482.3077480 chr8 53949349 N chr8 53949414 N DUP 18
SRR1766485.9463329 chr8 53949349 N chr8 53949414 N DUP 22
SRR1766486.11420708 chr8 53949349 N chr8 53949414 N DUP 17
SRR1766451.10491113 chr8 53949349 N chr8 53949414 N DUP 15
SRR1766479.1620539 chr8 53949349 N chr8 53949414 N DUP 15
SRR1766470.2756996 chr8 53949349 N chr8 53949414 N DUP 16
SRR1766465.9141214 chr8 53949349 N chr8 53949414 N DUP 17
SRR1766451.32847 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766451.3859206 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766474.8039837 chr8 53949349 N chr8 53949414 N DUP 19
SRR1766460.441049 chr8 53949349 N chr8 53949414 N DUP 21
SRR1766477.635213 chr8 53949349 N chr8 53949414 N DUP 22
SRR1766486.8335902 chr8 53949349 N chr8 53949414 N DUP 22
SRR1766448.4220291 chr8 53949349 N chr8 53949414 N DUP 24
SRR1766463.2129608 chr8 53949349 N chr8 53949414 N DUP 24
SRR1766469.8102695 chr8 53949349 N chr8 53949414 N DUP 24
SRR1766453.2819308 chr8 53949349 N chr8 53949414 N DUP 25
SRR1766481.11739291 chr8 53949193 N chr8 53949382 N DEL 12
SRR1766465.5298271 chr8 53949193 N chr8 53949382 N DEL 12
SRR1766472.3378987 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766448.8703754 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766478.3222391 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766452.5856556 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766458.6502372 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766481.6853877 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766442.39466710 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766455.4331222 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766476.5927921 chr8 53949162 N chr8 53949382 N DEL 12
SRR1766460.8989042 chr8 53948503 N chr8 53949382 N DEL 12
SRR1766478.231747 chr8 53947542 N chr8 53949383 N DEL 12
SRR1766442.2788552 chr8 53947544 N chr8 53949385 N DEL 12
SRR1766473.3207979 chr3 68370513 N chr3 68370588 N DUP 13
SRR1766463.4837440 chr3 68370481 N chr3 68370544 N DUP 10
SRR1766450.688529 chr1 193564085 N chr1 193564174 N DUP 1
SRR1766486.3462545 chr1 193564094 N chr1 193564157 N DUP 20
SRR1766471.8347138 chr1 193564152 N chr1 193564215 N DUP 24
SRR1766476.3882521 chr1 193564152 N chr1 193564215 N DUP 21
SRR1766475.4698443 chr1 193564152 N chr1 193564215 N DUP 18
SRR1766473.10071648 chr1 193564152 N chr1 193564215 N DUP 18
SRR1766442.25832369 chr1 193564152 N chr1 193564215 N DUP 18
SRR1766486.4843192 chr1 193564094 N chr1 193564157 N DUP 14
SRR1766483.11307293 chr1 193564152 N chr1 193564215 N DUP 17
SRR1766485.7714912 chr1 193564152 N chr1 193564215 N DUP 10
SRR1766451.4404855 chr1 193564152 N chr1 193564215 N DUP 11
SRR1766478.7697483 chr1 193564069 N chr1 193564152 N DEL 5
SRR1766442.26991531 chr1 193564115 N chr1 193564210 N DEL 3
SRR1766447.11444853 chr1 193564108 N chr1 193564235 N DEL 13
SRR1766457.8214793 chr1 193564109 N chr1 193564236 N DEL 12
SRR1766450.3142331 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766442.4206423 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766463.6903386 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766466.6520294 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766482.4059033 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766455.6058643 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766483.9242974 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766473.7538231 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766478.85808 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766485.11068888 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766464.7524560 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766476.8699710 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766442.36381810 chr1 193564447 N chr1 193564506 N DUP 14
SRR1766472.8079996 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766477.6387356 chr1 193564454 N chr1 193564513 N DUP 12
SRR1766451.7150110 chr1 193564447 N chr1 193564506 N DUP 10
SRR1766442.9353135 chr1 193564447 N chr1 193564506 N DUP 9
SRR1766485.11068888 chr1 193564447 N chr1 193564506 N DUP 8
SRR1766442.3212682 chr1 193564454 N chr1 193564513 N DUP 8
SRR1766482.7926549 chr1 193564447 N chr1 193564506 N DUP 10
SRR1766454.10975702 chr1 193564454 N chr1 193564513 N DUP 11
SRR1766443.8129339 chr1 193564447 N chr1 193564506 N DUP 8
SRR1766458.341289 chr1 193564447 N chr1 193564506 N DUP 8
SRR1766461.3014532 chr1 193564449 N chr1 193564508 N DUP 8
SRR1766473.7800479 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766485.11732669 chr1 193564447 N chr1 193564506 N DUP 10
SRR1766442.12520589 chr1 193564454 N chr1 193564513 N DUP 14
SRR1766474.8652019 chr1 193564447 N chr1 193564506 N DUP 11
SRR1766442.34783777 chr1 193564380 N chr1 193564447 N DEL 7
SRR1766451.318366 chr1 193564383 N chr1 193564450 N DEL 7
SRR1766442.4968880 chr1 193564356 N chr1 193564453 N DEL 7
SRR1766486.9867147 chr19 49064573 N chr19 49064651 N DUP 5
SRR1766479.9981107 chr19 49064619 N chr19 49064743 N DEL 5
SRR1766462.9034736 chr19 49064598 N chr19 49064801 N DEL 2
SRR1766442.9398036 chr4 47123595 N chr4 47123755 N DEL 4
SRR1766478.9799347 chr4 47123595 N chr4 47123755 N DEL 5
SRR1766445.8305075 chr4 47123595 N chr4 47123755 N DEL 5
SRR1766485.8423609 chr4 47123600 N chr4 47123802 N DUP 3
SRR1766457.1515191 chr4 47123601 N chr4 47123803 N DUP 2
SRR1766475.2271207 chr4 47123656 N chr4 47123728 N DEL 8
SRR1766476.5950297 chr4 47123656 N chr4 47123728 N DEL 10
SRR1766466.8043261 chr4 47123656 N chr4 47123728 N DEL 11
SRR1766481.6991814 chr4 47123656 N chr4 47123728 N DEL 12
SRR1766458.6776830 chr4 47123656 N chr4 47123728 N DEL 16
SRR1766462.5339398 chr4 47123656 N chr4 47123728 N DEL 16
SRR1766479.11486539 chr4 47123656 N chr4 47123728 N DEL 32
SRR1766468.7902720 chr4 47123656 N chr4 47123728 N DEL 28
SRR1766473.7989262 chr4 47123656 N chr4 47123728 N DEL 16
SRR1766469.668495 chr4 47123656 N chr4 47123728 N DEL 29
SRR1766461.7605809 chr4 47123591 N chr4 47123729 N DEL 14
SRR1766442.5011230 chr4 47123591 N chr4 47123729 N DEL 14
SRR1766447.8537721 chr4 47123615 N chr4 47123731 N DEL 12
SRR1766449.7330584 chr4 47123584 N chr4 47123739 N DEL 4
SRR1766453.7968916 chr4 47123584 N chr4 47123739 N DEL 4
SRR1766458.7859320 chr4 47123582 N chr4 47123737 N DEL 6
SRR1766460.4105720 chr4 47123618 N chr4 47123734 N DEL 4
SRR1766461.9421595 chr4 47123619 N chr4 47123735 N DEL 8
SRR1766463.2537939 chr4 47123619 N chr4 47123735 N DEL 8
SRR1766479.3554254 chr4 47123616 N chr4 47123732 N DEL 11
SRR1766447.2263748 chr4 47123616 N chr4 47123732 N DEL 11
SRR1766478.11765584 chr7 98548087 N chr7 98548224 N DEL 7
SRR1766486.7116022 chr7 98548101 N chr7 98548218 N DEL 10
SRR1766463.2227396 chr7 98548132 N chr7 98548749 N DEL 4
SRR1766463.7919771 chr7 98548140 N chr7 98548633 N DEL 9
SRR1766451.70958 chr7 98548129 N chr7 98548218 N DEL 9
SRR1766444.1218641 chr7 98548111 N chr7 98548200 N DEL 9
SRR1766466.2612322 chr7 98548115 N chr7 98548360 N DEL 10
SRR1766460.11162023 chr7 98548043 N chr7 98548146 N DUP 10
SRR1766461.6444505 chr7 98548147 N chr7 98548220 N DEL 10
SRR1766442.13887972 chr7 98548164 N chr7 98548669 N DEL 10
SRR1766461.9124717 chr7 98548157 N chr7 98548598 N DEL 15
SRR1766486.6817236 chr7 98548163 N chr7 98548768 N DEL 14
SRR1766476.461666 chr7 98548123 N chr7 98548208 N DEL 20
SRR1766442.27465266 chr7 98548139 N chr7 98548224 N DEL 15
SRR1766448.71091 chr7 98548139 N chr7 98548224 N DEL 15
SRR1766458.9403477 chr7 98548212 N chr7 98548309 N DEL 14
SRR1766471.264531 chr7 98548043 N chr7 98548214 N DUP 5
SRR1766471.10490373 chr7 98548043 N chr7 98548234 N DUP 3
SRR1766442.5942859 chr7 98548148 N chr7 98548243 N DUP 10
SRR1766467.11806918 chr7 98548247 N chr7 98548424 N DEL 4
SRR1766477.383737 chr7 98548043 N chr7 98548242 N DUP 10
SRR1766442.38352373 chr7 98548256 N chr7 98548729 N DEL 5
SRR1766470.5566145 chr7 98548268 N chr7 98548329 N DEL 10
SRR1766483.169293 chr7 98548200 N chr7 98548703 N DUP 17
SRR1766446.9791612 chr7 98548043 N chr7 98548278 N DUP 5
SRR1766471.11487128 chr7 98548208 N chr7 98548263 N DUP 14
SRR1766467.8889349 chr7 98548239 N chr7 98548344 N DEL 6
SRR1766442.40470313 chr7 98548220 N chr7 98548283 N DUP 12
SRR1766461.8064668 chr7 98548235 N chr7 98548690 N DUP 21
SRR1766466.4977195 chr7 98548186 N chr7 98548645 N DUP 17
SRR1766471.630374 chr7 98548186 N chr7 98548645 N DUP 16
SRR1766453.720103 chr7 98548296 N chr7 98548765 N DEL 16
SRR1766463.8036211 chr7 98548267 N chr7 98548344 N DEL 18
SRR1766461.948423 chr7 98548061 N chr7 98548202 N DEL 6
SRR1766446.8319032 chr7 98548045 N chr7 98548304 N DUP 12
SRR1766470.5739754 chr7 98548317 N chr7 98548766 N DEL 9
SRR1766484.3714467 chr7 98548322 N chr7 98548771 N DEL 12
SRR1766458.1981564 chr7 98548225 N chr7 98548276 N DUP 22
SRR1766484.11219731 chr7 98548225 N chr7 98548276 N DUP 28
SRR1766453.5406955 chr7 98548221 N chr7 98548324 N DUP 10
SRR1766466.8379930 chr7 98548190 N chr7 98548301 N DUP 10
SRR1766481.6867636 chr7 98548211 N chr7 98548326 N DUP 14
SRR1766460.1941494 chr7 98548116 N chr7 98548233 N DEL 4
SRR1766486.272339 chr7 98548208 N chr7 98548347 N DUP 6
SRR1766467.6559650 chr7 98548219 N chr7 98548350 N DUP 10
SRR1766460.1941494 chr7 98548025 N chr7 98548368 N DUP 9
SRR1766485.2766451 chr7 98548043 N chr7 98548366 N DUP 8
SRR1766457.5098205 chr7 98548200 N chr7 98548335 N DUP 12
SRR1766442.38352373 chr7 98548123 N chr7 98548256 N DEL 5
SRR1766470.10609240 chr7 98548376 N chr7 98548749 N DEL 17
SRR1766462.1249024 chr7 98548200 N chr7 98548307 N DUP 22
SRR1766458.8643213 chr7 98548395 N chr7 98548756 N DEL 10
SRR1766478.10878121 chr7 98548262 N chr7 98548347 N DEL 10
SRR1766460.9077210 chr7 98548144 N chr7 98548305 N DEL 5
SRR1766449.5729004 chr7 98548412 N chr7 98548757 N DEL 5
SRR1766481.11251140 chr7 98548244 N chr7 98548309 N DEL 11
SRR1766481.4296496 chr7 98548247 N chr7 98548332 N DEL 18
SRR1766467.6559650 chr7 98548162 N chr7 98548339 N DEL 10
SRR1766448.4562121 chr7 98548200 N chr7 98548407 N DUP 18
SRR1766442.18633094 chr7 98548274 N chr7 98548461 N DUP 5
SRR1766462.5733748 chr7 98548244 N chr7 98548381 N DEL 15
SRR1766476.4413794 chr7 98548362 N chr7 98548621 N DUP 5
SRR1766486.5726415 chr7 98548358 N chr7 98548441 N DUP 15
SRR1766485.6895961 chr7 98548039 N chr7 98548372 N DEL 1
SRR1766470.10609240 chr7 98548124 N chr7 98548381 N DEL 5
SRR1766451.6047935 chr7 98548488 N chr7 98548765 N DEL 13
SRR1766476.9806805 chr7 98548085 N chr7 98548484 N DUP 14
SRR1766448.2205439 chr7 98548205 N chr7 98548394 N DEL 9
SRR1766447.1335646 chr7 98548234 N chr7 98548509 N DUP 3
SRR1766478.5194205 chr7 98548043 N chr7 98548522 N DUP 13
SRR1766442.25488686 chr7 98548420 N chr7 98548523 N DUP 12
SRR1766458.6408914 chr7 98548061 N chr7 98548418 N DEL 5
SRR1766448.2205439 chr7 98548218 N chr7 98548525 N DUP 22
SRR1766475.3967999 chr7 98548245 N chr7 98548466 N DEL 26
SRR1766471.11487128 chr7 98548239 N chr7 98548444 N DEL 5
SRR1766484.10602199 chr7 98548218 N chr7 98548545 N DUP 6
SRR1766442.6855979 chr7 98548248 N chr7 98548473 N DEL 18
SRR1766453.8594256 chr7 98548274 N chr7 98548569 N DUP 7
SRR1766452.4814280 chr7 98548245 N chr7 98548466 N DEL 15
SRR1766484.2043011 chr7 98548472 N chr7 98548583 N DUP 15
SRR1766446.9127200 chr7 98548089 N chr7 98548474 N DEL 5
SRR1766460.4659647 chr7 98548106 N chr7 98548569 N DUP 10
SRR1766477.4790412 chr7 98548274 N chr7 98548593 N DUP 5
SRR1766445.8523246 chr7 98548244 N chr7 98548485 N DEL 5
SRR1766475.10506637 chr7 98548066 N chr7 98548499 N DEL 1
SRR1766443.9934761 chr7 98548244 N chr7 98548529 N DEL 5
SRR1766453.3255258 chr7 98548244 N chr7 98548529 N DEL 5
SRR1766481.620548 chr7 98548528 N chr7 98548843 N DUP 3
SRR1766442.5346174 chr7 98548472 N chr7 98548639 N DUP 5
SRR1766452.4814280 chr7 98548086 N chr7 98548539 N DEL 2
SRR1766484.3714467 chr7 98548270 N chr7 98548645 N DUP 4
SRR1766486.8758233 chr7 98548058 N chr7 98548539 N DEL 4
SRR1766464.8484214 chr7 98548472 N chr7 98548655 N DUP 5
SRR1766471.630374 chr7 98548477 N chr7 98548546 N DEL 5
SRR1766464.7088058 chr7 98548143 N chr7 98548564 N DEL 15
SRR1766442.4903226 chr7 98548423 N chr7 98548674 N DUP 14
SRR1766442.13408210 chr7 98548472 N chr7 98548639 N DUP 3
SRR1766452.2820528 chr7 98548488 N chr7 98548557 N DEL 15
SRR1766474.4111321 chr7 98548471 N chr7 98548560 N DEL 5
SRR1766477.8484845 chr7 98548043 N chr7 98548678 N DUP 7
SRR1766442.13408210 chr7 98548242 N chr7 98548571 N DEL 1
SRR1766466.4977195 chr7 98548282 N chr7 98548659 N DEL 7
SRR1766476.7130305 chr7 98548240 N chr7 98548589 N DEL 15
SRR1766462.7628201 chr7 98548106 N chr7 98548701 N DUP 10
SRR1766453.3469609 chr7 98548144 N chr7 98548627 N DUP 12
SRR1766452.3016551 chr7 98548186 N chr7 98548645 N DUP 31
SRR1766442.7191805 chr7 98548235 N chr7 98548690 N DUP 29
SRR1766482.8653878 chr7 98548245 N chr7 98548618 N DEL 5
SRR1766442.2809209 chr7 98548058 N chr7 98548619 N DEL 5
SRR1766477.9096937 chr7 98548376 N chr7 98548637 N DEL 5
SRR1766461.3998588 chr7 98548259 N chr7 98548640 N DEL 5
SRR1766453.3541418 chr7 98548100 N chr7 98548641 N DEL 6
SRR1766443.5165035 chr7 98548124 N chr7 98548669 N DEL 10
SRR1766449.5729004 chr7 98548121 N chr7 98548666 N DEL 2
SRR1766442.1388390 chr7 98548618 N chr7 98548711 N DEL 6
SRR1766486.6420781 chr7 98548086 N chr7 98548711 N DEL 6
SRR1766442.40470313 chr7 98548624 N chr7 98548749 N DEL 5
SRR1766450.673205 chr7 98548103 N chr7 98548876 N DEL 1
SRR1766479.1981210 chr20 33115619 N chr20 33115892 N DEL 1
SRR1766467.2633332 chr20 33115621 N chr20 33115817 N DEL 1
SRR1766445.4953721 chr20 33115533 N chr20 33116055 N DUP 5
SRR1766471.4531305 chr20 33115591 N chr20 33115822 N DUP 5
SRR1766483.3740123 chr20 33115683 N chr20 33115797 N DUP 3
SRR1766485.4716558 chr20 33115584 N chr20 33115740 N DEL 10
SRR1766444.428024 chr9 91132870 N chr9 91132999 N DEL 1
SRR1766475.10822230 chr8 72573730 N chr8 72573891 N DEL 5
SRR1766482.2577613 chr8 72573698 N chr8 72573779 N DEL 5
SRR1766472.1075631 chr8 72573698 N chr8 72573859 N DEL 15
SRR1766450.9008725 chr8 72573769 N chr8 72573890 N DEL 5
SRR1766451.290563 chr8 72573769 N chr8 72573890 N DEL 6
SRR1766450.4950739 chr8 72573821 N chr8 72573940 N DUP 5
SRR1766464.5436726 chr8 72573685 N chr8 72573964 N DUP 2
SRR1766468.5766139 chr8 72573821 N chr8 72573940 N DUP 5
SRR1766460.9278687 chr8 72573698 N chr8 72573939 N DEL 5
SRR1766477.8794052 chr10 123068735 N chr10 123068804 N DEL 2
SRR1766479.11684919 chr10 123068735 N chr10 123068804 N DEL 2
SRR1766485.11987279 chr10 123068733 N chr10 123068802 N DEL 4
SRR1766484.4937537 chr10 30500008 N chr10 30500276 N DEL 5
SRR1766458.4594203 chr19 51944740 N chr19 51944993 N DEL 15
SRR1766442.27426434 chr19 51944760 N chr19 51945013 N DEL 5
SRR1766468.783762 chr19 51944794 N chr19 51945047 N DEL 9
SRR1766476.5224973 chr19 51944879 N chr19 51945130 N DUP 5
SRR1766480.6838663 chr19 51944794 N chr19 51945047 N DEL 18
SRR1766466.2797376 chr19 51944903 N chr19 51945156 N DEL 25
SRR1766464.2882461 chr11 129671491 N chr11 129671694 N DUP 5
SRR1766466.8807604 chr11 129671511 N chr11 129671713 N DEL 5
SRR1766442.4047295 chr11 129671829 N chr11 129672176 N DEL 16
SRR1766462.7016405 chr11 129671834 N chr11 129672181 N DEL 10
SRR1766477.8915645 chr11 129671835 N chr11 129672182 N DEL 9
SRR1766474.2884312 chr11 129671831 N chr11 129672259 N DEL 6
SRR1766450.10255368 chr11 129671835 N chr11 129672263 N DEL 2
SRR1766482.8707106 chr11 129671832 N chr11 129672260 N DEL 5
SRR1766462.4809574 chr3 122252489 N chr3 122252560 N DEL 10
SRR1766469.10628670 chr3 122252509 N chr3 122252572 N DEL 2
SRR1766484.2031519 chr1 203500084 N chr1 203500341 N DEL 9
SRR1766471.7217889 chr3 47659267 N chr3 47659431 N DUP 5
SRR1766473.3170980 chr6 59360905 N chr6 59361226 N DEL 5
SRR1766485.9605830 chr6 59360896 N chr6 59361217 N DEL 20
SRR1766455.9178962 chr6 59360842 N chr6 59361010 N DUP 1
SRR1766457.6889164 chr6 59360836 N chr6 59361004 N DUP 10
SRR1766453.4173298 chr6 59360818 N chr6 59360986 N DUP 10
SRR1766457.483625 chr8 144670308 N chr8 144670381 N DUP 5
SRR1766442.21498640 chr11 131265291 N chr11 131265465 N DEL 15
SRR1766472.10859752 chr11 131265291 N chr11 131265465 N DEL 15
SRR1766451.10489424 chr11 131265291 N chr11 131265465 N DEL 16
SRR1766442.15356765 chr11 131265291 N chr11 131265465 N DEL 17
SRR1766465.2138958 chr11 131265291 N chr11 131265465 N DEL 17
SRR1766442.861060 chr11 131265291 N chr11 131265465 N DEL 17
SRR1766484.9393062 chr11 131265291 N chr11 131265465 N DEL 22
SRR1766442.22279736 chr11 131265291 N chr11 131265465 N DEL 24
SRR1766448.674019 chr11 131265291 N chr11 131265465 N DEL 24
SRR1766476.7224224 chr11 131265291 N chr11 131265465 N DEL 24
SRR1766485.10255151 chr11 131265325 N chr11 131265447 N DEL 30
SRR1766445.8661391 chr11 131265291 N chr11 131265465 N DEL 26
SRR1766458.1558429 chr11 131265291 N chr11 131265465 N DEL 26
SRR1766475.1156443 chr11 131265325 N chr11 131265447 N DEL 30
SRR1766448.6456425 chr11 131265325 N chr11 131265447 N DEL 30
SRR1766451.9100705 chr11 131265291 N chr11 131265465 N DEL 26
SRR1766485.9338154 chr11 131265291 N chr11 131265465 N DEL 26
SRR1766479.3546291 chr11 131265325 N chr11 131265447 N DEL 30
SRR1766467.219304 chr11 131265291 N chr11 131265465 N DEL 30
SRR1766454.2075922 chr11 131265284 N chr11 131265474 N DUP 4
SRR1766463.6385019 chr11 131265284 N chr11 131265474 N DUP 4
SRR1766479.13508971 chr11 131265284 N chr11 131265474 N DUP 4
SRR1766453.4034834 chr11 131265284 N chr11 131265474 N DUP 4
SRR1766477.3862137 chr11 131265284 N chr11 131265474 N DUP 4
SRR1766442.22279736 chr11 131265284 N chr11 131265474 N DUP 4
SRR1766446.7220201 chr11 131265284 N chr11 131265474 N DUP 4
SRR1766463.2421801 chr11 131265285 N chr11 131265475 N DUP 4
SRR1766459.6349939 chr11 131265287 N chr11 131265477 N DUP 2
SRR1766457.8210272 chr11 131265287 N chr11 131265477 N DUP 2
SRR1766451.4150346 chr11 131265352 N chr11 131265544 N DUP 21
SRR1766460.4871000 chr11 131265296 N chr11 131265357 N DEL 5
SRR1766467.5413266 chr11 131265368 N chr11 131265417 N DUP 11
SRR1766481.234453 chr11 131265352 N chr11 131265544 N DUP 11
SRR1766476.8218203 chr12 56557901 N chr12 56558202 N DUP 5
SRR1766481.11764772 chr12 56558030 N chr12 56558340 N DEL 5
SRR1766455.6746793 chr12 56558084 N chr12 56558393 N DUP 5
SRR1766472.2922658 chr4 15733379 N chr4 15733487 N DEL 5
SRR1766464.7571813 chr4 15733379 N chr4 15733487 N DEL 5
SRR1766466.445776 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766448.6861360 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766486.7403981 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766460.564753 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766456.6360332 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766466.2773231 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766459.6392920 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766442.43738583 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766478.9858646 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766464.4197082 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766447.7273899 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766467.7352371 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766465.1277132 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766482.13002681 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766459.4540238 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766476.10930185 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766485.7572244 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766462.3912399 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766442.33411782 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766466.9910422 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766468.2612794 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766445.1267 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766450.9650909 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766442.5546913 chr4 15733430 N chr4 15733538 N DEL 5
SRR1766470.9197282 chr4 15733452 N chr4 15733558 N DUP 5
SRR1766473.5689533 chr4 15733452 N chr4 15733558 N DUP 5
SRR1766444.5294263 chr4 15733454 N chr4 15733560 N DUP 3
SRR1766475.3597832 chr4 15733442 N chr4 15733548 N DUP 2
SRR1766474.3008217 chr4 15733484 N chr4 15733631 N DUP 5
SRR1766481.3520101 chr4 15733484 N chr4 15733631 N DUP 5
SRR1766485.8934153 chr4 15733484 N chr4 15733631 N DUP 5
SRR1766468.2007970 chr4 15733383 N chr4 15733532 N DEL 18
SRR1766481.12862453 chr4 15733484 N chr4 15733631 N DUP 5
SRR1766461.3951074 chr4 15733525 N chr4 15733633 N DEL 5
SRR1766467.7869835 chr4 15733525 N chr4 15733633 N DEL 5
SRR1766472.2922658 chr4 15733525 N chr4 15733633 N DEL 5
SRR1766483.10835780 chr4 15733525 N chr4 15733633 N DEL 5
SRR1766452.4088085 chr4 15733525 N chr4 15733633 N DEL 5
SRR1766447.8959949 chr4 15733525 N chr4 15733633 N DEL 5
SRR1766444.5486946 chr4 15733525 N chr4 15733633 N DEL 5
SRR1766472.7210017 chr4 15733525 N chr4 15733633 N DEL 5
SRR1766485.7649150 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766482.2902224 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766442.43743060 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766443.5310923 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766457.5709426 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766485.376141 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766454.7804134 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766475.1437449 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766442.28706715 chr4 15733418 N chr4 15733633 N DEL 5
SRR1766442.40611382 chr4 15733378 N chr4 15733634 N DEL 5
SRR1766468.2612794 chr4 15733378 N chr4 15733634 N DEL 5
SRR1766475.536004 chr4 15733420 N chr4 15733635 N DEL 5
SRR1766486.7403981 chr4 15733421 N chr4 15733636 N DEL 5
SRR1766464.8478121 chr4 15733498 N chr4 15733647 N DEL 1
SRR1766461.3839406 chr4 144058388 N chr4 144058472 N DUP 3
SRR1766482.8795333 chr4 144058388 N chr4 144058472 N DUP 5
SRR1766453.1964387 chr4 144058404 N chr4 144058502 N DEL 9
SRR1766448.9924526 chr4 144058406 N chr4 144058504 N DEL 7
SRR1766460.4593620 chr11 70119172 N chr11 70119469 N DUP 1
SRR1766482.1129829 chr11 70119213 N chr11 70119510 N DUP 5
SRR1766442.42863461 chr11 70119163 N chr11 70119388 N DUP 10
SRR1766474.8467699 chr11 70119427 N chr11 70119627 N DEL 5
SRR1766483.7050024 chr11 70119432 N chr11 70119632 N DEL 10
SRR1766472.8823127 chr11 70119320 N chr11 70119455 N DUP 5
SRR1766482.8676524 chr11 70119386 N chr11 70119521 N DUP 5
SRR1766442.27729275 chr11 70119350 N chr11 70119487 N DEL 3
SRR1766479.11067805 chr7 50459509 N chr7 50459780 N DUP 8
SRR1766476.7916920 chr7 50459756 N chr7 50459872 N DUP 5
SRR1766476.5278659 chr7 50459692 N chr7 50459884 N DUP 2
SRR1766486.4582198 chr7 50459932 N chr7 50460030 N DEL 5
SRR1766454.6137843 chr7 50459722 N chr7 50459916 N DEL 10
SRR1766478.10207624 chr15 58282915 N chr15 58282972 N DEL 8
SRR1766480.8791773 chr15 58282915 N chr15 58282972 N DEL 8
SRR1766480.1118635 chr2 16332758 N chr2 16332887 N DEL 5
SRR1766461.2220115 chr21 43160144 N chr21 43160222 N DUP 2
SRR1766442.2124340 chr21 43160258 N chr21 43160398 N DEL 5
SRR1766467.6930519 chr21 43160399 N chr21 43160463 N DEL 1
SRR1766456.6474595 chr21 43160576 N chr21 43160659 N DEL 1
SRR1766449.557086 chr21 43160468 N chr21 43160771 N DUP 5
SRR1766483.7554626 chr21 43160012 N chr21 43160686 N DEL 5
SRR1766481.6269075 chr21 43160620 N chr21 43160701 N DEL 5
SRR1766467.9106630 chrX 120374689 N chrX 120374755 N DUP 7
SRR1766459.3422271 chrX 120374689 N chrX 120374755 N DUP 7
SRR1766481.2162972 chrX 120374757 N chrX 120374845 N DEL 17
SRR1766458.6409505 chrX 120374674 N chrX 120374858 N DUP 9
SRR1766485.3273815 chrX 120374817 N chrX 120374925 N DUP 3
SRR1766465.10776256 chrX 120374820 N chrX 120374928 N DUP 2
SRR1766458.2264043 chrX 120374820 N chrX 120374928 N DUP 4
SRR1766446.9985693 chrX 120374820 N chrX 120374928 N DUP 6
SRR1766452.107015 chrX 120374810 N chrX 120374920 N DUP 15
SRR1766451.294699 chrX 120374788 N chrX 120374910 N DUP 16
SRR1766457.1377531 chrX 120374719 N chrX 120374907 N DEL 2
SRR1766471.8831086 chrX 120374719 N chrX 120374907 N DEL 7
SRR1766446.10099312 chrX 120374696 N chrX 120374907 N DEL 7
SRR1766485.4373049 chrX 120374696 N chrX 120374907 N DEL 16
SRR1766486.10324246 chr10 124306160 N chr10 124306300 N DUP 3
SRR1766450.7704233 chr10 124306160 N chr10 124306300 N DUP 5
SRR1766450.7380979 chr10 124306167 N chr10 124306307 N DUP 5
SRR1766445.39710 chr11 48956125 N chr11 48956242 N DEL 3
SRR1766453.3189876 chr11 48956132 N chr11 48956210 N DEL 4
SRR1766486.431758 chr11 2773264 N chr11 2773409 N DUP 2
SRR1766468.5013654 chr11 2773499 N chr11 2773638 N DUP 6
SRR1766470.7999481 chrX 54065527 N chrX 54065825 N DEL 2
SRR1766450.10847777 chrX 54065345 N chrX 54065860 N DEL 10
SRR1766466.6724924 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766483.8471184 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766484.10564141 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766454.8744575 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766468.1924063 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766485.4868547 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766442.11627177 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766447.4222320 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766484.9696450 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766465.1980891 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766475.6264890 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766475.9555954 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766461.6343354 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766442.27421955 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766484.12055572 chr1 162727366 N chr1 162727421 N DEL 5
SRR1766445.8753351 chr1 162727339 N chr1 162727421 N DEL 5
SRR1766450.8234669 chr1 162727339 N chr1 162727421 N DEL 5
SRR1766442.47343 chr1 162727339 N chr1 162727421 N DEL 5
SRR1766469.97096 chr1 162727339 N chr1 162727421 N DEL 5
SRR1766486.9621019 chr1 162727339 N chr1 162727421 N DEL 5
SRR1766462.7927521 chr1 162727339 N chr1 162727421 N DEL 5
SRR1766455.4439218 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766479.4388881 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766443.10354262 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766486.7199176 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766466.7073609 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766455.4791355 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766475.10743860 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766465.8455944 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766471.8115941 chr1 162727312 N chr1 162727421 N DEL 5
SRR1766480.7687492 chr10 87320563 N chr10 87320674 N DUP 1
SRR1766481.4209142 chr10 87320617 N chr10 87320730 N DEL 4
SRR1766466.4449911 chr7 155958254 N chr7 155958375 N DEL 5
SRR1766442.29239577 chr7 155958259 N chr7 155958380 N DEL 5
SRR1766444.5968899 chr7 155958165 N chr7 155958286 N DEL 1
SRR1766473.11385992 chr4 160662794 N chr4 160662928 N DEL 5
SRR1766482.5014329 chr4 160662812 N chr4 160662944 N DUP 5
SRR1766462.9581166 chr20 36976591 N chr20 36976765 N DUP 9
SRR1766472.6244029 chr20 36976590 N chr20 36976969 N DUP 6
SRR1766447.4140266 chr20 36976587 N chr20 36976712 N DUP 3
SRR1766482.5320126 chr20 36976587 N chr20 36976712 N DUP 6
SRR1766445.4310590 chr20 36976713 N chr20 36976966 N DUP 6
SRR1766459.7653812 chr20 36976537 N chr20 36976713 N DEL 6
SRR1766454.7343632 chr20 36976600 N chr20 36976727 N DEL 1
SRR1766466.7316142 chr20 36976600 N chr20 36976727 N DEL 1
SRR1766484.7672051 chr20 36976512 N chr20 36976860 N DUP 12
SRR1766442.33669736 chr20 36976713 N chr20 36976839 N DUP 5
SRR1766447.1968733 chr20 36976512 N chr20 36976860 N DUP 12
SRR1766457.807368 chr20 36976703 N chr20 36976831 N DEL 5
SRR1766475.10176252 chr20 36976713 N chr20 36976839 N DUP 5
SRR1766457.6491588 chr20 36976713 N chr20 36976839 N DUP 5
SRR1766472.3416332 chr20 36976713 N chr20 36976839 N DUP 5
SRR1766464.1302046 chr20 36976713 N chr20 36976839 N DUP 5
SRR1766485.4660086 chr20 36976713 N chr20 36976839 N DUP 5
SRR1766446.878032 chr20 36976713 N chr20 36976839 N DUP 5
SRR1766465.1364111 chr8 38508022 N chr8 38508089 N DEL 8
SRR1766458.2008137 chr8 38508022 N chr8 38508089 N DEL 9
SRR1766482.5858890 chr8 38508022 N chr8 38508089 N DEL 9
SRR1766478.660096 chr8 38508022 N chr8 38508089 N DEL 9
SRR1766473.4263025 chr8 38508022 N chr8 38508089 N DEL 12
SRR1766469.6961169 chr8 38508008 N chr8 38508090 N DEL 14
SRR1766486.9922501 chr17 72189556 N chr17 72189693 N DUP 3
SRR1766449.8636484 chr17 72189542 N chr17 72189697 N DUP 14
SRR1766472.2440465 chr9 43337167 N chr9 43337241 N DUP 12
SRR1766442.45733144 chr9 43337177 N chr9 43337300 N DUP 2
SRR1766450.8914783 chr9 43337194 N chr9 43337343 N DUP 3
SRR1766484.6622019 chr9 43337185 N chr9 43337334 N DUP 5
SRR1766474.6441472 chr9 43337185 N chr9 43337334 N DUP 5
SRR1766442.41433694 chr9 43337321 N chr9 43337397 N DEL 7
SRR1766459.11224855 chr9 43337229 N chr9 43337329 N DUP 3
SRR1766476.1772692 chr9 43337254 N chr9 43337328 N DUP 5
SRR1766460.1570980 chr9 43337254 N chr9 43337328 N DUP 5
SRR1766454.3094938 chr9 43337254 N chr9 43337328 N DUP 5
SRR1766462.4458553 chr9 43337254 N chr9 43337328 N DUP 5
SRR1766451.7594565 chr9 43337221 N chr9 43337396 N DUP 5
SRR1766442.21596347 chr9 43337221 N chr9 43337396 N DUP 8
SRR1766442.11017443 chr9 43337225 N chr9 43337400 N DUP 8
SRR1766447.2529256 chr17 73696955 N chr17 73697214 N DEL 3
SRR1766460.4041490 chr17 73697027 N chr17 73697110 N DUP 5
SRR1766449.3071390 chr17 73697028 N chr17 73697265 N DUP 4
SRR1766459.3573798 chr17 73697006 N chr17 73697174 N DUP 2
SRR1766445.1287922 chr17 73697114 N chr17 73697242 N DUP 5
SRR1766478.9649410 chr17 73697132 N chr17 73697218 N DEL 8
SRR1766460.6991982 chr17 73697164 N chr17 73697252 N DUP 3
SRR1766458.185366 chr17 73697033 N chr17 73697203 N DEL 5
SRR1766462.9722638 chr17 73697033 N chr17 73697203 N DEL 5
SRR1766477.4892721 chr17 73696967 N chr17 73697226 N DEL 3
SRR1766484.6706550 chr1 211219273 N chr1 211219417 N DUP 3
SRR1766482.12321221 chr5 280627 N chr5 280835 N DEL 5
SRR1766464.8222280 chr5 280668 N chr5 280952 N DEL 5
SRR1766466.292360 chr8 142205166 N chr8 142205237 N DEL 22
SRR1766453.4094 chr8 142205162 N chr8 142205229 N DEL 9
SRR1766486.4109640 chr8 142205162 N chr8 142205229 N DEL 9
SRR1766445.5686130 chr8 142205162 N chr8 142205229 N DEL 9
SRR1766442.20093800 chr8 142205162 N chr8 142205229 N DEL 9
SRR1766453.1741952 chr8 142205162 N chr8 142205229 N DEL 9
SRR1766466.2479373 chr6 157870670 N chr6 157870732 N DEL 5
SRR1766450.2426774 chr6 157870670 N chr6 157870940 N DEL 5
SRR1766442.15755755 chr6 157870686 N chr6 157870748 N DUP 8
SRR1766462.7000411 chr6 157870704 N chr6 157870913 N DEL 5
SRR1766460.5617959 chr6 157870610 N chr6 157870819 N DUP 10
SRR1766455.7348910 chr19 5774621 N chr19 5774946 N DEL 5
SRR1766467.7354583 chr19 5774672 N chr19 5775001 N DEL 2
SRR1766474.5561374 chr1 91140860 N chr1 91140915 N DUP 2
SRR1766474.2905388 chr12 31610114 N chr12 31610430 N DEL 5
SRR1766442.45318606 chrX 20559277 N chrX 20559598 N DEL 6
SRR1766466.6142338 chr10 27296559 N chr10 27296783 N DUP 15
SRR1766451.8314679 chr10 27296547 N chr10 27296722 N DUP 5
SRR1766476.10091523 chr10 27296590 N chr10 27296716 N DUP 10
SRR1766469.10364748 chr10 27296591 N chr10 27296768 N DEL 5
SRR1766471.10382996 chr8 26128390 N chr8 26128447 N DEL 2
SRR1766442.1572658 chr8 26128485 N chr8 26128538 N DEL 5
SRR1766460.1123600 chr8 26128358 N chr8 26128540 N DEL 5
SRR1766482.5402242 chr8 26128358 N chr8 26128540 N DEL 5
SRR1766467.9535631 chr12 34437113 N chr12 34437455 N DEL 2
SRR1766482.980916 chr4 43451137 N chr4 43451231 N DEL 14
SRR1766442.27703620 chr4 43450920 N chr4 43451088 N DEL 10
SRR1766476.535031 chr4 43451137 N chr4 43451231 N DEL 34
SRR1766453.5121668 chr4 43451137 N chr4 43451231 N DEL 42
SRR1766466.2585089 chr4 43451137 N chr4 43451231 N DEL 46
SRR1766481.4666068 chr4 43451137 N chr4 43451231 N DEL 46
SRR1766446.10223277 chr4 43451144 N chr4 43451238 N DEL 8
SRR1766477.11559707 chr4 43451144 N chr4 43451238 N DEL 8
SRR1766459.9894578 chr4 43452278 N chr4 43452343 N DEL 5
SRR1766464.783418 chr4 43452278 N chr4 43452343 N DEL 5
SRR1766463.8449283 chr4 43452150 N chr4 43452363 N DEL 3
SRR1766453.1432334 chr4 43452574 N chr4 43452653 N DUP 5
SRR1766470.1922316 chr4 43452574 N chr4 43452653 N DUP 5
SRR1766453.3537969 chr4 43452503 N chr4 43452668 N DUP 5
SRR1766457.7065825 chr4 43452503 N chr4 43452668 N DUP 5
SRR1766442.44638811 chr4 43452593 N chr4 43452674 N DEL 5
SRR1766453.9828256 chr21 46109188 N chr21 46109260 N DEL 5
SRR1766468.6833304 chr9 134115812 N chr9 134115989 N DEL 5
SRR1766484.8998653 chr9 134115720 N chr9 134115895 N DUP 5
SRR1766442.13103493 chr9 134115744 N chr9 134115921 N DEL 5
SRR1766443.6423881 chr9 134115757 N chr9 134115934 N DEL 5
SRR1766469.1730906 chr9 134115789 N chr9 134115968 N DEL 7
SRR1766486.6267016 chr10 123572702 N chr10 123572872 N DEL 3
SRR1766452.6849372 chr10 12345317 N chr10 12345646 N DUP 1
SRR1766465.10137073 chr10 12345347 N chr10 12345513 N DUP 6
SRR1766462.11108636 chr6 22836799 N chr6 22836928 N DEL 5
SRR1766477.221440 chr6 22836800 N chr6 22836929 N DEL 2
SRR1766483.11233226 chr6 22836813 N chr6 22836942 N DEL 5
SRR1766442.43901911 chr6 22836799 N chr6 22836928 N DEL 10
SRR1766443.5421022 chr6 22836800 N chr6 22836929 N DEL 5
SRR1766461.1534938 chr6 22836949 N chr6 22837204 N DEL 6
SRR1766451.2477563 chr6 22836918 N chr6 22837221 N DUP 5
SRR1766457.769618 chr6 22836727 N chr6 22837030 N DUP 10
SRR1766474.6762309 chr6 22836737 N chr6 22837089 N DUP 10
SRR1766482.12278866 chr6 22836769 N chr6 22837121 N DUP 1
SRR1766483.6957947 chr6 22836780 N chr6 22837036 N DEL 3
SRR1766447.1367030 chr6 22836753 N chr6 22837058 N DEL 9
SRR1766469.7077818 chr9 43321680 N chr9 43321829 N DUP 5
SRR1766443.4923669 chr9 43321687 N chr9 43321784 N DUP 5
SRR1766468.2838446 chr9 43321797 N chr9 43321850 N DEL 5
SRR1766445.9010177 chr9 43321797 N chr9 43321850 N DEL 6
SRR1766458.8358781 chr9 43321797 N chr9 43321850 N DEL 9
SRR1766464.6026045 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766460.1982169 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766453.7066482 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766442.12203348 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766451.6880040 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766447.2945355 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766453.6237945 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766450.1838200 chr9 43321797 N chr9 43321850 N DEL 10
SRR1766460.8339405 chr9 43321830 N chr9 43321923 N DUP 14
SRR1766445.8712223 chr9 43321647 N chr9 43321900 N DUP 5
SRR1766455.7921756 chr9 43321921 N chr9 43321974 N DEL 2
SRR1766448.7581432 chr9 43321731 N chr9 43321807 N DEL 5
SRR1766472.5866829 chr9 43321846 N chr9 43321897 N DUP 10
SRR1766483.669286 chr9 43321798 N chr9 43321849 N DUP 11
SRR1766470.2513747 chr9 43321843 N chr9 43321894 N DUP 11
SRR1766453.5350190 chr9 43321843 N chr9 43321894 N DUP 12
SRR1766484.5894344 chr9 43321779 N chr9 43321858 N DEL 5
SRR1766474.7568818 chr9 43321655 N chr9 43322058 N DUP 6
SRR1766473.5193450 chr9 43321842 N chr9 43322069 N DUP 4
SRR1766448.1113246 chr1 2960156 N chr1 2960247 N DEL 5
SRR1766445.9477328 chr1 2960163 N chr1 2960254 N DEL 5
SRR1766456.3931677 chr1 2960156 N chr1 2960247 N DEL 8
SRR1766452.7524072 chr1 2960156 N chr1 2960247 N DEL 10
SRR1766471.10812301 chr1 2960156 N chr1 2960247 N DEL 10
SRR1766465.1854512 chr1 2960156 N chr1 2960277 N DEL 12
SRR1766482.4026133 chr1 2960156 N chr1 2960277 N DEL 12
SRR1766443.1192417 chr1 2960156 N chr1 2960277 N DEL 13
SRR1766470.8564719 chr1 2960156 N chr1 2960277 N DEL 15
SRR1766479.9203261 chr1 2960156 N chr1 2960277 N DEL 15
SRR1766479.10388521 chr1 2960156 N chr1 2960277 N DEL 25
SRR1766461.7065754 chr1 2960162 N chr1 2960283 N DEL 5
SRR1766466.6253184 chr1 2960156 N chr1 2960277 N DEL 14
SRR1766458.7832198 chr1 2960163 N chr1 2960284 N DEL 5
SRR1766457.4757990 chr22 43737678 N chr22 43737799 N DUP 1
SRR1766457.6778094 chr22 43737664 N chr22 43737785 N DUP 5
SRR1766467.3828753 chr22 43737704 N chr22 43737825 N DUP 5
SRR1766473.7675464 chr22 43737704 N chr22 43737825 N DUP 5
SRR1766479.1652201 chr22 43737705 N chr22 43737826 N DUP 5
SRR1766477.1251589 chr22 43737706 N chr22 43737827 N DUP 5
SRR1766445.4621908 chr22 43737706 N chr22 43737827 N DUP 5
SRR1766477.5863205 chr22 43737707 N chr22 43737828 N DUP 5
SRR1766475.7133176 chr22 43737707 N chr22 43737828 N DUP 3
SRR1766481.11036162 chr22 43737843 N chr22 43737932 N DEL 5
SRR1766482.7198718 chr22 43737807 N chr22 43737918 N DUP 3
SRR1766467.2129123 chr2 3844442 N chr2 3844561 N DUP 5
SRR1766468.3661359 chr2 3844467 N chr2 3844526 N DUP 10
SRR1766469.4306334 chr2 3844488 N chr2 3844609 N DEL 5
SRR1766464.8546167 chr2 3844492 N chr2 3844613 N DEL 5
SRR1766454.10290652 chr2 3844489 N chr2 3844610 N DEL 5
SRR1766442.25242889 chr2 3844490 N chr2 3844611 N DEL 5
SRR1766484.523673 chr2 3844490 N chr2 3844611 N DEL 5
SRR1766485.958744 chrX 56725954 N chrX 56726025 N DEL 1
SRR1766478.10911501 chr17 51613716 N chr17 51613769 N DEL 5
SRR1766462.8979372 chr12 96104146 N chr12 96104247 N DEL 5
SRR1766452.5653115 chr1 38647379 N chr1 38647496 N DEL 6
SRR1766445.8725304 chr1 38647548 N chr1 38647623 N DUP 3
SRR1766480.8203682 chr1 38647375 N chr1 38647648 N DEL 5
SRR1766453.829135 chr10 42171825 N chr10 42171966 N DEL 10
SRR1766458.6292032 chr10 42171772 N chr10 42171883 N DUP 5
SRR1766475.5093522 chr10 42171772 N chr10 42171883 N DUP 5
SRR1766482.13089722 chr10 42171756 N chr10 42171919 N DUP 7
SRR1766459.4761453 chr10 42171756 N chr10 42171919 N DUP 8
SRR1766458.4299740 chr10 42171701 N chr10 42171840 N DEL 5
SRR1766470.5077822 chr10 42171845 N chr10 42171945 N DUP 3
SRR1766471.2631426 chr10 42171704 N chr10 42171843 N DEL 2
SRR1766448.6758659 chr10 42171865 N chr10 42171965 N DUP 6
SRR1766478.2377712 chr10 42171865 N chr10 42171965 N DUP 6
SRR1766458.8630276 chr10 42171865 N chr10 42171965 N DUP 7
SRR1766480.7533387 chrX 146259472 N chrX 146259617 N DEL 3
SRR1766472.11835266 chr11 62962001 N chr11 62962302 N DEL 19
SRR1766442.27904954 chr11 62962139 N chr11 62962440 N DEL 5
SRR1766442.6779404 chr11 62962001 N chr11 62962302 N DEL 10
SRR1766478.10273516 chr11 62962263 N chr11 62962575 N DEL 5
SRR1766478.3257918 chr6 4895431 N chr6 4895506 N DUP 16
SRR1766479.11434772 chr6 4895448 N chr6 4895611 N DUP 5
SRR1766471.2626782 chr6 4895499 N chr6 4895610 N DUP 5
SRR1766442.26579387 chr6 4895507 N chr6 4895622 N DEL 21
SRR1766442.22697217 chr6 4895555 N chr6 4895650 N DEL 4
SRR1766448.1234984 chr16 29060373 N chr16 29060424 N DEL 3
SRR1766442.26160586 chr16 29060308 N chr16 29060408 N DEL 5
SRR1766448.9962561 chr20 63871409 N chr20 63872001 N DEL 5
SRR1766444.1029360 chr20 63871760 N chr20 63872045 N DEL 32
SRR1766485.5298360 chr15 57075906 N chr15 57075980 N DUP 8
SRR1766462.885501 chr15 57075906 N chr15 57075980 N DUP 12
SRR1766474.4160485 chr15 57075906 N chr15 57075980 N DUP 12
SRR1766471.436829 chr15 57075906 N chr15 57075980 N DUP 13
SRR1766453.7001851 chr15 57075920 N chr15 57075992 N DUP 7
SRR1766474.9860200 chr15 57075924 N chr15 57075986 N DEL 14
SRR1766443.11231260 chr12 102973626 N chr12 102973859 N DUP 5
SRR1766476.1474661 chr3 21496582 N chr3 21496653 N DUP 1
SRR1766457.7847837 chr3 21496610 N chr3 21496685 N DEL 1
SRR1766457.7035441 chr3 21496544 N chr3 21496725 N DEL 9
SRR1766474.2533292 chr3 21496544 N chr3 21496725 N DEL 9
SRR1766472.11926361 chr3 21496544 N chr3 21496725 N DEL 9
SRR1766474.4584722 chr3 21496544 N chr3 21496725 N DEL 9
SRR1766469.3164683 chr3 21496544 N chr3 21496725 N DEL 9
SRR1766449.874617 chr3 21496544 N chr3 21496725 N DEL 9
SRR1766455.4983306 chr3 21496544 N chr3 21496725 N DEL 9
SRR1766451.1556417 chr3 21496544 N chr3 21496725 N DEL 9
SRR1766459.5590550 chr3 21496547 N chr3 21496728 N DEL 9
SRR1766483.494712 chr3 21496517 N chr3 21496730 N DEL 9
SRR1766486.4078943 chr3 21496622 N chr3 21496731 N DEL 9
SRR1766442.18690879 chr2 197473575 N chr2 197473658 N DEL 7
SRR1766476.806376 chr2 197473565 N chr2 197473642 N DUP 15
SRR1766457.6012039 chr6 170251963 N chr6 170252020 N DEL 2
SRR1766482.1419644 chr6 170251963 N chr6 170252020 N DEL 2
SRR1766453.7302443 chr6 170251963 N chr6 170252020 N DEL 3
SRR1766482.4756693 chr6 170251963 N chr6 170252020 N DEL 4
SRR1766465.6486597 chr6 170251963 N chr6 170252020 N DEL 5
SRR1766486.5541864 chr6 170251963 N chr6 170252020 N DEL 5
SRR1766465.2074941 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766474.847146 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766466.5773802 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766463.7230179 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766442.42341384 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766448.10181389 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766463.8311409 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766463.3368607 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766448.3603024 chr6 170251952 N chr6 170252007 N DUP 5
SRR1766463.3368607 chr6 170252020 N chr6 170252075 N DUP 5
SRR1766442.37142560 chr6 170252020 N chr6 170252075 N DUP 5
SRR1766470.10813181 chr6 170252020 N chr6 170252075 N DUP 5
SRR1766465.9070294 chr6 170252020 N chr6 170252075 N DUP 5
SRR1766452.4274191 chr6 170252020 N chr6 170252075 N DUP 5
SRR1766457.2986462 chr6 170252020 N chr6 170252075 N DUP 5
SRR1766457.7833498 chr6 170252020 N chr6 170252075 N DUP 5
SRR1766469.2047695 chr6 170251971 N chr6 170252028 N DEL 5
SRR1766478.8840627 chr6 170251977 N chr6 170252034 N DEL 1
SRR1766454.6495806 chr1 167506388 N chr1 167506459 N DEL 7
SRR1766476.8026585 chr1 167506384 N chr1 167506439 N DEL 7
SRR1766476.3939194 chr1 167506387 N chr1 167506442 N DEL 7
SRR1766469.7847890 chr1 167506384 N chr1 167506444 N DEL 7
SRR1766453.3874319 chr1 167506388 N chr1 167506448 N DEL 6
SRR1766452.8553403 chr1 167506387 N chr1 167506452 N DEL 2
SRR1766460.7446245 chr2 225783180 N chr2 225783338 N DEL 5
SRR1766477.7574171 chr2 225783280 N chr2 225783342 N DEL 5
SRR1766443.9604506 chr19 44730626 N chr19 44730949 N DEL 5
SRR1766446.7033783 chr19 44730626 N chr19 44730949 N DEL 7
SRR1766446.7033783 chr19 44730860 N chr19 44731163 N DUP 1
SRR1766481.2334976 chr19 44730636 N chr19 44730959 N DEL 5
SRR1766458.2870641 chr19 44730669 N chr19 44730992 N DEL 5
SRR1766484.9451400 chr19 44730682 N chr19 44731005 N DEL 5
SRR1766484.9790583 chr19 44730507 N chr19 44731134 N DUP 2
SRR1766450.2365068 chr19 44730710 N chr19 44731033 N DEL 5
SRR1766445.5323279 chr19 44730723 N chr19 44731046 N DEL 5
SRR1766452.285581 chr5 38862305 N chr5 38862663 N DUP 1
SRR1766463.5115647 chr5 38862255 N chr5 38862449 N DUP 3
SRR1766470.7760159 chr5 38862255 N chr5 38862449 N DUP 5
SRR1766469.1376196 chr5 38862271 N chr5 38862465 N DUP 5
SRR1766484.1543181 chr5 38862255 N chr5 38862449 N DUP 5
SRR1766480.7569849 chr5 38862255 N chr5 38862449 N DUP 5
SRR1766458.949337 chr5 38862285 N chr5 38862384 N DEL 5
SRR1766454.10077353 chr5 38862288 N chr5 38862387 N DEL 5
SRR1766455.1203447 chr5 38862390 N chr5 38862564 N DUP 5
SRR1766442.35164889 chr5 38862393 N chr5 38862567 N DUP 5
SRR1766479.2196465 chr5 38862285 N chr5 38862432 N DEL 5
SRR1766461.9688510 chr5 38862285 N chr5 38862432 N DEL 5
SRR1766465.1349538 chr5 38862432 N chr5 38862558 N DUP 7
SRR1766466.11251498 chr5 38862432 N chr5 38862558 N DUP 7
SRR1766477.10527439 chr5 38862291 N chr5 38862487 N DEL 1
SRR1766478.9918823 chr5 38862398 N chr5 38862573 N DEL 5
SRR1766463.9324214 chr16 89417849 N chr16 89417990 N DUP 1
SRR1766477.7942558 chr16 89417886 N chr16 89417955 N DUP 5
SRR1766445.2972041 chr16 89417889 N chr16 89417958 N DUP 2
SRR1766486.8105960 chr16 89417889 N chr16 89417958 N DUP 2
SRR1766459.2548269 chr1 143218305 N chr1 143218356 N DUP 5
SRR1766449.2373281 chr1 143218125 N chr1 143218316 N DUP 5
SRR1766479.1501246 chr1 143218258 N chr1 143218407 N DUP 1
SRR1766443.5346150 chr1 143218114 N chr1 143218256 N DUP 5
SRR1766443.1076977 chr1 143218137 N chr1 143218302 N DUP 5
SRR1766481.3915051 chr1 143218138 N chr1 143218303 N DUP 5
SRR1766461.5139701 chr1 143218190 N chr1 143218410 N DUP 5
SRR1766470.10516141 chr1 143218118 N chr1 143218283 N DUP 5
SRR1766461.1718841 chr1 143218114 N chr1 143218305 N DUP 5
SRR1766469.2657001 chr1 143218205 N chr1 143218298 N DUP 7
SRR1766470.2305551 chr1 143218205 N chr1 143218298 N DUP 22
SRR1766462.2447400 chr1 143218118 N chr1 143218283 N DUP 5
SRR1766442.29016697 chr1 143218133 N chr1 143218298 N DUP 5
SRR1766461.8444079 chr1 143218196 N chr1 143218416 N DUP 5
SRR1766479.8582843 chr1 143218133 N chr1 143218298 N DUP 5
SRR1766442.19447755 chr1 143218133 N chr1 143218298 N DUP 5
SRR1766474.1707019 chr1 143218133 N chr1 143218298 N DUP 5
SRR1766476.1620330 chr1 143218166 N chr1 143218308 N DUP 5
SRR1766446.10035376 chr1 143218139 N chr1 143218304 N DUP 5
SRR1766484.834890 chr1 143218135 N chr1 143218300 N DUP 5
SRR1766477.407659 chr1 143218135 N chr1 143218300 N DUP 5
SRR1766470.2298968 chr1 143218118 N chr1 143218283 N DUP 23
SRR1766443.1166908 chr1 143218142 N chr1 143218307 N DUP 5
SRR1766466.7452790 chr1 143218190 N chr1 143218410 N DUP 4
SRR1766452.5273182 chr1 143218196 N chr1 143218416 N DUP 6
SRR1766458.1081399 chr1 143218136 N chr1 143218301 N DUP 5
SRR1766446.6167637 chr1 143218258 N chr1 143218407 N DUP 1
SRR1766484.10173210 chr1 143218114 N chr1 143218305 N DUP 5
SRR1766452.746458 chr1 143218118 N chr1 143218283 N DUP 24
SRR1766467.2479671 chr1 143218190 N chr1 143218410 N DUP 8
SRR1766476.7671085 chr1 143218132 N chr1 143218297 N DUP 8
SRR1766470.9102549 chr1 143218190 N chr1 143218410 N DUP 8
SRR1766455.1240257 chr1 143218118 N chr1 143218283 N DUP 5
SRR1766451.2149196 chr15 65864322 N chr15 65864479 N DEL 6
SRR1766470.5034301 chr15 65864366 N chr15 65864523 N DEL 6
SRR1766442.14001716 chr15 65864256 N chr15 65864590 N DUP 4
SRR1766452.212756 chr15 65864298 N chr15 65864603 N DUP 7
SRR1766449.10680438 chr15 65864298 N chr15 65864603 N DUP 7
SRR1766474.374694 chr15 65864298 N chr15 65864603 N DUP 7
SRR1766451.10065634 chr15 65864546 N chr15 65864603 N DUP 7
SRR1766478.5113766 chr15 65864546 N chr15 65864603 N DUP 7
SRR1766444.3238798 chr15 65864546 N chr15 65864603 N DUP 7
SRR1766450.8830998 chr15 65864211 N chr15 65864551 N DEL 11
SRR1766442.13788801 chr15 65864213 N chr15 65864553 N DEL 9
SRR1766455.3422400 chr15 65864214 N chr15 65864554 N DEL 8
SRR1766474.1194395 chr15 65864271 N chr15 65864578 N DEL 5
SRR1766467.1812199 chr15 65864274 N chr15 65864581 N DEL 5
SRR1766442.30350383 chr15 65864192 N chr15 65864590 N DEL 1
SRR1766451.5135594 chr15 65864193 N chr15 65864623 N DEL 11
SRR1766484.10435606 chr15 65864193 N chr15 65864623 N DEL 11
SRR1766442.13637331 chr15 65864224 N chr15 65864623 N DEL 6
SRR1766460.9135129 chr15 65864224 N chr15 65864623 N DEL 6
SRR1766442.8043184 chr15 65864224 N chr15 65864623 N DEL 6
SRR1766442.26901111 chr15 65864224 N chr15 65864623 N DEL 6
SRR1766458.2858166 chr15 65864224 N chr15 65864623 N DEL 8
SRR1766463.7034056 chr15 65864224 N chr15 65864623 N DEL 8
SRR1766484.9713825 chr6 169923983 N chr6 169924381 N DUP 16
SRR1766478.10214154 chr6 169923983 N chr6 169924381 N DUP 16
SRR1766467.9996857 chr6 169924033 N chr6 169924140 N DUP 28
SRR1766469.5036537 chr6 169923983 N chr6 169924381 N DUP 12
SRR1766463.3411238 chr6 169923983 N chr6 169924381 N DUP 11
SRR1766454.1328482 chr6 169924070 N chr6 169924194 N DEL 7
SRR1766452.1811418 chr6 169923993 N chr6 169924109 N DUP 5
SRR1766479.5250248 chr6 169923959 N chr6 169924141 N DUP 14
SRR1766473.11177425 chr6 169923954 N chr6 169924136 N DUP 10
SRR1766442.17343206 chr6 169924033 N chr6 169924254 N DUP 24
SRR1766485.449032 chr6 169924065 N chr6 169924283 N DUP 16
SRR1766455.6704533 chr6 169924033 N chr6 169924140 N DUP 18
SRR1766458.1423171 chr6 169923954 N chr6 169924136 N DUP 16
SRR1766445.2206256 chr6 169924033 N chr6 169924140 N DUP 18
SRR1766462.1454658 chr6 169923954 N chr6 169924136 N DUP 17
SRR1766456.3733458 chr6 169923954 N chr6 169924136 N DUP 17
SRR1766467.6218822 chr6 169923954 N chr6 169924136 N DUP 17
SRR1766477.7915747 chr6 169923959 N chr6 169924141 N DUP 17
SRR1766481.11745449 chr6 169923959 N chr6 169924141 N DUP 18
SRR1766468.3918415 chr6 169923954 N chr6 169924136 N DUP 20
SRR1766482.4613517 chr6 169923954 N chr6 169924136 N DUP 22
SRR1766443.7775524 chr6 169923989 N chr6 169924065 N DEL 13
SRR1766450.10520590 chr6 169923920 N chr6 169924038 N DEL 7
SRR1766461.1697056 chr6 169923980 N chr6 169924056 N DEL 10
SRR1766467.2115205 chr6 169924004 N chr6 169924105 N DUP 24
SRR1766451.4867269 chr6 169923989 N chr6 169924065 N DEL 5
SRR1766454.3008047 chr6 169923989 N chr6 169924065 N DEL 5
SRR1766467.5248265 chr6 169923991 N chr6 169924067 N DEL 3
SRR1766442.5342272 chr6 169923994 N chr6 169924070 N DEL 1
SRR1766444.5700040 chr6 169924033 N chr6 169924140 N DUP 46
SRR1766442.938096 chr6 169923967 N chr6 169924091 N DEL 10
SRR1766453.4029098 chr6 169923923 N chr6 169924092 N DEL 5
SRR1766449.7222867 chr6 169924101 N chr6 169924382 N DUP 2
SRR1766460.5590422 chr6 169924014 N chr6 169924162 N DEL 6
SRR1766454.1846509 chr6 169923990 N chr6 169924304 N DUP 5
SRR1766442.33894225 chr12 42227872 N chr12 42228095 N DUP 5
SRR1766442.37606599 chr12 42228010 N chr12 42228312 N DUP 5
SRR1766467.1702631 chr12 42228137 N chr12 42228264 N DEL 2
SRR1766459.9942971 chr12 42227995 N chr12 42228169 N DUP 5
SRR1766457.2154291 chr12 42227916 N chr12 42228189 N DEL 4
SRR1766455.10007880 chr12 42228188 N chr12 42228315 N DUP 10
SRR1766467.877846 chr12 42228069 N chr12 42228245 N DEL 2
SRR1766472.878605 chr12 42228262 N chr12 42228360 N DUP 5
SRR1766475.4098700 chr12 42228309 N chr12 42228358 N DUP 8
SRR1766471.601216 chr12 42228262 N chr12 42228360 N DUP 6
SRR1766459.7695023 chr10 2392410 N chr10 2392566 N DEL 5
SRR1766452.3386821 chr10 2392410 N chr10 2392566 N DEL 5
SRR1766476.3897371 chr10 2392410 N chr10 2392566 N DEL 5
SRR1766477.2080943 chr10 2392451 N chr10 2392570 N DEL 10
SRR1766444.5589195 chr10 2392454 N chr10 2392573 N DEL 10
SRR1766485.4708893 chr10 2392458 N chr10 2392577 N DEL 10
SRR1766479.13518341 chr10 2392458 N chr10 2392663 N DEL 8
SRR1766458.4289321 chr10 2392482 N chr10 2392730 N DEL 12
SRR1766442.37383603 chr10 2392487 N chr10 2392647 N DUP 17
SRR1766469.1566032 chr10 2392515 N chr10 2392763 N DEL 11
SRR1766458.4056319 chr10 2392488 N chr10 2392648 N DUP 12
SRR1766456.2321708 chr10 2392488 N chr10 2392605 N DUP 16
SRR1766448.229427 chr10 2392488 N chr10 2392648 N DUP 12
SRR1766474.10375373 chr10 2392620 N chr10 2392783 N DUP 28
SRR1766483.3160667 chr10 2392482 N chr10 2392730 N DEL 16
SRR1766444.656851 chr10 2392488 N chr10 2392736 N DEL 11
SRR1766485.9920992 chr10 2392600 N chr10 2392730 N DEL 15
SRR1766466.10126575 chr10 2392600 N chr10 2392730 N DEL 15
SRR1766456.2978175 chr10 2392445 N chr10 2392730 N DEL 9
SRR1766464.8410264 chr10 2392445 N chr10 2392730 N DEL 6
SRR1766442.45502902 chr10 2392486 N chr10 2392734 N DEL 5
SRR1766466.11274297 chr10 2392493 N chr10 2392741 N DEL 4
SRR1766451.3213089 chr10 2392605 N chr10 2392774 N DEL 15
SRR1766480.1168746 chr10 60240183 N chr10 60240269 N DEL 1
SRR1766482.8864026 chr10 60240183 N chr10 60240269 N DEL 4
SRR1766477.7922198 chr10 60240183 N chr10 60240269 N DEL 5
SRR1766443.193253 chr10 60240259 N chr10 60240368 N DEL 1
SRR1766479.7995816 chr10 60240259 N chr10 60240368 N DEL 5
SRR1766486.1121972 chr10 60240259 N chr10 60240368 N DEL 13
SRR1766477.8986785 chr10 60240259 N chr10 60240368 N DEL 13
SRR1766447.460340 chr10 60240162 N chr10 60240282 N DUP 31
SRR1766457.6485003 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766461.10565373 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766451.8173222 chr10 60240162 N chr10 60240282 N DUP 32
SRR1766444.5590973 chr10 60240258 N chr10 60240359 N DUP 5
SRR1766443.2558803 chr10 60240271 N chr10 60240402 N DUP 20
SRR1766451.10459403 chr10 60240271 N chr10 60240402 N DUP 13
SRR1766474.7729092 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766442.20425156 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766467.6718301 chr10 60240205 N chr10 60240303 N DEL 15
SRR1766466.3883400 chr10 60240205 N chr10 60240303 N DEL 14
SRR1766482.7427773 chr10 60240205 N chr10 60240303 N DEL 13
SRR1766483.3981936 chr10 60240174 N chr10 60240314 N DEL 4
SRR1766477.8457743 chr10 60240352 N chr10 60240433 N DEL 7
SRR1766451.8156767 chr10 60240352 N chr10 60240433 N DEL 7
SRR1766486.498212 chr10 60240352 N chr10 60240433 N DEL 7
SRR1766458.242909 chr10 60240355 N chr10 60240436 N DEL 7
SRR1766466.8624685 chr12 50378710 N chr12 50378775 N DEL 9
SRR1766449.9449617 chr12 50378716 N chr12 50378779 N DEL 6
SRR1766442.15502095 chr12 50378718 N chr12 50378781 N DEL 4
SRR1766442.812296 chr17 4933971 N chr17 4934050 N DEL 13
SRR1766452.2466527 chr17 4933973 N chr17 4934052 N DEL 18
SRR1766462.8540546 chr17 4934005 N chr17 4934085 N DEL 6
SRR1766480.3290935 chr14 34897709 N chr14 34897909 N DUP 5
SRR1766465.10238656 chrX 72179169 N chrX 72179295 N DUP 5
SRR1766461.8066145 chrX 72179282 N chrX 72179448 N DUP 3
SRR1766452.440472 chrX 72179281 N chrX 72179447 N DUP 4
SRR1766450.3422374 chrX 72179206 N chrX 72179334 N DEL 5
SRR1766472.452723 chrX 72179207 N chrX 72179374 N DUP 7
SRR1766453.2661435 chrX 72179226 N chrX 72179392 N DUP 5
SRR1766457.9295456 chrX 72179346 N chrX 72179472 N DUP 5
SRR1766471.3266159 chrX 72179346 N chrX 72179472 N DUP 5
SRR1766447.9756145 chrX 72179346 N chrX 72179472 N DUP 5
SRR1766473.11825443 chrX 72179232 N chrX 72179400 N DEL 15
SRR1766475.8277335 chr21 8464564 N chr21 8464732 N DUP 5
SRR1766454.1824241 chr21 8464345 N chr21 8464792 N DEL 8
SRR1766458.9586774 chr21 8464379 N chr21 8464624 N DEL 10
SRR1766442.13676881 chr21 8464564 N chr21 8464736 N DUP 18
SRR1766442.17271852 chr21 8464305 N chr21 8464444 N DEL 5
SRR1766460.10003694 chr21 8464327 N chr21 8464809 N DUP 5
SRR1766471.5057437 chr21 8464360 N chr21 8464663 N DEL 5
SRR1766481.3451753 chr21 8464569 N chr21 8464932 N DUP 3
SRR1766445.9717491 chr21 8464376 N chr21 8464882 N DEL 10
SRR1766455.7199638 chr21 8464297 N chr21 8464997 N DUP 5
SRR1766459.9134128 chr21 8464542 N chr21 8464712 N DEL 5
SRR1766451.7395397 chr21 8464513 N chr21 8464870 N DEL 5
SRR1766473.7180514 chr21 8464308 N chr21 8464968 N DEL 5
SRR1766442.7475928 chr21 8464340 N chr21 8464665 N DEL 5
SRR1766470.591325 chr21 8464512 N chr21 8464599 N DUP 4
SRR1766460.7110250 chr21 8464276 N chr21 8464374 N DUP 5
SRR1766483.2960922 chr21 8464389 N chr21 8464931 N DUP 9
SRR1766455.3184500 chr21 8464276 N chr21 8464996 N DUP 7
SRR1766442.24267580 chr21 8464841 N chr21 8464900 N DUP 13
SRR1766442.10665647 chr21 8464524 N chr21 8464746 N DEL 11
SRR1766473.9914864 chr21 8464346 N chr21 8464737 N DEL 9
SRR1766476.8394631 chr21 8464661 N chr21 8464931 N DUP 5
SRR1766486.4409072 chr21 8464377 N chr21 8464881 N DEL 9
SRR1766480.1786082 chr21 8464326 N chr21 8464926 N DUP 9
SRR1766484.7204063 chr21 8464341 N chr21 8464835 N DEL 9
SRR1766485.2390290 chr21 8464327 N chr21 8464803 N DEL 4
SRR1766478.685978 chr21 8464464 N chr21 8464923 N DEL 5
SRR1766442.46570216 chr21 8464378 N chr21 8464878 N DEL 7
SRR1766450.670091 chr21 8464326 N chr21 8464866 N DUP 5
SRR1766458.2189670 chr21 8464762 N chr21 8464854 N DUP 10
SRR1766461.34003 chr21 8464792 N chr21 8464898 N DUP 21
SRR1766469.8387807 chr21 8464574 N chr21 8464847 N DUP 5
SRR1766484.2942527 chr21 8464558 N chr21 8464728 N DEL 5
SRR1766472.10445186 chr21 8464276 N chr21 8464893 N DUP 3
SRR1766473.3235767 chr21 8464715 N chr21 8464897 N DUP 24
SRR1766471.2392060 chr21 8464341 N chr21 8464796 N DEL 13
SRR1766467.1222354 chr21 8464515 N chr21 8464886 N DUP 2
SRR1766449.2432414 chr21 8464354 N chr21 8464846 N DEL 9
SRR1766446.4101725 chr21 8464369 N chr21 8464869 N DEL 12
SRR1766450.4272693 chr21 8464378 N chr21 8464703 N DEL 2
SRR1766482.7714200 chr21 8464343 N chr21 8464841 N DEL 10
SRR1766444.721342 chr21 8464763 N chr21 8464907 N DUP 8
SRR1766455.9913124 chr21 8464339 N chr21 8464664 N DEL 6
SRR1766442.8810644 chr21 8464343 N chr21 8464712 N DEL 12
SRR1766442.28179648 chr21 8464343 N chr21 8464811 N DEL 9
SRR1766465.3959404 chr21 8464378 N chr21 8464882 N DEL 8
SRR1766455.6929771 chr21 8464380 N chr21 8464884 N DEL 6
SRR1766481.9529702 chr21 8464309 N chr21 8464884 N DEL 3
SRR1766456.711271 chr21 8464345 N chr21 8464599 N DEL 5
SRR1766483.4348363 chr21 8464400 N chr21 8464876 N DEL 12
SRR1766468.3617512 chr21 8464377 N chr21 8464883 N DEL 9
SRR1766443.6673159 chr21 8464587 N chr21 8464701 N DEL 5
SRR1766470.9672461 chr21 8464360 N chr21 8464878 N DEL 6
SRR1766460.8874286 chr21 8464532 N chr21 8464690 N DEL 13
SRR1766451.6536886 chr21 8464792 N chr21 8464894 N DUP 20
SRR1766448.7939414 chr21 8464341 N chr21 8464873 N DEL 7
SRR1766486.2980316 chr21 8464276 N chr21 8464712 N DUP 13
SRR1766477.9428816 chr21 8464386 N chr21 8464866 N DUP 5
SRR1766442.23940742 chr21 8464340 N chr21 8464850 N DEL 6
SRR1766467.4832535 chr21 8464789 N chr21 8464855 N DUP 10
SRR1766481.659836 chr21 8464341 N chr21 8464477 N DEL 7
SRR1766471.7694111 chr21 8464378 N chr21 8464703 N DEL 2
SRR1766479.626147 chr21 8464341 N chr21 8464668 N DEL 5
SRR1766452.21346 chr21 8464821 N chr21 8464969 N DUP 10
SRR1766442.11262696 chr21 8464309 N chr21 8464566 N DEL 14
SRR1766480.5361683 chr21 8464763 N chr21 8464907 N DUP 3
SRR1766465.5434200 chr21 8464386 N chr21 8464868 N DUP 1
SRR1766446.4705173 chr21 8464381 N chr21 8464881 N DEL 5
SRR1766453.862850 chr21 8464837 N chr21 8464896 N DUP 8
SRR1766479.4969022 chr21 8464581 N chr21 8464872 N DUP 5
SRR1766442.620304 chr21 8464833 N chr21 8464942 N DUP 21
SRR1766475.4098489 chr21 8464356 N chr21 8464685 N DEL 2
SRR1766442.15595324 chr21 8464317 N chr21 8464946 N DUP 4
SRR1766446.630456 chr21 8464377 N chr21 8464921 N DEL 5
SRR1766442.46989117 chr21 8464346 N chr21 8464429 N DEL 5
SRR1766466.5418269 chr21 8464830 N chr21 8464982 N DUP 5
SRR1766449.6438939 chr21 8464334 N chr21 8464763 N DEL 7
SRR1766464.3757429 chr21 8464532 N chr21 8464690 N DEL 13
SRR1766449.5213487 chr21 8464836 N chr21 8464905 N DUP 5
SRR1766464.1938123 chr21 8464564 N chr21 8464732 N DUP 5
SRR1766455.10015014 chr21 8464299 N chr21 8464562 N DUP 5
SRR1766465.11254159 chr21 8464351 N chr21 8464994 N DEL 5
SRR1766469.10703780 chr21 8464405 N chr21 8464903 N DEL 5
SRR1766465.1058562 chr21 8464384 N chr21 8464870 N DEL 1
SRR1766449.2873499 chr21 8464841 N chr21 8464894 N DUP 10
SRR1766479.12120908 chr21 8464386 N chr21 8464671 N DUP 14
SRR1766472.4060817 chr21 8464499 N chr21 8464763 N DUP 5
SRR1766442.1157181 chr21 8464317 N chr21 8464946 N DUP 5
SRR1766473.694178 chr21 8464386 N chr21 8464868 N DUP 1
SRR1766450.6683608 chr21 8464366 N chr21 8464604 N DEL 1
SRR1766459.1611681 chr21 8464457 N chr21 8464830 N DEL 21
SRR1766442.745341 chr21 8464330 N chr21 8464926 N DUP 2
SRR1766476.605959 chr21 8464340 N chr21 8464671 N DEL 3
SRR1766461.6805265 chr21 8464525 N chr21 8464743 N DEL 10
SRR1766447.963571 chr21 8464339 N chr21 8464891 N DEL 1
SRR1766460.2018822 chr21 8464377 N chr21 8464869 N DEL 2
SRR1766445.10115037 chr21 8464334 N chr21 8464413 N DUP 5
SRR1766481.4904471 chr21 8464584 N chr21 8464990 N DEL 4
SRR1766466.613870 chr21 8464377 N chr21 8464881 N DEL 9
SRR1766442.37524806 chr21 8464346 N chr21 8464618 N DEL 5
SRR1766473.4130301 chr21 8464524 N chr21 8464851 N DEL 1
SRR1766474.3908746 chr21 8464344 N chr21 8464830 N DEL 5
SRR1766480.3699048 chr21 8464841 N chr21 8464894 N DUP 10
SRR1766463.5777243 chr21 8464496 N chr21 8464692 N DEL 1
SRR1766467.7924805 chr21 8464405 N chr21 8464903 N DEL 5
SRR1766461.6723246 chr21 8464316 N chr21 8464581 N DEL 13
SRR1766481.12563641 chr21 8464341 N chr21 8464790 N DEL 10
SRR1766460.1772583 chr21 8464820 N chr21 8464935 N DUP 11
SRR1766482.5440054 chr21 8464330 N chr21 8464926 N DUP 2
SRR1766445.8867467 chr21 8464560 N chr21 8464642 N DUP 5
SRR1766442.33858989 chr21 8464542 N chr21 8464712 N DEL 2
SRR1766446.6490081 chr21 8464792 N chr21 8464900 N DUP 25
SRR1766446.2261520 chr21 8464576 N chr21 8464881 N DUP 1
SRR1766485.5818323 chr21 8464742 N chr21 8465013 N DUP 10
SRR1766463.8530599 chr21 8464399 N chr21 8464527 N DEL 2
SRR1766444.1655131 chr21 8464385 N chr21 8464919 N DUP 10
SRR1766458.5269397 chr21 8464277 N chr21 8464695 N DUP 1
SRR1766478.11848773 chr21 8464395 N chr21 8464841 N DEL 10
SRR1766482.3258177 chr21 8464603 N chr21 8464890 N DEL 5
SRR1766453.7794336 chr21 8464794 N chr21 8464902 N DUP 34
SRR1766475.8472962 chr21 8464340 N chr21 8464882 N DEL 2
SRR1766461.8239120 chr21 8464399 N chr21 8464780 N DEL 14
SRR1766459.2654123 chr21 8464450 N chr21 8464998 N DEL 9
SRR1766452.9773891 chr21 8464324 N chr21 8464882 N DEL 5
SRR1766484.5282827 chr10 120793074 N chr10 120793440 N DEL 5
SRR1766453.2495297 chr3 9822857 N chr3 9822924 N DEL 7
SRR1766457.6639652 chr21 34670028 N chr21 34670329 N DEL 11
SRR1766455.4043273 chr21 34670048 N chr21 34670169 N DEL 5
SRR1766451.6958305 chr21 34670050 N chr21 34670171 N DEL 5
SRR1766474.9565566 chr21 34670048 N chr21 34670169 N DEL 8
SRR1766447.6241773 chr21 34670048 N chr21 34670169 N DEL 5
SRR1766467.1224372 chr21 34670028 N chr21 34670327 N DUP 4
SRR1766442.4241701 chr21 34670067 N chr21 34670338 N DEL 6
SRR1766466.5498767 chr6 16616704 N chr6 16616761 N DEL 11
SRR1766464.5343103 chr12 59486432 N chr12 59486505 N DUP 7
SRR1766485.365663 chr12 59486432 N chr12 59486505 N DUP 7
SRR1766454.6793110 chr12 5929418 N chr12 5929493 N DEL 5
SRR1766455.408025 chr12 5929430 N chr12 5929653 N DEL 5
SRR1766477.4271506 chr12 5929427 N chr12 5929650 N DEL 5
SRR1766451.6226572 chr12 5929464 N chr12 5929613 N DEL 1
SRR1766460.9137463 chr12 5929427 N chr12 5929650 N DEL 5
SRR1766442.14279952 chr12 5929310 N chr12 5929453 N DUP 10
SRR1766442.11314633 chr12 5929310 N chr12 5929453 N DUP 10
SRR1766459.10593179 chr12 5929310 N chr12 5929453 N DUP 11
SRR1766453.1126053 chr12 5929481 N chr12 5929704 N DEL 4
SRR1766442.40349687 chr12 5929481 N chr12 5929704 N DEL 2
SRR1766472.8895753 chr12 5929310 N chr12 5929453 N DUP 15
SRR1766452.3700988 chr12 5929310 N chr12 5929453 N DUP 15
SRR1766473.529077 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766465.6848241 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766481.4209435 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766474.9457543 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766485.11783333 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766443.1801683 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766469.1366437 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766448.8597871 chr12 5929427 N chr12 5929650 N DEL 5
SRR1766481.7697176 chr12 5929419 N chr12 5929492 N DUP 5
SRR1766458.7161007 chr12 5929487 N chr12 5929782 N DUP 10
SRR1766454.7436758 chr12 5929419 N chr12 5929492 N DUP 5
SRR1766442.6809372 chr12 5929419 N chr12 5929492 N DUP 5
SRR1766477.2409670 chr12 5929419 N chr12 5929492 N DUP 5
SRR1766464.5984668 chr12 5929501 N chr12 5929650 N DEL 10
SRR1766447.8588736 chr12 5929419 N chr12 5929492 N DUP 6
SRR1766443.286116 chr12 5929566 N chr12 5929641 N DEL 5
SRR1766443.2697334 chr12 5929403 N chr12 5929550 N DUP 10
SRR1766464.1168502 chr12 5929599 N chr12 5929746 N DUP 10
SRR1766485.6063647 chr12 5929599 N chr12 5929746 N DUP 10
SRR1766476.2299154 chr12 5929380 N chr12 5929599 N DEL 5
SRR1766477.11129207 chr12 5929380 N chr12 5929599 N DEL 5
SRR1766442.10393556 chr12 5929310 N chr12 5929675 N DUP 4
SRR1766478.2533654 chr12 5929310 N chr12 5929675 N DUP 5
SRR1766483.11302872 chr12 5929386 N chr12 5929605 N DEL 5
SRR1766442.23668787 chr12 5929395 N chr12 5929614 N DEL 5
SRR1766465.696922 chr12 5929413 N chr12 5929782 N DUP 18
SRR1766442.36054067 chr12 5929630 N chr12 5929703 N DUP 5
SRR1766469.6104689 chr12 5929402 N chr12 5929621 N DEL 5
SRR1766466.2117814 chr12 5929337 N chr12 5929630 N DEL 5
SRR1766442.42200809 chr12 5929413 N chr12 5929782 N DUP 15
SRR1766465.3969839 chr12 5929413 N chr12 5929782 N DUP 15
SRR1766467.692760 chr12 5929492 N chr12 5929641 N DEL 5
SRR1766484.9151315 chr12 5929635 N chr12 5929782 N DUP 10
SRR1766448.6711066 chr12 5929413 N chr12 5929782 N DUP 15
SRR1766469.9006952 chr12 5929310 N chr12 5929675 N DUP 5
SRR1766460.2502789 chr12 5929310 N chr12 5929675 N DUP 5
SRR1766445.4204844 chr12 5929492 N chr12 5929641 N DEL 5
SRR1766456.3939774 chr12 5929413 N chr12 5929782 N DUP 10
SRR1766463.5892525 chr12 5929418 N chr12 5929713 N DUP 5
SRR1766448.8184556 chr12 5929492 N chr12 5929641 N DEL 5
SRR1766470.250806 chr12 5929492 N chr12 5929641 N DEL 5
SRR1766474.9591594 chr12 5929492 N chr12 5929641 N DEL 5
SRR1766443.1801683 chr12 5929429 N chr12 5929652 N DEL 10
SRR1766482.6561632 chr12 5929337 N chr12 5929630 N DEL 5
SRR1766445.8424435 chr12 5929492 N chr12 5929641 N DEL 5
SRR1766476.6140423 chr12 5929630 N chr12 5929703 N DUP 10
SRR1766466.621726 chr12 5929487 N chr12 5929782 N DUP 15
SRR1766477.10533136 chr12 5929310 N chr12 5929383 N DUP 15
SRR1766482.2985557 chr12 5929506 N chr12 5929655 N DEL 5
SRR1766446.1555345 chr12 5929418 N chr12 5929713 N DUP 5
SRR1766449.1295593 chr12 5929348 N chr12 5929641 N DEL 10
SRR1766466.10933280 chr12 5929492 N chr12 5929641 N DEL 5
SRR1766469.6428948 chr12 5929498 N chr12 5929647 N DEL 5
SRR1766464.694524 chr12 5929427 N chr12 5929650 N DEL 5
SRR1766442.36126599 chr12 5929481 N chr12 5929704 N DEL 10
SRR1766456.2078241 chr12 5929501 N chr12 5929650 N DEL 10
SRR1766469.2484114 chr12 5929481 N chr12 5929704 N DEL 6
SRR1766448.10418503 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766470.10141030 chr12 5929413 N chr12 5929782 N DUP 15
SRR1766481.11343330 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766442.46155632 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766482.10295176 chr12 5929413 N chr12 5929782 N DUP 10
SRR1766442.29850140 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766478.1657900 chr12 5929413 N chr12 5929782 N DUP 9
SRR1766482.11883983 chr12 5929317 N chr12 5929703 N DUP 1
SRR1766473.4342316 chr12 5929413 N chr12 5929782 N DUP 12
SRR1766454.2961043 chr12 5929413 N chr12 5929782 N DUP 12
SRR1766451.6561987 chr11 71098183 N chr11 71098435 N DUP 2
SRR1766443.94490 chr10 132980543 N chr10 132980609 N DEL 9
SRR1766471.7033430 chr10 132980594 N chr10 132980836 N DEL 1
SRR1766459.9979723 chr10 132980583 N chr10 132980781 N DEL 1
SRR1766442.31065082 chr10 132980618 N chr10 132980772 N DEL 10
SRR1766454.2308710 chr10 132980531 N chr10 132980847 N DUP 5
SRR1766463.9952196 chr10 132980618 N chr10 132980825 N DUP 5
SRR1766461.7176706 chr10 132980758 N chr10 132980836 N DEL 10
SRR1766481.4141272 chr10 132980702 N chr10 132980909 N DUP 10
SRR1766442.47100771 chr10 132980715 N chr10 132980779 N DUP 5
SRR1766473.10628996 chr10 132980780 N chr10 132980954 N DUP 10
SRR1766460.9222259 chr10 132980592 N chr10 132980876 N DUP 10
SRR1766459.4747082 chr10 132980780 N chr10 132980954 N DUP 5
SRR1766485.9369820 chr10 132980622 N chr10 132980927 N DUP 4
SRR1766443.4889964 chr10 132980602 N chr10 132980940 N DUP 5
SRR1766460.7856237 chr10 132980591 N chr10 132980962 N DUP 5
SRR1766464.610714 chr10 132980639 N chr10 132980870 N DEL 10
SRR1766455.5502769 chr10 132980928 N chr10 132980993 N DUP 4
SRR1766479.10310734 chr10 132980692 N chr10 132980890 N DEL 17
SRR1766447.10545792 chr10 132980648 N chr10 132980955 N DEL 10
SRR1766483.8506841 chr10 132980919 N chr10 132981018 N DEL 6
SRR1766473.3961923 chr10 132980919 N chr10 132981018 N DEL 5
SRR1766468.3414348 chr10 132980919 N chr10 132981018 N DEL 5
SRR1766465.3087414 chrX 107204842 N chrX 107205043 N DEL 2
SRR1766458.5361336 chrX 107204842 N chrX 107205043 N DEL 3
SRR1766473.4107834 chrX 107204842 N chrX 107205043 N DEL 12
SRR1766483.2792806 chrX 107204842 N chrX 107205043 N DEL 13
SRR1766486.3641391 chrX 107204870 N chrX 107205043 N DEL 21
SRR1766468.1757784 chrX 107204870 N chrX 107205043 N DEL 24
SRR1766462.2979910 chrX 107204870 N chrX 107205043 N DEL 26
SRR1766478.3051211 chrX 107204827 N chrX 107204882 N DUP 26
SRR1766442.9865723 chrX 107204827 N chrX 107204882 N DUP 26
SRR1766443.4347326 chrX 107204827 N chrX 107205110 N DUP 33
SRR1766454.3763868 chrX 107204827 N chrX 107205110 N DUP 30
SRR1766471.9933313 chrX 107204827 N chrX 107205110 N DUP 31
SRR1766486.1230929 chrX 107204847 N chrX 107204902 N DUP 26
SRR1766463.2942810 chrX 107204827 N chrX 107204882 N DUP 26
SRR1766466.9635048 chrX 107204870 N chrX 107204967 N DEL 13
SRR1766471.7817743 chrX 107204870 N chrX 107204967 N DEL 13
SRR1766473.3981399 chrX 107204922 N chrX 107205043 N DEL 20
SRR1766462.9059923 chrX 107204827 N chrX 107204882 N DUP 19
SRR1766484.7167012 chrX 107204827 N chrX 107204882 N DUP 19
SRR1766478.11061727 chrX 107204922 N chrX 107205043 N DEL 15
SRR1766480.8300932 chrX 107204922 N chrX 107205043 N DEL 14
SRR1766470.4514772 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766457.6266848 chrX 107204827 N chrX 107205110 N DUP 34
SRR1766464.7782581 chrX 107204898 N chrX 107205019 N DEL 13
SRR1766457.7288802 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766466.4236866 chrX 107204898 N chrX 107205043 N DEL 27
SRR1766485.724969 chrX 107204898 N chrX 107205043 N DEL 27
SRR1766486.3641391 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766453.6069706 chrX 107204827 N chrX 107204906 N DUP 15
SRR1766465.2348161 chrX 107204898 N chrX 107205043 N DEL 26
SRR1766447.6559092 chrX 107204898 N chrX 107205043 N DEL 26
SRR1766475.5690233 chrX 107204827 N chrX 107204906 N DUP 19
SRR1766467.9269252 chrX 107204922 N chrX 107205043 N DEL 21
SRR1766459.5660222 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766465.2885075 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766477.6988972 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766462.11206093 chrX 107204922 N chrX 107205043 N DEL 13
SRR1766468.4946384 chrX 107204842 N chrX 107205043 N DEL 13
SRR1766447.6559092 chrX 107204846 N chrX 107205047 N DEL 11
SRR1766462.11206093 chrX 107204853 N chrX 107205054 N DEL 4
SRR1766477.11794956 chrX 107204866 N chrX 107205071 N DEL 9
SRR1766443.10307533 chrX 54607144 N chrX 54607209 N DEL 3
SRR1766453.1693973 chrX 54607144 N chrX 54607209 N DEL 7
SRR1766463.5104021 chrX 54607144 N chrX 54607209 N DEL 7
SRR1766470.5027380 chr19 40377188 N chr19 40377495 N DEL 6
SRR1766460.4998436 chr19 40377071 N chr19 40377273 N DUP 5
SRR1766454.4028571 chr19 40377443 N chr19 40377511 N DUP 30
SRR1766476.4176311 chr21 8244412 N chr21 8244478 N DUP 4
SRR1766466.1923431 chr21 8244409 N chr21 8244479 N DUP 1
SRR1766472.5999522 chr3 887332 N chr3 887388 N DEL 10
SRR1766476.8866578 chr3 887332 N chr3 887388 N DEL 10
SRR1766483.2546936 chr3 887342 N chr3 887402 N DEL 1
SRR1766473.7521504 chr14 105327922 N chr14 105328111 N DEL 5
SRR1766481.11573596 chr15 32417583 N chr15 32417635 N DUP 5
SRR1766470.2461658 chr16 88831839 N chr16 88832042 N DEL 5
SRR1766455.7284046 chr1 34102722 N chr1 34102780 N DEL 5
SRR1766448.8725288 chr1 34102722 N chr1 34102818 N DEL 5
SRR1766447.11066493 chr1 34102722 N chr1 34102818 N DEL 5
SRR1766453.7127672 chr1 34102722 N chr1 34102818 N DEL 19
SRR1766477.4047385 chr1 34102728 N chr1 34102784 N DUP 15
SRR1766481.12021832 chr1 34102728 N chr1 34102784 N DUP 19
SRR1766484.5433352 chr1 34102766 N chr1 34102824 N DEL 34
SRR1766453.3143994 chr1 34102766 N chr1 34102824 N DEL 30
SRR1766443.8046965 chr1 34102766 N chr1 34102824 N DEL 28
SRR1766443.1788655 chr1 34102722 N chr1 34102818 N DEL 18
SRR1766457.6683676 chr1 34102722 N chr1 34102818 N DEL 17
SRR1766475.5642958 chr1 34102722 N chr1 34102818 N DEL 20
SRR1766464.5833726 chr1 34102722 N chr1 34102818 N DEL 17
SRR1766452.4723694 chr1 34102766 N chr1 34102824 N DEL 25
SRR1766478.3716221 chr1 34102766 N chr1 34102824 N DEL 25
SRR1766465.4371388 chr1 34102722 N chr1 34102818 N DEL 5
SRR1766481.5713646 chr1 34102766 N chr1 34102824 N DEL 21
SRR1766486.2116935 chr1 34102724 N chr1 34102820 N DEL 5
SRR1766475.2411998 chr1 34102712 N chr1 34102827 N DEL 12
SRR1766459.3958705 chr1 34102721 N chr1 34102836 N DEL 3
SRR1766459.10498539 chr1 34102714 N chr1 34102829 N DEL 10
SRR1766478.5525424 chr1 34102714 N chr1 34102829 N DEL 10
SRR1766467.2872865 chr1 118225744 N chr1 118225860 N DEL 1
SRR1766458.7095308 chr8 28463387 N chr8 28463520 N DEL 10
SRR1766456.2343785 chr8 28463307 N chr8 28463460 N DEL 5
SRR1766468.1945978 chr8 28463492 N chr8 28463549 N DEL 1
SRR1766473.1646758 chr16 77713959 N chr16 77714021 N DEL 5
SRR1766473.1646758 chr16 77713966 N chr16 77714026 N DUP 5
SRR1766447.2056282 chr16 77713960 N chr16 77714020 N DUP 5
SRR1766485.1236663 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766461.7417626 chr16 77713978 N chr16 77714221 N DUP 14
SRR1766452.4185721 chr16 77713974 N chr16 77714217 N DUP 7
SRR1766471.5530269 chr16 77713978 N chr16 77714221 N DUP 11
SRR1766447.6561819 chr16 77713974 N chr16 77714034 N DUP 1
SRR1766468.1127984 chr16 77713974 N chr16 77714217 N DUP 10
SRR1766470.4539864 chr16 77714034 N chr16 77714279 N DEL 10
SRR1766479.7692193 chr16 77713960 N chr16 77714264 N DUP 8
SRR1766475.4264379 chr16 77713916 N chr16 77713991 N DEL 2
SRR1766456.5828534 chr16 77713960 N chr16 77714020 N DUP 5
SRR1766482.4415151 chr16 77713960 N chr16 77714020 N DUP 5
SRR1766483.11854027 chr16 77714071 N chr16 77714375 N DUP 5
SRR1766442.6683352 chr16 77713988 N chr16 77714048 N DUP 2
SRR1766464.3285261 chr16 77713960 N chr16 77714081 N DUP 4
SRR1766479.1270044 chr16 77714071 N chr16 77714375 N DUP 5
SRR1766477.8245138 chr16 77713960 N chr16 77714081 N DUP 5
SRR1766442.14867442 chr16 77713960 N chr16 77714081 N DUP 5
SRR1766444.115041 chr16 77713960 N chr16 77714081 N DUP 5
SRR1766452.6609368 chr16 77714009 N chr16 77714071 N DEL 5
SRR1766472.3059684 chr16 77714009 N chr16 77714071 N DEL 5
SRR1766458.4030495 chr16 77713960 N chr16 77714081 N DUP 5
SRR1766445.4851760 chr16 77713888 N chr16 77713963 N DEL 2
SRR1766475.1924080 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766471.7393756 chr16 77713945 N chr16 77714249 N DUP 14
SRR1766479.12483281 chr16 77713974 N chr16 77714217 N DUP 5
SRR1766466.3808934 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766477.461687 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766470.2704532 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766448.5973104 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766442.26447917 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766459.5599482 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766447.3685595 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766484.5039321 chr16 77713885 N chr16 77714143 N DEL 5
SRR1766459.5389597 chr16 77713887 N chr16 77714145 N DEL 5
SRR1766451.2528521 chr16 77714038 N chr16 77714222 N DEL 7
SRR1766462.3000269 chr16 77714038 N chr16 77714222 N DEL 8
SRR1766448.7793587 chr16 77713977 N chr16 77714222 N DEL 4
SRR1766477.10337537 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766448.3695286 chr16 77714034 N chr16 77714218 N DEL 5
SRR1766464.8336984 chr16 77713974 N chr16 77714278 N DUP 5
SRR1766477.461687 chr16 77714157 N chr16 77714217 N DUP 5
SRR1766477.9694789 chr16 77714218 N chr16 77714339 N DUP 5
SRR1766449.3850380 chr16 77714034 N chr16 77714218 N DEL 5
SRR1766467.587397 chr16 77714157 N chr16 77714217 N DUP 5
SRR1766470.4669954 chr16 77714034 N chr16 77714218 N DEL 5
SRR1766471.3247598 chr16 77714034 N chr16 77714218 N DEL 5
SRR1766479.4585769 chr16 77714034 N chr16 77714218 N DEL 5
SRR1766449.5567257 chr16 77714157 N chr16 77714217 N DUP 5
SRR1766477.11329342 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766457.4679150 chr16 77714038 N chr16 77714222 N DEL 9
SRR1766445.8151642 chr16 77714034 N chr16 77714218 N DEL 5
SRR1766458.7741035 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766446.7094752 chr16 77713978 N chr16 77714221 N DUP 15
SRR1766471.3247598 chr16 77713974 N chr16 77714278 N DUP 5
SRR1766449.9990780 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766485.2350102 chr16 77714062 N chr16 77714246 N DEL 10
SRR1766442.8319229 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766442.8142213 chr16 77714038 N chr16 77714222 N DEL 10
SRR1766465.3766743 chr16 77713977 N chr16 77714222 N DEL 10
SRR1766476.4967565 chr16 77713845 N chr16 77714225 N DEL 10
SRR1766451.3253584 chr16 77713960 N chr16 77714264 N DUP 5
SRR1766453.8368872 chr16 77714228 N chr16 77714587 N DUP 5
SRR1766479.12483281 chr16 77714034 N chr16 77714279 N DEL 9
SRR1766480.602535 chr16 77714279 N chr16 77714339 N DUP 5
SRR1766457.8639579 chr16 77714034 N chr16 77714279 N DEL 7
SRR1766442.20225464 chr16 77714034 N chr16 77714279 N DEL 6
SRR1766458.5014427 chr16 77714071 N chr16 77714253 N DUP 1
SRR1766469.10886800 chr16 77714071 N chr16 77714253 N DUP 1
SRR1766447.6917605 chr16 77714071 N chr16 77714253 N DUP 2
SRR1766453.10968362 chr16 77714071 N chr16 77714253 N DUP 4
SRR1766442.4623241 chr16 77713974 N chr16 77714217 N DUP 4
SRR1766469.362655 chr16 77714071 N chr16 77714253 N DUP 5
SRR1766442.34248598 chr16 77713978 N chr16 77714221 N DUP 9
SRR1766449.3850380 chr16 77714071 N chr16 77714253 N DUP 5
SRR1766449.9995154 chr16 77714034 N chr16 77714279 N DEL 5
SRR1766468.3943243 chr16 77713978 N chr16 77714221 N DUP 10
SRR1766472.11653910 chr16 77714100 N chr16 77714221 N DUP 10
SRR1766455.1866751 chr16 77713974 N chr16 77714217 N DUP 5
SRR1766461.7417626 chr16 77713960 N chr16 77714264 N DUP 5
SRR1766449.1647445 chr16 77714034 N chr16 77714279 N DEL 5
SRR1766482.4415151 chr16 77714275 N chr16 77714457 N DUP 5
SRR1766485.10259289 chr16 77713960 N chr16 77714264 N DUP 5
SRR1766450.8966939 chr16 77714034 N chr16 77714279 N DEL 5
SRR1766464.3547367 chr16 77714034 N chr16 77714279 N DEL 5
SRR1766470.928911 chr16 77713974 N chr16 77714217 N DUP 5
SRR1766449.2884125 chr16 77714034 N chr16 77714279 N DEL 5
SRR1766442.22500358 chr16 77713978 N chr16 77714221 N DUP 10
SRR1766473.5310134 chr16 77713978 N chr16 77714221 N DUP 10
SRR1766443.1932068 chr16 77713960 N chr16 77714264 N DUP 5
SRR1766463.7277456 chr16 77713960 N chr16 77714264 N DUP 5
SRR1766451.2448077 chr16 77713960 N chr16 77714264 N DUP 5
SRR1766442.8319229 chr16 77713960 N chr16 77714264 N DUP 5
SRR1766464.9869033 chr16 77713978 N chr16 77714221 N DUP 11
SRR1766476.1684303 chr16 77714034 N chr16 77714279 N DEL 5
SRR1766467.8685699 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766446.9313097 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766464.9869033 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766452.2336657 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766453.7909117 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766474.6044085 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766453.7217103 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766442.14867442 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766476.8151780 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766480.1609384 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766450.554946 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766467.10385950 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766486.469049 chr16 77714218 N chr16 77714339 N DUP 10
SRR1766480.59524 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766484.4081816 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766482.4856079 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766474.4073984 chr16 77714143 N chr16 77714264 N DUP 5
SRR1766467.293977 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766448.1705051 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766461.8854497 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766480.7444091 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766467.9079179 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766480.1609384 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766467.4919345 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766442.27455245 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766482.5868814 chr16 77714020 N chr16 77714143 N DEL 5
SRR1766477.8245138 chr16 77714133 N chr16 77714378 N DEL 5
SRR1766473.11219750 chr16 77714133 N chr16 77714378 N DEL 5
SRR1766442.43139 chr16 77714133 N chr16 77714378 N DEL 5
SRR1766442.15390481 chr16 77714133 N chr16 77714378 N DEL 5
SRR1766443.1932068 chr16 77714133 N chr16 77714378 N DEL 5
SRR1766454.596053 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766458.7946766 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766477.2710984 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766479.11971227 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766470.2976153 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766475.10402152 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766472.4292333 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766464.3285261 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766454.10932212 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766479.7692193 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766465.1623954 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766461.5411160 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766462.3000269 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766445.7680878 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766461.1614457 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766463.7277456 chr16 77714011 N chr16 77714378 N DEL 5
SRR1766455.6059336 chr16 77713881 N chr16 77714383 N DEL 5
SRR1766462.10955584 chr7 108585315 N chr7 108585388 N DUP 2
SRR1766472.11431254 chr7 108585315 N chr7 108585388 N DUP 2
SRR1766465.333060 chr22 48584648 N chr22 48585059 N DEL 1
SRR1766480.6266090 chr22 48584654 N chr22 48585050 N DEL 4
SRR1766455.7563926 chr22 48584486 N chr22 48584686 N DUP 6
SRR1766467.4542356 chr22 48584634 N chr22 48584771 N DUP 1
SRR1766482.4874365 chr22 48584504 N chr22 48584673 N DEL 9
SRR1766452.974154 chr22 48584689 N chr22 48584812 N DUP 5
SRR1766477.5691124 chr22 48584658 N chr22 48584744 N DEL 5
SRR1766453.10861472 chr19 50377009 N chr19 50377083 N DUP 3
SRR1766476.9806305 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766447.7674177 chr16 46401604 N chr16 46401925 N DUP 6
SRR1766478.5936796 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766477.5248982 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766478.9651247 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766463.8502224 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766454.5040531 chr16 46401600 N chr16 46401746 N DUP 5
SRR1766447.1417977 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766483.10549275 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766462.1753586 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766442.19645423 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766484.5739339 chr16 46401590 N chr16 46401713 N DUP 3
SRR1766483.12512599 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766448.481280 chr16 46401603 N chr16 46401921 N DUP 4
SRR1766476.3684383 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766459.713195 chr16 46401598 N chr16 46401893 N DUP 4
SRR1766461.7961472 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766457.182032 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766472.594471 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766486.751975 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766465.8651395 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766475.5327683 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766463.7023723 chr16 46401619 N chr16 46401742 N DUP 5
SRR1766470.9621184 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766476.5660747 chr16 46401622 N chr16 46401790 N DUP 8
SRR1766442.24138561 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766475.9701027 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766466.373593 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766442.32715017 chr16 46401623 N chr16 46401746 N DUP 1
SRR1766446.9490615 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766466.241010 chr16 46401708 N chr16 46401804 N DUP 5
SRR1766486.9465990 chr16 46401643 N chr16 46401814 N DUP 2
SRR1766479.2731281 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766483.2953988 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766451.3840824 chr16 46401754 N chr16 46401879 N DEL 5
SRR1766454.1227289 chr1 205830853 N chr1 205830918 N DEL 3
SRR1766484.11919070 chr9 24100001 N chr9 24100138 N DEL 5
SRR1766484.6934444 chr9 24100027 N chr9 24100088 N DUP 10
SRR1766459.141951 chr9 24100087 N chr9 24100163 N DEL 15
SRR1766482.10868281 chr9 24100087 N chr9 24100163 N DEL 9
SRR1766469.6932174 chr3 22379370 N chr3 22379649 N DEL 9
SRR1766465.5448123 chr3 22379368 N chr3 22379427 N DUP 5
SRR1766468.2231961 chr3 22379396 N chr3 22379459 N DUP 5
SRR1766466.6479193 chr3 22379366 N chr3 22379481 N DUP 5
SRR1766464.7146132 chr3 22379398 N chr3 22379489 N DUP 10
SRR1766457.1895463 chr3 22379397 N chr3 22379472 N DUP 12
SRR1766484.633396 chr3 22379429 N chr3 22379674 N DUP 7
SRR1766443.4299081 chr5 1272674 N chr5 1272743 N DEL 2
SRR1766474.7432449 chr5 1272674 N chr5 1273690 N DEL 3
SRR1766460.4027190 chr5 1272722 N chr5 1273234 N DEL 10
SRR1766451.4601320 chr5 1272674 N chr5 1273690 N DEL 5
SRR1766465.11290015 chr5 1272674 N chr5 1273690 N DEL 5
SRR1766486.9056919 chr5 1272674 N chr5 1273724 N DEL 25
SRR1766464.9101210 chr5 1272674 N chr5 1273724 N DEL 33
SRR1766448.9611073 chr5 1272688 N chr5 1272901 N DEL 14
SRR1766476.8657152 chr5 1272674 N chr5 1273724 N DEL 28
SRR1766482.8219950 chr5 1272688 N chr5 1273270 N DEL 14
SRR1766452.1353494 chr5 1272828 N chr5 1273883 N DEL 10
SRR1766455.188779 chr5 1273738 N chr5 1273850 N DUP 14
SRR1766462.10635448 chr5 1272759 N chr5 1273117 N DUP 10
SRR1766482.3332762 chr5 1272761 N chr5 1273673 N DUP 13
SRR1766451.10431201 chr5 1272898 N chr5 1273234 N DEL 4
SRR1766476.4105952 chr5 1272854 N chr5 1273258 N DUP 5
SRR1766482.7756251 chr5 1272974 N chr5 1273238 N DEL 5
SRR1766451.6609716 chr5 1272974 N chr5 1273238 N DEL 5
SRR1766464.6504791 chr5 1272833 N chr5 1272976 N DEL 1
SRR1766446.3537281 chr5 1272990 N chr5 1273218 N DEL 3
SRR1766476.3700204 chr5 1272770 N chr5 1273246 N DUP 5
SRR1766476.4105952 chr5 1272762 N chr5 1273120 N DUP 6
SRR1766464.866160 chr5 1273146 N chr5 1273258 N DUP 2
SRR1766464.10805325 chr5 1272702 N chr5 1273171 N DEL 1
SRR1766482.11112772 chr5 1272921 N chr5 1273217 N DUP 12
SRR1766469.6686642 chr5 1272915 N chr5 1273095 N DUP 12
SRR1766456.4037959 chr5 1272758 N chr5 1273157 N DUP 5
SRR1766443.4299081 chr5 1272984 N chr5 1273135 N DEL 7
SRR1766486.3429159 chr5 1272722 N chr5 1272829 N DEL 2
SRR1766467.10309732 chr5 1272878 N chr5 1273979 N DEL 5
SRR1766453.976552 chr5 1272878 N chr5 1273979 N DEL 5
SRR1766471.11449076 chr5 1272678 N chr5 1272957 N DUP 1
SRR1766482.11883006 chr5 1272880 N chr5 1273940 N DEL 10
SRR1766456.6498723 chr5 1272808 N chr5 1273650 N DEL 7
SRR1766454.4863295 chr5 1272688 N chr5 1272899 N DUP 5
SRR1766483.4279854 chr5 1272723 N chr5 1272970 N DUP 5
SRR1766474.5045022 chr5 1272950 N chr5 1273940 N DEL 12
SRR1766446.5732889 chr5 1272926 N chr5 1273106 N DUP 8
SRR1766454.8034845 chr5 1272688 N chr5 1273039 N DUP 5
SRR1766463.3371660 chr5 1272744 N chr5 1272957 N DEL 5
SRR1766461.10313243 chr5 1272833 N chr5 1273010 N DEL 4
SRR1766459.9700305 chr5 1273137 N chr5 1273285 N DUP 8
SRR1766467.4058410 chr5 1272802 N chr5 1273526 N DEL 9
SRR1766451.4002328 chr5 1272646 N chr5 1272824 N DUP 18
SRR1766474.6306011 chr5 1272828 N chr5 1273738 N DEL 20
SRR1766486.5221576 chr5 1272792 N chr5 1273738 N DEL 9
SRR1766478.6070231 chr5 1272828 N chr5 1273738 N DEL 11
SRR1766463.10454938 chr5 1272857 N chr5 1273699 N DEL 5
SRR1766462.1593480 chr5 1272950 N chr5 1273940 N DEL 33
SRR1766453.8101317 chr5 1272844 N chr5 1273940 N DEL 29
SRR1766460.8119854 chr5 1272950 N chr5 1273940 N DEL 36
SRR1766459.4436321 chr5 1272844 N chr5 1273940 N DEL 29
SRR1766483.2079340 chr5 1272950 N chr5 1273940 N DEL 36
SRR1766472.437435 chr5 1272950 N chr5 1273940 N DEL 36
SRR1766461.10590260 chr5 1272950 N chr5 1273940 N DEL 35
SRR1766452.1640759 chr5 1272844 N chr5 1273940 N DEL 24
SRR1766476.9508035 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766480.5186410 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766442.12661975 chr5 1272817 N chr5 1273951 N DEL 27
SRR1766442.43499975 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766468.5427890 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766480.8591848 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766460.8119854 chr5 1272772 N chr5 1273940 N DEL 27
SRR1766449.7348751 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766481.1203964 chr5 1272808 N chr5 1273940 N DEL 20
SRR1766448.8659739 chr5 1272705 N chr5 1273941 N DEL 14
SRR1766462.11127400 chr5 1272709 N chr5 1273945 N DEL 10
SRR1766450.6397588 chr5 1272707 N chr5 1273943 N DEL 12
SRR1766452.1028794 chr5 1272706 N chr5 1273942 N DEL 13
SRR1766460.7266798 chr5 1272712 N chr5 1273948 N DEL 7
SRR1766468.653379 chr5 1272716 N chr5 1273952 N DEL 3
SRR1766442.12861091 chr7 1295473 N chr7 1295557 N DUP 12
SRR1766442.19980291 chr7 1295515 N chr7 1295601 N DUP 8
SRR1766480.6512380 chr7 1295517 N chr7 1295603 N DUP 13
SRR1766460.10594615 chr7 1295478 N chr7 1295564 N DEL 2
SRR1766474.6466550 chr7 1295491 N chr7 1295575 N DEL 5
SRR1766485.4631770 chr7 1295512 N chr7 1295592 N DEL 22
SRR1766451.1278231 chr7 1295428 N chr7 1295702 N DEL 14
SRR1766442.2573565 chr7 1295448 N chr7 1295722 N DEL 5
SRR1766478.11455743 chr7 1295443 N chr7 1295717 N DEL 10
SRR1766486.7928276 chr7 1295451 N chr7 1295725 N DEL 3
SRR1766474.6047719 chr15 72396428 N chr15 72396585 N DEL 1
SRR1766442.41742928 chr15 72396594 N chr15 72396709 N DUP 2
SRR1766452.6331120 chr7 45813283 N chr7 45813382 N DEL 10
SRR1766444.91059 chr7 45813324 N chr7 45813505 N DEL 18
SRR1766482.488163 chr7 45813249 N chr7 45813444 N DUP 11
SRR1766462.1769388 chr7 45813276 N chr7 45813586 N DUP 1
SRR1766470.6002787 chr7 45813488 N chr7 45813602 N DUP 6
SRR1766453.8521863 chr19 57138063 N chr19 57138228 N DEL 6
SRR1766449.4570193 chr19 57137989 N chr19 57138060 N DUP 8
SRR1766469.10089654 chr19 57137989 N chr19 57138068 N DUP 5
SRR1766442.15979870 chr19 57138034 N chr19 57138141 N DUP 2
SRR1766445.3513444 chr19 57138016 N chr19 57138178 N DUP 14
SRR1766465.6743129 chr19 57138060 N chr19 57138116 N DUP 13
SRR1766475.7586315 chr19 57137986 N chr19 57138146 N DUP 12
SRR1766469.5791321 chr19 57137992 N chr19 57138139 N DUP 5
SRR1766469.10762129 chr19 57138052 N chr19 57138155 N DUP 10
SRR1766474.60635 chr19 57138024 N chr19 57138099 N DUP 13
SRR1766463.3412795 chr19 57138057 N chr19 57138133 N DUP 12
SRR1766481.5417566 chr19 57138007 N chr19 57138134 N DUP 4
SRR1766448.10590751 chr19 57137994 N chr19 57138067 N DEL 2
SRR1766457.8388299 chr19 57137986 N chr19 57138130 N DUP 7
SRR1766442.35089032 chr19 57138028 N chr19 57138152 N DUP 12
SRR1766463.4717118 chr19 57138033 N chr19 57138098 N DEL 4
SRR1766453.8693804 chr19 57138038 N chr19 57138139 N DEL 6
SRR1766442.38839232 chr19 57138011 N chr19 57138242 N DUP 14
SRR1766470.9249561 chr19 57138052 N chr19 57138231 N DUP 15
SRR1766470.4003522 chr3 198168301 N chr3 198169088 N DEL 10
SRR1766467.3206215 chr3 198168361 N chr3 198168770 N DEL 5
SRR1766463.9035814 chr3 198168256 N chr3 198168411 N DUP 2
SRR1766443.9176099 chr3 198168293 N chr3 198169015 N DUP 3
SRR1766482.9253841 chr3 198168416 N chr3 198168888 N DEL 10
SRR1766486.5983349 chr3 198168324 N chr3 198169046 N DUP 12
SRR1766479.7923151 chr3 198168324 N chr3 198169046 N DUP 11
SRR1766480.1763470 chr3 198168320 N chr3 198169546 N DUP 5
SRR1766447.6382140 chr3 198168328 N chr3 198169050 N DUP 10
SRR1766473.4993679 chr3 198168364 N chr3 198168836 N DEL 15
SRR1766459.2845767 chr3 198168429 N chr3 198168838 N DEL 6
SRR1766482.9747560 chr3 198168406 N chr3 198168752 N DEL 23
SRR1766459.10979788 chr3 198168266 N chr3 198168484 N DUP 4
SRR1766468.5502777 chr3 198168486 N chr3 198168865 N DEL 5
SRR1766463.821138 chr3 198168513 N chr3 198169396 N DEL 5
SRR1766451.1827322 chr3 198168513 N chr3 198169396 N DEL 5
SRR1766464.7279379 chr3 198168513 N chr3 198169396 N DEL 5
SRR1766460.2885429 chr3 198168513 N chr3 198169396 N DEL 5
SRR1766450.4387738 chr3 198168562 N chr3 198168626 N DEL 5
SRR1766451.1147388 chr3 198168513 N chr3 198169396 N DEL 10
SRR1766442.2697693 chr3 198168513 N chr3 198169396 N DEL 10
SRR1766479.11570173 chr3 198168281 N chr3 198168625 N DUP 5
SRR1766475.2265742 chr3 198168562 N chr3 198168626 N DEL 5
SRR1766450.5701804 chr3 198168533 N chr3 198168595 N DUP 5
SRR1766447.11059853 chr3 198168533 N chr3 198168595 N DUP 5
SRR1766463.10014911 chr3 198168312 N chr3 198168532 N DEL 2
SRR1766464.4819138 chr3 198168595 N chr3 198168974 N DEL 5
SRR1766466.6705235 chr3 198168576 N chr3 198169396 N DEL 6
SRR1766458.8507277 chr3 198168595 N chr3 198169100 N DEL 10
SRR1766474.8032473 chr3 198168313 N chr3 198168533 N DEL 3
SRR1766474.8032473 chr3 198168533 N chr3 198168595 N DUP 5
SRR1766461.6124205 chr3 198168595 N chr3 198169415 N DEL 5
SRR1766470.1585656 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766462.2218794 chr3 198168595 N chr3 198169415 N DEL 5
SRR1766462.2847133 chr3 198169225 N chr3 198169415 N DEL 10
SRR1766454.7751465 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766449.1855363 chr3 198168595 N chr3 198169415 N DEL 5
SRR1766466.1238624 chr3 198168584 N chr3 198168898 N DUP 5
SRR1766458.149025 chr3 198168595 N chr3 198169415 N DEL 5
SRR1766476.3553924 chr3 198168533 N chr3 198168595 N DUP 5
SRR1766483.7964676 chr3 198168595 N chr3 198169415 N DEL 10
SRR1766466.1238624 chr3 198168533 N chr3 198168595 N DUP 5
SRR1766479.9453824 chr3 198168639 N chr3 198169396 N DEL 5
SRR1766450.8295568 chr3 198168639 N chr3 198169396 N DEL 5
SRR1766465.8869808 chr3 198168639 N chr3 198169396 N DEL 5
SRR1766442.7091515 chr3 198168626 N chr3 198168877 N DUP 5
SRR1766443.3857864 chr3 198168626 N chr3 198169129 N DUP 10
SRR1766455.3342924 chr3 198168646 N chr3 198168773 N DEL 5
SRR1766453.7421237 chr3 198168626 N chr3 198168877 N DUP 9
SRR1766457.6923399 chr3 198168689 N chr3 198168877 N DUP 5
SRR1766461.7582032 chr3 198168530 N chr3 198168783 N DEL 5
SRR1766475.2265742 chr3 198168532 N chr3 198168596 N DEL 5
SRR1766471.429066 chr3 198168562 N chr3 198168689 N DEL 5
SRR1766442.40805581 chr3 198168355 N chr3 198168701 N DEL 10
SRR1766464.8444301 chr3 198168292 N chr3 198168701 N DEL 10
SRR1766480.8407238 chr3 198168752 N chr3 198169129 N DUP 10
SRR1766481.10912235 chr3 198168521 N chr3 198168772 N DUP 5
SRR1766442.34123755 chr3 198168406 N chr3 198168752 N DEL 12
SRR1766454.5730456 chr3 198168521 N chr3 198168772 N DUP 5
SRR1766454.5089271 chr3 198168521 N chr3 198168772 N DUP 5
SRR1766478.8185470 chr3 198168752 N chr3 198168940 N DUP 10
SRR1766484.9415166 chr3 198168752 N chr3 198168940 N DUP 10
SRR1766452.2061604 chr3 198168772 N chr3 198168962 N DEL 5
SRR1766458.8145277 chr3 198168315 N chr3 198168724 N DEL 1
SRR1766466.3350993 chr3 198168802 N chr3 198169307 N DEL 9
SRR1766448.1998186 chr3 198168802 N chr3 198169307 N DEL 10
SRR1766454.684991 chr3 198168779 N chr3 198169410 N DEL 5
SRR1766450.6283041 chr3 198168432 N chr3 198168652 N DEL 5
SRR1766482.5096010 chr3 198168773 N chr3 198169150 N DUP 15
SRR1766442.25227893 chr3 198168773 N chr3 198169150 N DUP 15
SRR1766442.18645038 chr3 198168773 N chr3 198169150 N DUP 13
SRR1766475.5999820 chr3 198168511 N chr3 198168764 N DEL 3
SRR1766442.34274820 chr3 198168511 N chr3 198168764 N DEL 3
SRR1766445.4493860 chr3 198168773 N chr3 198169150 N DUP 11
SRR1766450.3427921 chr3 198168772 N chr3 198169403 N DEL 5
SRR1766477.1888262 chr3 198168898 N chr3 198169403 N DEL 9
SRR1766475.2686149 chr3 198168898 N chr3 198169403 N DEL 7
SRR1766448.4566268 chr3 198168772 N chr3 198169403 N DEL 5
SRR1766460.2252981 chr3 198168775 N chr3 198169152 N DUP 7
SRR1766470.8162279 chr3 198168776 N chr3 198169407 N DEL 5
SRR1766444.738799 chr3 198168780 N chr3 198169411 N DEL 5
SRR1766442.30573396 chr3 198168780 N chr3 198169411 N DEL 5
SRR1766452.2755246 chr3 198168815 N chr3 198168940 N DUP 5
SRR1766450.5701804 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766451.4579689 chr3 198168702 N chr3 198169396 N DEL 5
SRR1766442.23240159 chr3 198168688 N chr3 198169319 N DEL 15
SRR1766448.10026155 chr3 198168702 N chr3 198169396 N DEL 5
SRR1766448.578390 chr3 198168603 N chr3 198168793 N DEL 5
SRR1766486.5983349 chr3 198168420 N chr3 198168829 N DEL 10
SRR1766454.1401927 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766455.4999360 chr3 198169151 N chr3 198169528 N DUP 6
SRR1766471.1101035 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766442.8618175 chr3 198168428 N chr3 198168837 N DEL 10
SRR1766442.34414733 chr3 198168702 N chr3 198169396 N DEL 5
SRR1766465.4324141 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766444.6857119 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766455.6253367 chr3 198168428 N chr3 198168837 N DEL 10
SRR1766444.3699360 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766480.6787953 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766467.9442482 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766464.832250 chr3 198168591 N chr3 198169535 N DUP 10
SRR1766475.624834 chr3 198168639 N chr3 198169396 N DEL 5
SRR1766442.34604789 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766484.4291198 chr3 198168639 N chr3 198169396 N DEL 5
SRR1766477.7101214 chr3 198168815 N chr3 198169066 N DUP 10
SRR1766465.6269768 chr3 198168639 N chr3 198169396 N DEL 5
SRR1766446.4642990 chr3 198168595 N chr3 198168848 N DEL 10
SRR1766442.6537885 chr3 198168898 N chr3 198169151 N DEL 5
SRR1766485.776469 chr3 198168355 N chr3 198168827 N DEL 10
SRR1766471.2064196 chr3 198168353 N chr3 198168825 N DEL 10
SRR1766462.1723348 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766442.32097902 chr3 198168345 N chr3 198168817 N DEL 5
SRR1766442.46537276 chr3 198168345 N chr3 198168817 N DEL 5
SRR1766464.4819138 chr3 198168345 N chr3 198168817 N DEL 5
SRR1766463.7625470 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766482.3827695 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766470.420736 chr3 198168521 N chr3 198168898 N DUP 4
SRR1766473.1681528 chr3 198168848 N chr3 198168910 N DUP 10
SRR1766477.1343927 chr3 198168299 N chr3 198169525 N DUP 10
SRR1766485.12100895 chr3 198168836 N chr3 198168898 N DUP 10
SRR1766482.7183837 chr3 198168881 N chr3 198169071 N DEL 5
SRR1766459.1218682 chr3 198168888 N chr3 198169139 N DUP 10
SRR1766461.3325996 chr3 198168572 N chr3 198168825 N DEL 5
SRR1766479.7923151 chr3 198169093 N chr3 198169155 N DUP 5
SRR1766446.9440374 chr3 198168898 N chr3 198169088 N DEL 5
SRR1766486.246178 chr3 198168836 N chr3 198168898 N DUP 9
SRR1766469.9171054 chr3 198168372 N chr3 198168905 N DUP 4
SRR1766459.2845767 chr3 198168292 N chr3 198168951 N DUP 4
SRR1766484.4162833 chr3 198168794 N chr3 198169047 N DEL 10
SRR1766444.1157143 chr3 198168362 N chr3 198168895 N DUP 5
SRR1766452.9115284 chr3 198168802 N chr3 198168866 N DEL 3
SRR1766450.1379613 chr3 198168314 N chr3 198168849 N DEL 2
SRR1766472.2526073 chr3 198168762 N chr3 198168950 N DUP 10
SRR1766482.9253841 chr3 198168636 N chr3 198168950 N DUP 10
SRR1766452.6384526 chr3 198168762 N chr3 198168950 N DUP 10
SRR1766453.10082429 chr3 198168338 N chr3 198169186 N DUP 15
SRR1766463.182813 chr3 198168583 N chr3 198168899 N DEL 5
SRR1766453.10158119 chr3 198168978 N chr3 198169546 N DEL 2
SRR1766442.31879319 chr3 198168825 N chr3 198168950 N DUP 10
SRR1766452.1092783 chr3 198168522 N chr3 198168901 N DEL 5
SRR1766480.3685199 chr3 198168772 N chr3 198169088 N DEL 5
SRR1766457.1125682 chr3 198168825 N chr3 198168950 N DUP 2
SRR1766446.8889376 chr3 198168591 N chr3 198168907 N DEL 5
SRR1766454.6879471 chr3 198168513 N chr3 198168953 N DUP 10
SRR1766453.910504 chr3 198168310 N chr3 198168908 N DEL 5
SRR1766442.45189830 chr3 198168529 N chr3 198168908 N DEL 5
SRR1766480.4875857 chr3 198168513 N chr3 198168953 N DUP 5
SRR1766447.9921110 chr3 198168427 N chr3 198168836 N DEL 10
SRR1766462.4508420 chr3 198168580 N chr3 198168959 N DEL 10
SRR1766470.9600531 chr3 198168972 N chr3 198169288 N DEL 10
SRR1766477.9009449 chr3 198168961 N chr3 198169403 N DEL 5
SRR1766451.1147388 chr3 198168580 N chr3 198168959 N DEL 10
SRR1766449.9015426 chr3 198168991 N chr3 198169307 N DEL 5
SRR1766484.6834473 chr3 198168991 N chr3 198169307 N DEL 5
SRR1766483.1634676 chr3 198169013 N chr3 198169140 N DEL 5
SRR1766479.12862958 chr3 198169035 N chr3 198169288 N DEL 5
SRR1766451.10354665 chr3 198168314 N chr3 198168975 N DEL 2
SRR1766484.4352583 chr3 198168594 N chr3 198169288 N DEL 5
SRR1766442.14859936 chr3 198169063 N chr3 198169566 N DUP 5
SRR1766480.3509420 chr3 198169053 N chr3 198169432 N DEL 5
SRR1766452.1424623 chr3 198169224 N chr3 198169288 N DEL 10
SRR1766459.7820729 chr3 198168594 N chr3 198169288 N DEL 5
SRR1766445.9260066 chr3 198168555 N chr3 198169058 N DUP 1
SRR1766449.3403725 chr3 198169047 N chr3 198169487 N DUP 5
SRR1766486.147745 chr3 198168594 N chr3 198169288 N DEL 9
SRR1766457.503391 chr3 198168428 N chr3 198168837 N DEL 10
SRR1766469.2879404 chr3 198169046 N chr3 198169425 N DEL 5
SRR1766443.1188513 chr3 198169046 N chr3 198169425 N DEL 5
SRR1766448.2303111 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766453.1085413 chr3 198169047 N chr3 198169487 N DUP 5
SRR1766474.2192381 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766478.11096723 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766475.4682199 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766473.4683580 chr3 198169048 N chr3 198169362 N DUP 10
SRR1766468.2547939 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766486.7845216 chr3 198169047 N chr3 198169361 N DUP 10
SRR1766469.10805515 chr3 198168335 N chr3 198168996 N DEL 1
SRR1766450.4387738 chr3 198169047 N chr3 198169487 N DUP 5
SRR1766464.9935684 chr3 198169047 N chr3 198169487 N DUP 5
SRR1766459.3172453 chr3 198168594 N chr3 198169288 N DEL 5
SRR1766454.6879471 chr3 198169369 N chr3 198169433 N DEL 9
SRR1766449.3403725 chr3 198169369 N chr3 198169433 N DEL 10
SRR1766473.9311745 chr3 198169055 N chr3 198169117 N DUP 10
SRR1766442.16936494 chr3 198168794 N chr3 198169047 N DEL 10
SRR1766453.5629003 chr3 198168513 N chr3 198168890 N DUP 5
SRR1766474.7853394 chr3 198168668 N chr3 198169047 N DEL 5
SRR1766447.3271600 chr3 198168668 N chr3 198169047 N DEL 5
SRR1766448.4465461 chr3 198168668 N chr3 198169047 N DEL 5
SRR1766475.8232298 chr3 198168668 N chr3 198169047 N DEL 5
SRR1766451.7300931 chr3 198168921 N chr3 198169046 N DUP 5
SRR1766471.2197121 chr3 198168668 N chr3 198169047 N DEL 5
SRR1766459.9461813 chr3 198168668 N chr3 198169047 N DEL 5
SRR1766469.8352623 chr3 198168513 N chr3 198169079 N DUP 5
SRR1766458.8507277 chr3 198168676 N chr3 198169055 N DEL 10
SRR1766464.5011680 chr3 198169180 N chr3 198169433 N DEL 9
SRR1766446.2005536 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766442.37051932 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766462.8845260 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766459.7820729 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766478.8149081 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766448.10141482 chr3 198168762 N chr3 198168950 N DUP 10
SRR1766443.3217929 chr3 198168394 N chr3 198169055 N DEL 10
SRR1766442.5783748 chr3 198168762 N chr3 198168950 N DUP 10
SRR1766465.9837079 chr3 198169117 N chr3 198169307 N DEL 5
SRR1766443.7510034 chr3 198168457 N chr3 198169055 N DEL 10
SRR1766457.8951768 chr3 198168393 N chr3 198169054 N DEL 5
SRR1766475.9502882 chr3 198169117 N chr3 198169307 N DEL 5
SRR1766456.619137 chr3 198169055 N chr3 198169180 N DUP 5
SRR1766445.3857965 chr3 198168625 N chr3 198169067 N DEL 5
SRR1766467.4594022 chr3 198168395 N chr3 198169056 N DEL 10
SRR1766470.11000823 chr3 198169059 N chr3 198169184 N DUP 3
SRR1766479.810973 chr3 198168398 N chr3 198169059 N DEL 8
SRR1766452.380541 chr3 198169060 N chr3 198169185 N DUP 2
SRR1766442.9264084 chr3 198168825 N chr3 198168950 N DUP 5
SRR1766460.4744481 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766484.9025942 chr3 198169117 N chr3 198169307 N DEL 5
SRR1766446.9440374 chr3 198169098 N chr3 198169288 N DEL 10
SRR1766450.6116059 chr3 198169098 N chr3 198169288 N DEL 10
SRR1766465.10534219 chr3 198169098 N chr3 198169288 N DEL 10
SRR1766482.11356723 chr3 198169117 N chr3 198169307 N DEL 5
SRR1766459.1218682 chr3 198168344 N chr3 198169068 N DEL 2
SRR1766460.4744481 chr3 198168843 N chr3 198168905 N DUP 10
SRR1766460.9798777 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766470.4827455 chr3 198168825 N chr3 198169139 N DUP 5
SRR1766464.3904924 chr3 198169078 N chr3 198169142 N DEL 5
SRR1766466.1909684 chr3 198168332 N chr3 198169180 N DUP 2
SRR1766479.9645029 chr3 198169077 N chr3 198169139 N DUP 2
SRR1766442.14859936 chr3 198169124 N chr3 198169375 N DUP 5
SRR1766453.10082429 chr3 198168900 N chr3 198169090 N DEL 5
SRR1766442.9781420 chr3 198168353 N chr3 198169077 N DEL 5
SRR1766464.9935684 chr3 198168992 N chr3 198169369 N DUP 5
SRR1766457.3720400 chr3 198169140 N chr3 198169517 N DUP 5
SRR1766446.10204673 chr3 198168898 N chr3 198169088 N DEL 5
SRR1766454.9378363 chr3 198168992 N chr3 198169369 N DUP 5
SRR1766477.10850804 chr3 198168260 N chr3 198169077 N DEL 5
SRR1766444.6298511 chr3 198168825 N chr3 198168950 N DUP 10
SRR1766484.2970205 chr3 198168825 N chr3 198168950 N DUP 10
SRR1766449.1855363 chr3 198168825 N chr3 198169139 N DUP 5
SRR1766451.10354665 chr3 198168992 N chr3 198169369 N DUP 5
SRR1766455.4999360 chr3 198168992 N chr3 198169369 N DUP 5
SRR1766454.870693 chr3 198168365 N chr3 198169150 N DUP 6
SRR1766482.11356723 chr3 198168992 N chr3 198169369 N DUP 5
SRR1766442.19270100 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766442.46920417 chr3 198168513 N chr3 198169142 N DUP 5
SRR1766442.12012906 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766470.7841674 chr3 198168772 N chr3 198169088 N DEL 5
SRR1766454.4115906 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766450.9303779 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766456.4679184 chr3 198168513 N chr3 198169142 N DUP 5
SRR1766469.1169436 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766454.7751465 chr3 198168992 N chr3 198169369 N DUP 5
SRR1766473.1681528 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766451.5914311 chr3 198168513 N chr3 198169142 N DUP 5
SRR1766453.1680305 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766479.13019236 chr3 198168825 N chr3 198168950 N DUP 10
SRR1766464.7672523 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766445.9276662 chr3 198168774 N chr3 198169090 N DEL 5
SRR1766460.7941418 chr3 198168774 N chr3 198169090 N DEL 5
SRR1766464.9399280 chr3 198168513 N chr3 198169142 N DUP 5
SRR1766455.2914168 chr3 198168515 N chr3 198168892 N DUP 5
SRR1766486.147745 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766467.10458266 chr3 198168975 N chr3 198169163 N DUP 1
SRR1766444.738799 chr3 198168775 N chr3 198169091 N DEL 5
SRR1766466.2502959 chr3 198168513 N chr3 198169142 N DUP 5
SRR1766453.6561226 chr3 198168958 N chr3 198169148 N DEL 10
SRR1766445.9260066 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766455.7254789 chr3 198168514 N chr3 198169143 N DUP 5
SRR1766464.3904924 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766473.7100442 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766450.5785015 chr3 198169143 N chr3 198169396 N DEL 7
SRR1766450.8295568 chr3 198168887 N chr3 198169140 N DEL 5
SRR1766454.6331897 chr3 198168513 N chr3 198169142 N DUP 5
SRR1766451.5885465 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766455.3342924 chr3 198168572 N chr3 198169140 N DEL 5
SRR1766471.9903279 chr3 198168815 N chr3 198169192 N DUP 6
SRR1766457.3720400 chr3 198168594 N chr3 198169288 N DEL 9
SRR1766442.22748149 chr3 198168513 N chr3 198168953 N DUP 9
SRR1766453.6561226 chr3 198168594 N chr3 198169288 N DEL 7
SRR1766460.5977806 chr3 198168594 N chr3 198169288 N DEL 6
SRR1766467.5880320 chr3 198168572 N chr3 198169140 N DEL 5
SRR1766454.9378363 chr3 198168594 N chr3 198169288 N DEL 6
SRR1766442.13409660 chr3 198168420 N chr3 198169396 N DEL 10
SRR1766453.10136296 chr3 198168418 N chr3 198168638 N DEL 10
SRR1766470.6730709 chr3 198168613 N chr3 198169055 N DEL 10
SRR1766484.9748975 chr3 198168357 N chr3 198169396 N DEL 10
SRR1766483.10467038 chr3 198168594 N chr3 198169288 N DEL 5
SRR1766447.10449885 chr3 198168420 N chr3 198169396 N DEL 10
SRR1766486.3461517 chr3 198169047 N chr3 198169172 N DUP 9
SRR1766466.2801333 chr3 198168416 N chr3 198168825 N DEL 10
SRR1766442.28744001 chr3 198169181 N chr3 198169495 N DUP 10
SRR1766442.27572363 chr3 198168418 N chr3 198168638 N DEL 10
SRR1766446.8068417 chr3 198169047 N chr3 198169172 N DUP 10
SRR1766445.2284530 chr3 198168866 N chr3 198169180 N DUP 15
SRR1766459.1534905 chr3 198168572 N chr3 198169140 N DEL 5
SRR1766471.747624 chr3 198169047 N chr3 198169172 N DUP 10
SRR1766473.7100442 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766479.6955620 chr3 198169047 N chr3 198169172 N DUP 10
SRR1766486.1130915 chr3 198169047 N chr3 198169172 N DUP 10
SRR1766451.5914311 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766473.6114207 chr3 198168550 N chr3 198169242 N DUP 2
SRR1766472.2095336 chr3 198169180 N chr3 198169433 N DEL 15
SRR1766460.9485661 chr3 198168865 N chr3 198169242 N DUP 5
SRR1766447.9827794 chr3 198168497 N chr3 198169252 N DUP 10
SRR1766465.671698 chr3 198169369 N chr3 198169433 N DEL 13
SRR1766466.2502959 chr3 198168513 N chr3 198169205 N DUP 10
SRR1766469.185018 chr3 198168676 N chr3 198169181 N DEL 5
SRR1766461.6124205 chr3 198168550 N chr3 198169181 N DEL 5
SRR1766485.9932434 chr3 198168394 N chr3 198169181 N DEL 5
SRR1766449.6993317 chr3 198169151 N chr3 198169276 N DUP 5
SRR1766448.1998186 chr3 198168396 N chr3 198169183 N DEL 5
SRR1766481.9241269 chr3 198169226 N chr3 198169351 N DUP 5
SRR1766481.10912235 chr3 198169036 N chr3 198169226 N DEL 10
SRR1766466.1909684 chr3 198169099 N chr3 198169226 N DEL 5
SRR1766448.578390 chr3 198168638 N chr3 198169206 N DEL 2
SRR1766450.10028515 chr3 198169151 N chr3 198169276 N DUP 5
SRR1766484.4291198 chr3 198168612 N chr3 198169243 N DEL 5
SRR1766454.5089271 chr3 198168549 N chr3 198169243 N DEL 10
SRR1766478.8688477 chr3 198168549 N chr3 198169243 N DEL 10
SRR1766450.6135126 chr3 198168320 N chr3 198169233 N DEL 5
SRR1766479.3581095 chr3 198168909 N chr3 198169288 N DEL 12
SRR1766465.1965398 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766452.2248917 chr3 198168909 N chr3 198169288 N DEL 15
SRR1766459.4870445 chr3 198168594 N chr3 198169288 N DEL 10
SRR1766476.8882488 chr3 198168928 N chr3 198169307 N DEL 15
SRR1766467.5347130 chr3 198168531 N chr3 198169288 N DEL 5
SRR1766477.9288504 chr3 198168802 N chr3 198169307 N DEL 15
SRR1766458.2705722 chr3 198168588 N chr3 198169282 N DEL 5
SRR1766461.4066443 chr3 198168571 N chr3 198169389 N DUP 5
SRR1766460.8661718 chr3 198168676 N chr3 198169307 N DEL 15
SRR1766442.34414733 chr3 198168783 N chr3 198169288 N DEL 5
SRR1766450.252618 chr3 198169140 N chr3 198169328 N DUP 10
SRR1766442.23240159 chr3 198168394 N chr3 198169307 N DEL 10
SRR1766446.10204673 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766459.4870445 chr3 198168815 N chr3 198169192 N DUP 10
SRR1766478.10398491 chr3 198168386 N chr3 198169299 N DEL 4
SRR1766466.1988026 chr3 198168389 N chr3 198169302 N DEL 1
SRR1766460.5977806 chr3 198169224 N chr3 198169288 N DEL 14
SRR1766443.1207970 chr3 198169047 N chr3 198169361 N DUP 10
SRR1766443.1207970 chr3 198169047 N chr3 198169361 N DUP 5
SRR1766447.3271600 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766464.1224651 chr3 198168394 N chr3 198169307 N DEL 5
SRR1766449.9644855 chr3 198169047 N chr3 198169361 N DUP 10
SRR1766448.391205 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766453.1085413 chr3 198169224 N chr3 198169288 N DEL 15
SRR1766474.2192381 chr3 198169224 N chr3 198169288 N DEL 15
SRR1766442.38264626 chr3 198169224 N chr3 198169288 N DEL 15
SRR1766452.1424623 chr3 198169224 N chr3 198169288 N DEL 13
SRR1766442.12012906 chr3 198168866 N chr3 198169369 N DUP 15
SRR1766473.572903 chr3 198168345 N chr3 198169321 N DEL 1
SRR1766465.6269768 chr3 198168823 N chr3 198169389 N DUP 5
SRR1766465.10534219 chr3 198169369 N chr3 198169433 N DEL 10
SRR1766442.27618723 chr3 198168823 N chr3 198169389 N DUP 5
SRR1766479.10326344 chr3 198169180 N chr3 198169433 N DEL 15
SRR1766449.9644855 chr3 198169369 N chr3 198169433 N DEL 7
SRR1766461.2947535 chr3 198169369 N chr3 198169433 N DEL 10
SRR1766443.3745812 chr3 198169369 N chr3 198169433 N DEL 7
SRR1766455.8789366 chr3 198168668 N chr3 198169047 N DEL 5
SRR1766474.11583667 chr3 198168668 N chr3 198169047 N DEL 5
SRR1766463.182813 chr3 198168676 N chr3 198169370 N DEL 5
SRR1766479.9714261 chr3 198168676 N chr3 198169370 N DEL 5
SRR1766443.10162366 chr3 198168992 N chr3 198169369 N DUP 5
SRR1766459.1759401 chr3 198168626 N chr3 198169192 N DUP 12
SRR1766459.10902306 chr3 198169140 N chr3 198169202 N DUP 10
SRR1766464.5484446 chr3 198168889 N chr3 198169394 N DEL 10
SRR1766475.1988528 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766452.10032623 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766452.10032623 chr3 198169224 N chr3 198169288 N DEL 12
SRR1766477.10850804 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766442.33436551 chr3 198169224 N chr3 198169288 N DEL 15
SRR1766486.1810069 chr3 198169224 N chr3 198169288 N DEL 13
SRR1766445.54561 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766447.1649448 chr3 198169206 N chr3 198169396 N DEL 10
SRR1766483.6483256 chr3 198168829 N chr3 198169395 N DUP 5
SRR1766461.2947535 chr3 198169224 N chr3 198169288 N DEL 10
SRR1766474.3597978 chr3 198168394 N chr3 198169370 N DEL 5
SRR1766456.3346227 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766478.10155535 chr3 198168959 N chr3 198169462 N DUP 5
SRR1766472.7814779 chr3 198168829 N chr3 198169395 N DUP 5
SRR1766444.3699360 chr3 198168829 N chr3 198169395 N DUP 5
SRR1766469.7577147 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766472.10629820 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766448.391205 chr3 198168829 N chr3 198169395 N DUP 5
SRR1766465.266139 chr3 198169200 N chr3 198169390 N DEL 5
SRR1766452.4383822 chr3 198168626 N chr3 198169192 N DUP 10
SRR1766467.9003657 chr3 198169080 N chr3 198169396 N DEL 10
SRR1766463.1766669 chr3 198168823 N chr3 198169389 N DUP 10
SRR1766442.22820724 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766466.11183284 chr3 198168343 N chr3 198169382 N DEL 1
SRR1766464.7279379 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766479.9714261 chr3 198168351 N chr3 198169390 N DEL 7
SRR1766451.9781443 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766466.8926755 chr3 198168351 N chr3 198169390 N DEL 5
SRR1766451.6884696 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766452.1509551 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766470.5199415 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766479.3818572 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766443.7224086 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766469.8352623 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766475.4068630 chr3 198168825 N chr3 198169139 N DUP 5
SRR1766473.2918984 chr3 198168294 N chr3 198169396 N DEL 11
SRR1766461.1662885 chr3 198168575 N chr3 198169395 N DEL 5
SRR1766473.6114207 chr3 198168297 N chr3 198169399 N DEL 11
SRR1766474.3597978 chr3 198168513 N chr3 198169457 N DUP 1
SRR1766442.34082399 chr3 198168295 N chr3 198169397 N DEL 14
SRR1766454.6331897 chr3 198168295 N chr3 198169397 N DEL 14
SRR1766480.4875857 chr3 198168513 N chr3 198168890 N DUP 10
SRR1766463.6602952 chr3 198168581 N chr3 198169401 N DEL 9
SRR1766442.47182058 chr3 198168513 N chr3 198169457 N DUP 5
SRR1766461.1662885 chr3 198168853 N chr3 198168915 N DUP 1
SRR1766464.5484446 chr3 198168762 N chr3 198168950 N DUP 6
SRR1766481.6445683 chr3 198168584 N chr3 198168774 N DEL 5
SRR1766454.3656345 chr3 198168513 N chr3 198169457 N DUP 5
SRR1766459.3172453 chr3 198168513 N chr3 198168890 N DUP 9
SRR1766460.9485661 chr3 198168676 N chr3 198169055 N DEL 10
SRR1766461.828113 chr3 198168513 N chr3 198168890 N DUP 9
SRR1766466.8926755 chr3 198168291 N chr3 198169517 N DUP 5
SRR1766482.659967 chr3 198168513 N chr3 198168890 N DUP 9
SRR1766484.9748975 chr3 198168291 N chr3 198169517 N DUP 5
SRR1766451.9039239 chr3 198168588 N chr3 198168778 N DEL 3
SRR1766442.45189830 chr3 198168825 N chr3 198169139 N DUP 7
SRR1766450.3205339 chr3 198169180 N chr3 198169433 N DEL 13
SRR1766472.3204706 chr3 198168842 N chr3 198168904 N DUP 5
SRR1766443.10162366 chr3 198168594 N chr3 198169414 N DEL 4
SRR1766449.1687252 chr3 198168836 N chr3 198168898 N DUP 9
SRR1766449.10184815 chr3 198168780 N chr3 198169411 N DEL 5
SRR1766452.9769942 chr3 198169369 N chr3 198169433 N DEL 10
SRR1766457.1125682 chr3 198168824 N chr3 198169201 N DUP 9
SRR1766473.6968027 chr3 198168898 N chr3 198168962 N DEL 10
SRR1766475.5999820 chr3 198168576 N chr3 198169396 N DEL 5
SRR1766481.943450 chr3 198169046 N chr3 198169425 N DEL 5
SRR1766448.4465461 chr3 198168576 N chr3 198169396 N DEL 6
SRR1766446.8889376 chr3 198168595 N chr3 198168974 N DEL 5
SRR1766450.9303779 chr3 198168576 N chr3 198169396 N DEL 7
SRR1766454.684991 chr3 198168562 N chr3 198168815 N DEL 2
SRR1766448.4054466 chr3 198168689 N chr3 198169192 N DUP 9
SRR1766482.2232758 chr3 198168576 N chr3 198169396 N DEL 9
SRR1766481.7178966 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766442.8103666 chr3 198168310 N chr3 198169412 N DEL 6
SRR1766450.10028515 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766446.9974041 chr3 198168410 N chr3 198168819 N DEL 5
SRR1766447.433975 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766474.8529549 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766453.6544433 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766461.6468289 chr3 198168576 N chr3 198169396 N DEL 10
SRR1766473.4683580 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766474.9001137 chr3 198168866 N chr3 198169180 N DUP 5
SRR1766485.4680483 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766462.8845260 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766455.3401312 chr3 198169050 N chr3 198169429 N DEL 5
SRR1766459.9461813 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766442.9781420 chr3 198168406 N chr3 198168815 N DEL 5
SRR1766467.10458266 chr3 198168866 N chr3 198169369 N DUP 10
SRR1766464.1224651 chr3 198168343 N chr3 198168815 N DEL 5
SRR1766449.6993317 chr3 198168343 N chr3 198168815 N DEL 5
SRR1766452.2023421 chr3 198169307 N chr3 198169495 N DUP 10
SRR1766453.3870843 chr3 198168343 N chr3 198168815 N DEL 5
SRR1766477.9288504 chr3 198168815 N chr3 198169066 N DUP 8
SRR1766445.3058538 chr3 198169117 N chr3 198169307 N DEL 7
SRR1766475.9242745 chr3 198168576 N chr3 198169396 N DEL 5
SRR1766453.5629003 chr3 198168583 N chr3 198169529 N DEL 5
SRR1766446.2336999 chr10 101730845 N chr10 101731152 N DUP 5
SRR1766442.7859557 chr10 101730848 N chr10 101731155 N DUP 2
SRR1766479.8333017 chr10 101730849 N chr10 101731155 N DUP 2
SRR1766476.8469361 chr10 101731102 N chr10 101731411 N DEL 1
SRR1766482.8035956 chr12 129388154 N chr12 129388238 N DEL 5
SRR1766466.2235694 chr12 129388109 N chr12 129388274 N DUP 5
SRR1766442.23051347 chr12 129388109 N chr12 129388191 N DUP 5
SRR1766473.10023952 chr12 129388211 N chr12 129388295 N DEL 5
SRR1766469.5921891 chr12 129388159 N chr12 129388241 N DUP 5
SRR1766456.790203 chr12 129388084 N chr12 129388168 N DEL 6
SRR1766448.622219 chr12 129388110 N chr12 129388275 N DUP 8
SRR1766455.5441327 chr12 129388142 N chr12 129388226 N DEL 9
SRR1766445.5448984 chr12 129388085 N chr12 129388169 N DEL 5
SRR1766450.10181560 chr12 129388109 N chr12 129388274 N DUP 5
SRR1766484.2144915 chr12 129388110 N chr12 129388275 N DUP 10
SRR1766471.10932933 chr12 129388132 N chr12 129388297 N DUP 2
SRR1766481.855447 chr12 129388132 N chr12 129388297 N DUP 4
SRR1766460.4324622 chr12 129388060 N chr12 129388308 N DUP 5
SRR1766442.36291067 chr12 129388060 N chr12 129388142 N DUP 5
SRR1766464.10054632 chr12 129388060 N chr12 129388308 N DUP 5
SRR1766460.616440 chr5 149226090 N chr5 149226178 N DEL 5
SRR1766467.1530237 chr2 88012368 N chr2 88012675 N DUP 5
SRR1766459.5794712 chr11 16888060 N chr11 16888294 N DEL 4
SRR1766446.3306 chr19 55630951 N chr19 55631130 N DEL 4
SRR1766457.6837236 chr19 55630951 N chr19 55631130 N DEL 4
SRR1766485.8172498 chr19 47802745 N chr19 47802842 N DEL 6
SRR1766466.10585236 chr19 47802655 N chr19 47802708 N DUP 5
SRR1766463.5850450 chr19 47802684 N chr19 47802767 N DUP 5
SRR1766474.1605081 chr19 47802619 N chr19 47802734 N DEL 9
SRR1766442.29120378 chr19 47802575 N chr19 47802756 N DEL 3
SRR1766482.2166763 chr19 47802706 N chr19 47802815 N DEL 12
SRR1766450.1557372 chr19 47802544 N chr19 47802839 N DEL 5
SRR1766463.3898758 chr19 47802679 N chr19 47802842 N DEL 5
SRR1766465.10994267 chr11 59632741 N chr11 59632802 N DUP 8
SRR1766463.7577776 chr11 59632741 N chr11 59632802 N DUP 8
SRR1766452.1172948 chr11 59632741 N chr11 59632802 N DUP 10
SRR1766472.11009848 chr11 59632741 N chr11 59632802 N DUP 11
SRR1766442.31034937 chr11 59632741 N chr11 59632802 N DUP 11
SRR1766479.2848175 chr11 59632741 N chr11 59632802 N DUP 11
SRR1766450.635471 chr11 59632741 N chr11 59632810 N DUP 5
SRR1766443.4708134 chr11 59632741 N chr11 59632810 N DUP 8
SRR1766475.3515252 chr11 59632733 N chr11 59632862 N DUP 6
SRR1766442.15789467 chr11 59632758 N chr11 59632896 N DUP 3
SRR1766447.4691360 chr11 59632758 N chr11 59632896 N DUP 3
SRR1766452.617377 chr11 59632758 N chr11 59632896 N DUP 5
SRR1766475.7201960 chr11 59632758 N chr11 59632896 N DUP 7
SRR1766460.2572116 chr11 59632758 N chr11 59632896 N DUP 9
SRR1766462.1996609 chr11 59632758 N chr11 59632896 N DUP 4
SRR1766446.1282549 chr11 59632758 N chr11 59632896 N DUP 5
SRR1766456.1667761 chr11 59632758 N chr11 59632896 N DUP 5
SRR1766454.7510045 chr11 59632758 N chr11 59632896 N DUP 11
SRR1766453.10320305 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766450.7426073 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766464.8162357 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766449.2984884 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766475.10377551 chr11 59632745 N chr11 59632905 N DUP 10
SRR1766472.11075332 chr11 59632758 N chr11 59632896 N DUP 17
SRR1766447.891614 chr11 59632758 N chr11 59632896 N DUP 10
SRR1766451.1611213 chr11 59632758 N chr11 59632896 N DUP 11
SRR1766476.6201423 chr11 59632758 N chr11 59632896 N DUP 14
SRR1766465.8666844 chr11 59632758 N chr11 59632896 N DUP 14
SRR1766468.526664 chr11 59632752 N chr11 59632817 N DEL 7
SRR1766461.4250550 chr11 59632752 N chr11 59632819 N DEL 5
SRR1766443.6420253 chr11 59632779 N chr11 59632848 N DEL 2
SRR1766450.71018 chr11 59632780 N chr11 59632849 N DEL 1
SRR1766479.5032663 chr11 59632755 N chr11 59632897 N DEL 15
SRR1766461.10365712 chr11 59632747 N chr11 59632903 N DEL 9
SRR1766442.36269242 chr11 59632749 N chr11 59632905 N DEL 7
SRR1766442.2571777 chr11 59632782 N chr11 59632912 N DEL 6
SRR1766465.6828250 chr11 59632776 N chr11 59632906 N DEL 6
SRR1766455.7866531 chr11 59632759 N chr11 59632911 N DEL 1
SRR1766447.2500321 chr11 59632759 N chr11 59632911 N DEL 1
SRR1766473.10277643 chr11 59632780 N chr11 59632910 N DEL 2
SRR1766443.1565522 chr10 27443056 N chr10 27443130 N DUP 8
SRR1766457.2999084 chr10 1160912 N chr10 1161025 N DUP 1
SRR1766464.10648971 chr10 132055033 N chr10 132055170 N DUP 1
SRR1766480.2696508 chr10 132055067 N chr10 132055158 N DUP 5
SRR1766460.1192209 chr14 91044488 N chr14 91044543 N DEL 1
SRR1766459.7519141 chr14 91044491 N chr14 91044542 N DEL 17
SRR1766484.11474737 chr1 81747030 N chr1 81747113 N DEL 14
SRR1766458.55022 chr1 231733659 N chr1 231733732 N DEL 7
SRR1766460.2202570 chr1 231733668 N chr1 231733741 N DEL 8
SRR1766463.1005663 chr1 231733473 N chr1 231733616 N DEL 3
SRR1766480.2312389 chr1 231733413 N chr1 231733613 N DEL 5
SRR1766475.8965645 chr14 104325061 N chr14 104325190 N DUP 10
SRR1766442.39536390 chr14 104325087 N chr14 104325216 N DUP 5
SRR1766477.1099365 chr14 104325126 N chr14 104325191 N DUP 14
SRR1766455.4718250 chr14 104325139 N chr14 104325266 N DUP 1
SRR1766449.5620478 chr14 104325139 N chr14 104325266 N DUP 10
SRR1766466.8296672 chr14 104325139 N chr14 104325266 N DUP 10
SRR1766442.8660600 chr14 104325139 N chr14 104325266 N DUP 10
SRR1766479.12956037 chr14 104325140 N chr14 104325267 N DUP 10
SRR1766465.3677512 chr14 104325124 N chr14 104325213 N DEL 6
SRR1766459.971536 chr14 104325247 N chr14 104325312 N DUP 1
SRR1766442.28702323 chr21 14261869 N chr21 14261948 N DEL 5
SRR1766475.6067563 chr21 14261869 N chr21 14261948 N DEL 5
SRR1766481.323076 chr21 14261869 N chr21 14261948 N DEL 5
SRR1766461.7271949 chr21 14261869 N chr21 14261948 N DEL 5
SRR1766454.8861020 chr21 14261869 N chr21 14261948 N DEL 5
SRR1766463.1337243 chr21 14261869 N chr21 14261948 N DEL 5
SRR1766479.4725377 chr21 14261869 N chr21 14261948 N DEL 5
SRR1766455.671730 chr21 14261871 N chr21 14261948 N DUP 1
SRR1766451.6949817 chr21 14261871 N chr21 14261948 N DUP 5
SRR1766445.760832 chr21 14261871 N chr21 14261948 N DUP 5
SRR1766459.2284506 chr21 14261871 N chr21 14261948 N DUP 5
SRR1766442.9005132 chr21 14261871 N chr21 14261948 N DUP 13
SRR1766443.5580810 chr21 14261873 N chr21 14261950 N DUP 13
SRR1766446.1585090 chr21 14261873 N chr21 14261950 N DUP 13
SRR1766449.1360291 chr21 14261871 N chr21 14261948 N DUP 13
SRR1766474.8544762 chr21 14261874 N chr21 14261951 N DUP 12
SRR1766460.18178 chr21 14261872 N chr21 14261949 N DUP 14
SRR1766452.6758425 chr21 14261871 N chr21 14261948 N DUP 17
SRR1766485.11016921 chr21 14261871 N chr21 14261948 N DUP 18
SRR1766447.9259204 chr21 14261871 N chr21 14261948 N DUP 23
SRR1766475.132202 chr19 6343693 N chr19 6343810 N DUP 5
SRR1766451.8352191 chr19 6343617 N chr19 6343739 N DEL 8
SRR1766479.1666874 chr19 33506268 N chr19 33506566 N DUP 5
SRR1766484.9732498 chr19 33506281 N chr19 33506482 N DUP 1
SRR1766459.5278527 chr19 33506281 N chr19 33506482 N DUP 3
SRR1766457.675379 chr19 33506390 N chr19 33506493 N DUP 5
SRR1766468.6198411 chr19 33506491 N chr19 33506589 N DEL 5
SRR1766484.7065748 chr19 33506497 N chr19 33506595 N DEL 5
SRR1766464.9266769 chr19 33506311 N chr19 33506410 N DEL 4
SRR1766484.5426429 chr19 33506497 N chr19 33506595 N DEL 7
SRR1766486.8632295 chr19 33506599 N chr19 33506783 N DUP 5
SRR1766473.6475918 chr4 4219978 N chr4 4220223 N DEL 2
SRR1766461.858923 chr4 4220141 N chr4 4220206 N DEL 2
SRR1766442.41054206 chr4 4220180 N chr4 4220245 N DUP 14
SRR1766452.7690436 chr4 4219993 N chr4 4220202 N DEL 7
SRR1766448.912489 chr4 4219964 N chr4 4220213 N DEL 2
SRR1766461.3961946 chr3 11057696 N chr3 11057861 N DUP 5
SRR1766462.10518422 chrX 649100 N chrX 649153 N DEL 10
SRR1766446.10003 chrX 649094 N chrX 649167 N DUP 11
SRR1766481.7302533 chrX 649071 N chrX 649196 N DEL 11
SRR1766464.6320556 chrX 649077 N chrX 649202 N DEL 6
SRR1766479.2828963 chrX 649080 N chrX 649205 N DEL 3
SRR1766484.5494232 chr2 30263826 N chr2 30264145 N DEL 1
SRR1766448.10642261 chr2 30263892 N chr2 30264211 N DEL 10
SRR1766466.7746883 chr21 45501807 N chr21 45502023 N DEL 2
SRR1766479.11284121 chr21 45501807 N chr21 45502023 N DEL 4
SRR1766458.2690898 chr21 45501821 N chr21 45501951 N DEL 1
SRR1766463.6131966 chr21 45501821 N chr21 45501951 N DEL 1
SRR1766476.4692302 chr21 45501821 N chr21 45501951 N DEL 9
SRR1766467.2321013 chr21 45501821 N chr21 45501951 N DEL 9
SRR1766471.7340057 chr21 45501821 N chr21 45501951 N DEL 9
SRR1766485.10433661 chr21 45501821 N chr21 45501951 N DEL 10
SRR1766480.8242211 chr21 45501849 N chr21 45502109 N DEL 5
SRR1766449.2761965 chr21 45501821 N chr21 45501951 N DEL 10
SRR1766460.4391164 chr21 45501797 N chr21 45501883 N DUP 7
SRR1766475.1586005 chr21 45501821 N chr21 45501951 N DEL 10
SRR1766454.7234472 chr21 45501849 N chr21 45502109 N DEL 5
SRR1766464.8914009 chr21 45501864 N chr21 45501951 N DEL 3
SRR1766462.5933631 chr21 45501821 N chr21 45501951 N DEL 10
SRR1766478.7185330 chr21 45501935 N chr21 45502109 N DEL 6
SRR1766449.10881995 chr21 45501840 N chr21 45502097 N DUP 10
SRR1766470.3741626 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766469.4529495 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766442.33116854 chr21 45502086 N chr21 45502218 N DEL 22
SRR1766468.5392343 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766465.5211463 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766481.187727 chr21 45501802 N chr21 45502102 N DUP 10
SRR1766469.8292411 chr21 45501864 N chr21 45501951 N DEL 5
SRR1766442.37980265 chr21 45501864 N chr21 45501951 N DEL 5
SRR1766469.3093661 chr21 45501821 N chr21 45501951 N DEL 5
SRR1766462.792828 chr21 45501821 N chr21 45501951 N DEL 5
SRR1766442.6124986 chr21 45501822 N chr21 45501952 N DEL 5
SRR1766476.1237475 chr21 45501822 N chr21 45501952 N DEL 5
SRR1766449.1035916 chr21 45501824 N chr21 45501954 N DEL 5
SRR1766484.6914247 chr21 45501831 N chr21 45501961 N DEL 5
SRR1766482.6656983 chr21 45501832 N chr21 45501962 N DEL 4
SRR1766455.1198918 chr21 45501808 N chr21 45502022 N DUP 3
SRR1766455.5073324 chr21 45501808 N chr21 45502022 N DUP 3
SRR1766455.9740757 chr21 45501808 N chr21 45502022 N DUP 5
SRR1766442.35278987 chr21 45501808 N chr21 45502022 N DUP 14
SRR1766462.884109 chr21 45501990 N chr21 45502119 N DUP 4
SRR1766471.11294967 chr21 45501850 N chr21 45502023 N DEL 10
SRR1766475.10758435 chr21 45501850 N chr21 45502023 N DEL 10
SRR1766449.1431250 chr21 45501850 N chr21 45502023 N DEL 10
SRR1766465.2663227 chr21 45501849 N chr21 45502109 N DEL 13
SRR1766477.4743806 chr21 45501849 N chr21 45502109 N DEL 15
SRR1766447.3396728 chr21 45502086 N chr21 45502218 N DEL 31
SRR1766448.1960208 chr21 45501914 N chr21 45502218 N DEL 16
SRR1766456.4267116 chr21 45502086 N chr21 45502218 N DEL 30
SRR1766474.2654014 chr21 45502086 N chr21 45502218 N DEL 24
SRR1766454.6352513 chr21 45502086 N chr21 45502218 N DEL 23
SRR1766471.12028313 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766477.4370754 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766461.5320310 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766473.7606447 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766448.840955 chr21 45502108 N chr21 45502239 N DEL 38
SRR1766443.9979007 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766472.8823673 chr21 45502108 N chr21 45502239 N DEL 38
SRR1766452.863021 chr21 45501871 N chr21 45502218 N DEL 21
SRR1766454.7710972 chr21 45502108 N chr21 45502239 N DEL 38
SRR1766474.4879850 chr21 45501871 N chr21 45502218 N DEL 15
SRR1766469.4529495 chr21 45502108 N chr21 45502239 N DEL 22
SRR1766464.4951487 chr21 45502108 N chr21 45502239 N DEL 22
SRR1766448.9862027 chr21 45502108 N chr21 45502239 N DEL 22
SRR1766483.8762190 chr21 45502108 N chr21 45502239 N DEL 22
SRR1766446.10458244 chr21 45501834 N chr21 45502224 N DEL 5
SRR1766483.7124964 chr21 45501834 N chr21 45502224 N DEL 5
SRR1766450.9359300 chr21 45501835 N chr21 45502225 N DEL 5
SRR1766483.10694395 chr21 45501839 N chr21 45502229 N DEL 4
SRR1766442.44674105 chr21 45502108 N chr21 45502239 N DEL 15
SRR1766469.6628223 chr21 45502112 N chr21 45502243 N DEL 11
SRR1766446.4480242 chr21 45502116 N chr21 45502247 N DEL 7
SRR1766470.1702057 chr21 45502117 N chr21 45502248 N DEL 6
SRR1766471.5322620 chr6 34683570 N chr6 34683627 N DUP 1
SRR1766485.7649540 chr6 34683567 N chr6 34683648 N DUP 9
SRR1766470.912384 chr6 34683567 N chr6 34683648 N DUP 11
SRR1766473.688089 chr6 34683567 N chr6 34683648 N DUP 11
SRR1766442.8348651 chr6 34683567 N chr6 34683648 N DUP 13
SRR1766443.3159768 chr10 46490102 N chr10 46490358 N DUP 2
SRR1766454.9560192 chr10 46490196 N chr10 46490340 N DUP 5
SRR1766455.6150538 chr10 46490119 N chr10 46490364 N DUP 5
SRR1766461.2198585 chr3 106074817 N chr3 106075069 N DUP 5
SRR1766468.2770024 chr3 106074815 N chr3 106074942 N DEL 4
SRR1766480.5579308 chr17 68834726 N chr17 68834826 N DEL 9
SRR1766480.2772431 chr18 49003377 N chr18 49003429 N DEL 8
SRR1766450.2828145 chr12 42501 N chr12 42929 N DUP 1
SRR1766474.10865485 chr12 42611 N chr12 42738 N DEL 5
SRR1766451.489135 chr12 42613 N chr12 42740 N DEL 7
SRR1766442.31433185 chr12 42548 N chr12 42724 N DEL 4
SRR1766471.966372 chr12 42511 N chr12 42814 N DEL 1
SRR1766465.9762385 chr15 61098258 N chr15 61098363 N DEL 1
SRR1766442.1034664 chr15 61098202 N chr15 61098358 N DEL 1
SRR1766466.8943973 chr20 35539467 N chr20 35539807 N DUP 5
SRR1766476.9605911 chr20 35539467 N chr20 35539807 N DUP 5
SRR1766476.2167019 chr20 35539469 N chr20 35539815 N DUP 6
SRR1766464.6886620 chr20 35539493 N chr20 35539583 N DUP 5
SRR1766446.4881816 chr20 35539493 N chr20 35539583 N DUP 5
SRR1766446.3713520 chr20 35539552 N chr20 35539680 N DUP 2
SRR1766464.10567720 chr20 35539681 N chr20 35539732 N DEL 12
SRR1766463.9499511 chr20 35539681 N chr20 35539732 N DEL 12
SRR1766455.9831150 chr20 35539681 N chr20 35539732 N DEL 6
SRR1766445.2516648 chr20 35539681 N chr20 35539732 N DEL 9
SRR1766453.6345054 chr20 35539681 N chr20 35539732 N DEL 9
SRR1766470.7981031 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766481.6709691 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766469.8182093 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766477.5894362 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766482.7814309 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766476.9366379 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766468.8036179 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766445.3171783 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766470.155980 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766449.7488778 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766466.11070763 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766472.253939 chr20 35539681 N chr20 35539732 N DEL 5
SRR1766442.42229746 chr20 35539486 N chr20 35539732 N DEL 5
SRR1766449.6875547 chr20 35539486 N chr20 35539732 N DEL 5
SRR1766447.10462480 chr20 35539486 N chr20 35539732 N DEL 5
SRR1766485.9304955 chr20 35539486 N chr20 35539732 N DEL 5
SRR1766478.2690806 chr20 35539486 N chr20 35539732 N DEL 5
SRR1766442.34887087 chr20 35539486 N chr20 35539732 N DEL 5
SRR1766484.929094 chr20 35539461 N chr20 35539732 N DEL 5
SRR1766447.8332153 chr20 35539471 N chr20 35539742 N DEL 5
SRR1766448.4362979 chr20 35539474 N chr20 35539745 N DEL 2
SRR1766454.11029363 chr16 58598156 N chr16 58598290 N DUP 5
SRR1766445.4742696 chr10 41779141 N chr10 41779389 N DEL 5
SRR1766474.11674361 chr10 41779427 N chr10 41779601 N DEL 4
SRR1766471.9899354 chr1 39869761 N chr1 39869841 N DEL 4
SRR1766485.3080118 chr19 621074 N chr19 621137 N DEL 22
SRR1766449.3144827 chr19 621074 N chr19 621137 N DEL 23
SRR1766458.1133797 chr19 621074 N chr19 621137 N DEL 26
SRR1766482.5533032 chr12 132317078 N chr12 132317264 N DEL 1
SRR1766462.9828690 chr12 132317085 N chr12 132317140 N DEL 1
SRR1766461.2564736 chr12 132317140 N chr12 132317242 N DUP 36
SRR1766471.4959538 chr1 162760614 N chr1 162760687 N DEL 7
SRR1766445.6924633 chr1 162760616 N chr1 162760689 N DEL 7
SRR1766444.7132994 chr1 162760617 N chr1 162760690 N DEL 7
SRR1766456.2841284 chr1 162760643 N chr1 162760696 N DEL 6
SRR1766446.2961395 chr1 162760646 N chr1 162760699 N DEL 3
SRR1766457.7681890 chr14 22888991 N chr14 22889147 N DUP 3
SRR1766481.9912671 chr6 1542157 N chr6 1542410 N DEL 7
SRR1766448.9099191 chr6 1542134 N chr6 1542359 N DEL 36
SRR1766442.39847886 chr6 1542137 N chr6 1542455 N DEL 2
SRR1766451.10700839 chr7 126373391 N chr7 126373451 N DEL 7
SRR1766450.3929579 chr7 126373396 N chr7 126373500 N DEL 3
SRR1766442.21438920 chr5 86032860 N chr5 86032911 N DEL 2
SRR1766468.1279516 chr19 42370669 N chr19 42370780 N DEL 1
SRR1766453.7456609 chr1 11522689 N chr1 11522844 N DEL 5
SRR1766481.10819592 chr1 11522679 N chr1 11522801 N DEL 1
SRR1766459.5517392 chr1 11522690 N chr1 11522911 N DEL 11
SRR1766448.4861640 chr1 11522690 N chr1 11522911 N DEL 18
SRR1766456.3063338 chr1 11522690 N chr1 11522911 N DEL 20
SRR1766445.6787493 chr1 11522701 N chr1 11522790 N DEL 18
SRR1766471.4990592 chr1 11522701 N chr1 11522790 N DEL 25
SRR1766462.9815771 chr1 11522701 N chr1 11522834 N DEL 23
SRR1766455.766176 chr1 11522739 N chr1 11522828 N DEL 5
SRR1766459.6434565 chr1 11522701 N chr1 11522790 N DEL 37
SRR1766442.13372194 chr1 11522672 N chr1 11522981 N DEL 20
SRR1766464.906067 chr1 11522745 N chr1 11522834 N DEL 5
SRR1766469.6336979 chr1 11522911 N chr1 11522976 N DUP 15
SRR1766482.3461498 chr1 11522745 N chr1 11522944 N DEL 21
SRR1766460.10284557 chr1 11522777 N chr1 11522866 N DEL 16
SRR1766442.11033935 chr1 11522733 N chr1 11522864 N DUP 9
SRR1766448.2677992 chr1 11522766 N chr1 11523020 N DEL 18
SRR1766468.3122618 chr1 11522771 N chr1 11522836 N DUP 16
SRR1766474.11193977 chr1 11522832 N chr1 11522888 N DEL 6
SRR1766444.3020589 chr1 11522932 N chr1 11522997 N DUP 20
SRR1766476.3342138 chr1 11522723 N chr1 11522779 N DEL 16
SRR1766481.6948997 chr1 11522800 N chr1 11522856 N DEL 15
SRR1766459.11097738 chr1 11522789 N chr1 11522964 N DUP 26
SRR1766474.2416296 chr1 11522778 N chr1 11522865 N DUP 15
SRR1766467.2864822 chr1 11522757 N chr1 11522855 N DUP 14
SRR1766471.12301012 chr1 11522690 N chr1 11522790 N DEL 4
SRR1766442.47184389 chr1 11522705 N chr1 11522761 N DEL 10
SRR1766482.7986008 chr1 11522811 N chr1 11522964 N DUP 13
SRR1766455.766176 chr1 11522855 N chr1 11522999 N DEL 15
SRR1766469.9457784 chr1 11522763 N chr1 11523081 N DUP 9
SRR1766462.1403498 chr1 11522722 N chr1 11522778 N DEL 12
SRR1766460.10284557 chr1 11522856 N chr1 11523020 N DUP 11
SRR1766476.7871370 chr1 11522801 N chr1 11523042 N DUP 5
SRR1766477.3418572 chr1 11522801 N chr1 11522899 N DUP 11
SRR1766447.1021930 chr1 11522847 N chr1 11522901 N DUP 15
SRR1766482.3461498 chr1 11522833 N chr1 11522898 N DUP 15
SRR1766449.10815081 chr1 11522867 N chr1 11522954 N DUP 15
SRR1766474.2416296 chr1 11522724 N chr1 11522877 N DUP 14
SRR1766472.11932065 chr1 11522845 N chr1 11522945 N DEL 5
SRR1766448.8745751 chr1 11522680 N chr1 11522976 N DUP 32
SRR1766444.5884168 chr1 11522844 N chr1 11522911 N DEL 15
SRR1766442.36692428 chr1 11522778 N chr1 11523008 N DUP 20
SRR1766459.11097738 chr1 11522837 N chr1 11522968 N DUP 10
SRR1766481.6698992 chr1 11522690 N chr1 11522909 N DUP 9
SRR1766472.1438968 chr1 11522673 N chr1 11522914 N DUP 20
SRR1766447.10571861 chr1 11522790 N chr1 11522912 N DEL 13
SRR1766477.3418572 chr1 11522834 N chr1 11522965 N DUP 10
SRR1766457.759551 chr1 11522834 N chr1 11522899 N DUP 15
SRR1766465.4579191 chr1 11522790 N chr1 11523064 N DUP 10
SRR1766444.1242946 chr1 11522889 N chr1 11522987 N DUP 10
SRR1766466.1601608 chr1 11522778 N chr1 11522865 N DUP 9
SRR1766458.3373386 chr1 11522779 N chr1 11522921 N DUP 15
SRR1766481.3241932 chr1 11522878 N chr1 11523042 N DUP 25
SRR1766467.2534300 chr1 11522789 N chr1 11522887 N DUP 20
SRR1766475.7604249 chr1 11522722 N chr1 11522833 N DEL 5
SRR1766462.9391873 chr1 11522887 N chr1 11522943 N DEL 17
SRR1766467.2534300 chr1 11522833 N chr1 11522898 N DUP 10
SRR1766447.966989 chr1 11522795 N chr1 11522871 N DUP 19
SRR1766458.598827 chr1 11522759 N chr1 11522958 N DEL 20
SRR1766483.3694014 chr1 11522833 N chr1 11522887 N DUP 6
SRR1766468.1363934 chr1 11522833 N chr1 11522898 N DUP 25
SRR1766457.759551 chr1 11522688 N chr1 11522843 N DEL 6
SRR1766445.2206400 chr1 11522756 N chr1 11522953 N DUP 16
SRR1766447.3775181 chr1 11522833 N chr1 11522898 N DUP 14
SRR1766458.8995500 chr1 11522682 N chr1 11522978 N DUP 11
SRR1766477.8399597 chr1 11522782 N chr1 11522990 N DUP 15
SRR1766446.2022640 chr1 11522690 N chr1 11522845 N DEL 9
SRR1766476.7871370 chr1 11522673 N chr1 11522892 N DUP 20
SRR1766472.2718692 chr1 11522728 N chr1 11522839 N DEL 11
SRR1766482.7986008 chr1 11522833 N chr1 11522920 N DUP 20
SRR1766449.318750 chr1 11522811 N chr1 11522909 N DUP 20
SRR1766450.5199216 chr1 11522833 N chr1 11522964 N DUP 5
SRR1766460.1744327 chr1 11522844 N chr1 11522900 N DEL 20
SRR1766458.598827 chr1 11522834 N chr1 11522910 N DUP 10
SRR1766463.715839 chr1 11522857 N chr1 11522944 N DUP 5
SRR1766482.1406693 chr1 11522733 N chr1 11522864 N DUP 31
SRR1766468.1363934 chr1 11522789 N chr1 11522964 N DUP 20
SRR1766447.966989 chr1 11522789 N chr1 11522898 N DUP 20
SRR1766472.11932065 chr1 11522689 N chr1 11522888 N DEL 10
SRR1766461.2232196 chr1 11522757 N chr1 11522921 N DUP 21
SRR1766457.1623244 chr1 11522933 N chr1 11522987 N DUP 10
SRR1766478.4754 chr1 11522877 N chr1 11522955 N DEL 20
SRR1766447.9072749 chr1 11522878 N chr1 11523009 N DUP 20
SRR1766482.10486760 chr1 11522800 N chr1 11522900 N DEL 10
SRR1766471.7637015 chr1 11522673 N chr1 11522892 N DUP 15
SRR1766484.5106505 chr1 11522899 N chr1 11522999 N DEL 14
SRR1766483.3694014 chr1 11522801 N chr1 11522899 N DUP 20
SRR1766471.2626925 chr1 11522876 N chr1 11522943 N DEL 10
SRR1766464.906067 chr1 11522683 N chr1 11522946 N DUP 16
SRR1766480.4017982 chr1 11522867 N chr1 11522954 N DUP 15
SRR1766484.5106505 chr1 11522713 N chr1 11522822 N DUP 15
SRR1766463.9240650 chr1 11522893 N chr1 11523004 N DEL 10
SRR1766448.2677992 chr1 11522778 N chr1 11523010 N DEL 20
SRR1766460.1744327 chr1 11522746 N chr1 11522833 N DUP 10
SRR1766467.4875381 chr1 11522733 N chr1 11523029 N DUP 11
SRR1766442.32466797 chr1 11522943 N chr1 11523063 N DUP 10
SRR1766449.9867223 chr1 11522723 N chr1 11522977 N DEL 20
SRR1766447.9072749 chr1 11522680 N chr1 11522976 N DUP 26
SRR1766469.1635488 chr1 11522779 N chr1 11523042 N DUP 20
SRR1766469.550113 chr1 11522909 N chr1 11522998 N DEL 12
SRR1766483.8843556 chr1 11522783 N chr1 11523103 N DEL 25
SRR1766477.6118014 chr1 11522768 N chr1 11523053 N DUP 25
SRR1766483.11554571 chr1 11522866 N chr1 11523087 N DEL 10
SRR1766442.36692428 chr1 11522807 N chr1 11523072 N DEL 10
SRR1766477.1710911 chr1 11522866 N chr1 11523087 N DEL 15
SRR1766442.10152581 chr1 11522783 N chr1 11523103 N DEL 20
SRR1766446.6835560 chr1 11522877 N chr1 11523087 N DEL 15
SRR1766470.3235227 chr1 11522717 N chr1 11523103 N DEL 18
SRR1766479.4367259 chr1 11522888 N chr1 11523087 N DEL 17
SRR1766475.2047625 chr1 11522871 N chr1 11523136 N DEL 26
SRR1766442.40938459 chr1 11522717 N chr1 11523103 N DEL 5
SRR1766481.10793214 chr1 11522794 N chr1 11523103 N DEL 6
SRR1766460.1469741 chr1 11522854 N chr1 11523108 N DEL 9
SRR1766478.3144285 chr6 35196095 N chr6 35196209 N DEL 5
SRR1766474.7916384 chr6 35196112 N chr6 35196224 N DUP 5
SRR1766484.6098070 chr8 1912454 N chr8 1912521 N DUP 5
SRR1766444.4167185 chr8 1912360 N chr8 1912495 N DUP 6
SRR1766458.4178085 chr8 1912454 N chr8 1912521 N DUP 5
SRR1766485.5642650 chr8 1912454 N chr8 1912521 N DUP 5
SRR1766462.5583317 chr8 1912454 N chr8 1912521 N DUP 5
SRR1766461.6546037 chr8 1912454 N chr8 1912521 N DUP 5
SRR1766454.5087424 chr8 1912454 N chr8 1912521 N DUP 5
SRR1766455.6227646 chr8 1912533 N chr8 1912600 N DUP 5
SRR1766450.4827719 chr8 1912533 N chr8 1912600 N DUP 5
SRR1766448.3080713 chr8 1912359 N chr8 1912641 N DEL 5
SRR1766444.4167185 chr8 1912377 N chr8 1912659 N DEL 22
SRR1766464.9306979 chr8 1912669 N chr8 1912736 N DUP 5
SRR1766465.3998850 chr10 1377070 N chr10 1377298 N DUP 1
SRR1766465.8277673 chr10 1377136 N chr10 1377297 N DEL 5
SRR1766446.546244 chr10 1377185 N chr10 1377383 N DEL 5
SRR1766458.5797418 chr4 6512034 N chr4 6512659 N DEL 26
SRR1766467.580406 chr4 6512027 N chr4 6512430 N DEL 2
SRR1766462.1512512 chr4 6512078 N chr4 6512181 N DEL 10
SRR1766462.7526382 chr4 6511915 N chr4 6512055 N DUP 25
SRR1766443.5814116 chr4 6511768 N chr4 6512007 N DUP 21
SRR1766473.7629812 chr4 6511991 N chr4 6512443 N DUP 25
SRR1766479.12325215 chr4 6511668 N chr4 6511969 N DEL 4
SRR1766464.1845413 chr4 6512032 N chr4 6512685 N DUP 17
SRR1766462.7118319 chr4 6511969 N chr4 6512046 N DUP 10
SRR1766442.17040874 chr4 6511764 N chr4 6512008 N DEL 1
SRR1766451.4246617 chr4 6511751 N chr4 6512788 N DUP 15
SRR1766442.37250888 chr4 6511696 N chr4 6511964 N DEL 10
SRR1766442.32331045 chr4 6512514 N chr4 6512803 N DEL 17
SRR1766453.7211894 chr4 6512049 N chr4 6512641 N DEL 20
SRR1766442.26404495 chr4 6512051 N chr4 6512712 N DEL 21
SRR1766466.6951659 chr4 6511660 N chr4 6512715 N DUP 2
SRR1766467.6755552 chr4 6511549 N chr4 6511937 N DEL 2
SRR1766464.6617698 chr4 6512005 N chr4 6512174 N DEL 15
SRR1766443.946713 chr4 6511751 N chr4 6512059 N DUP 19
SRR1766480.44355 chr4 6511672 N chr4 6512157 N DUP 15
SRR1766462.1106642 chr4 6511695 N chr4 6511870 N DEL 20
SRR1766463.9707609 chr4 6512061 N chr4 6512587 N DEL 15
SRR1766445.6525602 chr4 6512005 N chr4 6512793 N DUP 6
SRR1766479.4778171 chr4 6511987 N chr4 6512391 N DUP 12
SRR1766462.1998124 chr4 6512040 N chr4 6512404 N DEL 16
SRR1766470.8707988 chr4 6511789 N chr4 6512139 N DUP 9
SRR1766479.9659673 chr4 6512511 N chr4 6512803 N DEL 11
SRR1766482.7953450 chr4 6511565 N chr4 6512146 N DUP 15
SRR1766481.9635619 chr4 6512072 N chr4 6512595 N DEL 10
SRR1766486.4322751 chr4 6512011 N chr4 6512085 N DUP 11
SRR1766459.2358773 chr4 6511803 N chr4 6511909 N DEL 15
SRR1766449.9487334 chr4 6511719 N chr4 6512686 N DEL 15
SRR1766473.7629812 chr4 6512154 N chr4 6512515 N DEL 23
SRR1766443.6249558 chr4 6511900 N chr4 6511967 N DEL 19
SRR1766470.1436507 chr4 6511773 N chr4 6512806 N DEL 24
SRR1766484.11942807 chr4 6511443 N chr4 6512801 N DUP 4
SRR1766465.5187428 chr4 6511714 N chr4 6511863 N DUP 23
SRR1766480.1557525 chr4 6512001 N chr4 6512092 N DEL 10
SRR1766457.5541988 chr4 6511985 N chr4 6512719 N DUP 7
SRR1766449.9019694 chr4 6512042 N chr4 6512166 N DEL 10
SRR1766442.17603216 chr4 6511789 N chr4 6512079 N DUP 26
SRR1766476.884049 chr4 6511783 N chr4 6512681 N DEL 16
SRR1766467.7134931 chr4 6512055 N chr4 6512662 N DEL 9
SRR1766464.7167864 chr4 6512163 N chr4 6512662 N DEL 21
SRR1766474.11273852 chr4 6511751 N chr4 6512038 N DUP 18
SRR1766478.7571584 chr4 6512036 N chr4 6512310 N DEL 15
SRR1766444.2166882 chr4 6511719 N chr4 6512233 N DEL 26
SRR1766479.13279782 chr4 6511684 N chr4 6512076 N DUP 15
SRR1766467.6755552 chr4 6512267 N chr4 6512625 N DEL 16
SRR1766483.9041336 chr4 6511675 N chr4 6511988 N DEL 2
SRR1766461.4800950 chr4 6511540 N chr4 6511679 N DEL 2
SRR1766483.11286513 chr4 6512436 N chr4 6512674 N DEL 17
SRR1766481.8785133 chr4 6511659 N chr4 6512053 N DUP 25
SRR1766455.4043507 chr4 6511719 N chr4 6511840 N DEL 20
SRR1766477.8968558 chr4 6511751 N chr4 6512068 N DUP 19
SRR1766484.3012884 chr4 6511688 N chr4 6512838 N DEL 10
SRR1766474.7706815 chr4 6511699 N chr4 6512073 N DUP 10
SRR1766442.46992958 chr4 6512445 N chr4 6512641 N DEL 18
SRR1766462.5307146 chr4 6512041 N chr4 6512390 N DEL 15
SRR1766483.11530087 chr4 6511670 N chr4 6512817 N DEL 1
SRR1766467.2766808 chr4 6512334 N chr4 6512803 N DEL 17
SRR1766471.729973 chr4 6511727 N chr4 6512022 N DUP 11
SRR1766442.36245973 chr4 6511452 N chr4 6512809 N DEL 9
SRR1766472.643150 chr4 6512238 N chr4 6512803 N DEL 17
SRR1766460.3690639 chr4 6511522 N chr4 6511655 N DEL 12
SRR1766472.2957428 chr4 6512014 N chr4 6512805 N DUP 7
SRR1766463.7471291 chr4 6512034 N chr4 6512803 N DEL 30
SRR1766480.1267692 chr4 6512054 N chr4 6512298 N DEL 7
SRR1766474.10163277 chr4 6511660 N chr4 6512025 N DUP 5
SRR1766454.1081355 chr4 6511859 N chr4 6512074 N DUP 20
SRR1766481.5943877 chr4 6512014 N chr4 6512670 N DUP 12
SRR1766479.5221559 chr4 6511719 N chr4 6512728 N DEL 20
SRR1766442.21849030 chr4 6511794 N chr4 6512069 N DUP 21
SRR1766462.9182089 chr4 6512103 N chr4 6512833 N DEL 4
SRR1766454.4584699 chr4 6511774 N chr4 6512067 N DUP 18
SRR1766442.18117396 chr4 6511963 N chr4 6512553 N DUP 17
SRR1766476.7413809 chr4 6511689 N chr4 6512509 N DEL 20
SRR1766467.924225 chr4 6511666 N chr4 6511971 N DUP 20
SRR1766474.3663873 chr4 6511977 N chr4 6512075 N DUP 17
SRR1766485.7028537 chr4 6511904 N chr4 6512107 N DUP 1
SRR1766484.1532911 chr4 6512238 N chr4 6512803 N DEL 17
SRR1766452.6525913 chr4 6512122 N chr4 6512642 N DEL 17
SRR1766458.6656436 chr4 6512064 N chr4 6512662 N DEL 15
SRR1766469.10460161 chr4 6512008 N chr4 6512079 N DUP 10
SRR1766448.3200470 chr4 6511719 N chr4 6512116 N DEL 5
SRR1766442.15562102 chr4 6511800 N chr4 6512159 N DUP 14
SRR1766444.1067630 chr4 6511948 N chr4 6512442 N DUP 20
SRR1766473.9112661 chr4 6511751 N chr4 6512551 N DUP 21
SRR1766483.11340352 chr4 6512511 N chr4 6512803 N DEL 11
SRR1766476.8828890 chr4 6511972 N chr4 6512421 N DUP 7
SRR1766478.5148229 chr4 6512029 N chr4 6512115 N DUP 17
SRR1766450.7007537 chr4 6511789 N chr4 6512015 N DEL 5
SRR1766446.10068454 chr4 6511672 N chr4 6512064 N DUP 15
SRR1766447.6177714 chr4 6512603 N chr4 6512832 N DEL 26
SRR1766449.10862705 chr4 6511522 N chr4 6511691 N DEL 10
SRR1766454.1580500 chr4 6512244 N chr4 6512812 N DEL 6
SRR1766483.9989377 chr4 6511719 N chr4 6512311 N DEL 23
SRR1766442.22326896 chr4 6511933 N chr4 6511983 N DUP 11
SRR1766466.4087488 chr4 6511541 N chr4 6512235 N DEL 16
SRR1766471.3979794 chr4 6512051 N chr4 6512682 N DEL 25
SRR1766458.6656436 chr4 6511459 N chr4 6511844 N DEL 5
SRR1766472.6267779 chr4 6512004 N chr4 6512326 N DEL 12
SRR1766479.4778171 chr4 6511670 N chr4 6512811 N DEL 7
SRR1766473.6780587 chr4 6511981 N chr4 6512658 N DUP 5
SRR1766444.2734046 chr4 6511722 N chr4 6512662 N DEL 10
SRR1766476.7290640 chr4 6512078 N chr4 6512628 N DEL 10
SRR1766474.3016922 chr4 6511761 N chr4 6512075 N DUP 11
SRR1766452.5242026 chr4 6512511 N chr4 6512803 N DEL 11
SRR1766442.22389402 chr4 6511751 N chr4 6512062 N DUP 20
SRR1766480.1267692 chr4 6512040 N chr4 6512695 N DEL 20
SRR1766454.1913741 chr4 6511756 N chr4 6512076 N DUP 18
SRR1766442.6046883 chr4 6512010 N chr4 6512695 N DEL 33
SRR1766467.3829509 chr4 6511718 N chr4 6512238 N DEL 25
SRR1766476.5210159 chr4 6511987 N chr4 6512040 N DUP 20
SRR1766452.6525913 chr4 6512054 N chr4 6512475 N DEL 15
SRR1766443.8001581 chr4 6511966 N chr4 6512030 N DEL 2
SRR1766486.11962074 chr11 134738846 N chr11 134739165 N DEL 4
SRR1766486.8968326 chr11 134738854 N chr11 134739079 N DEL 9
SRR1766460.6596792 chr11 134738821 N chr11 134738982 N DEL 5
SRR1766442.25782208 chr11 134738880 N chr11 134739013 N DEL 19
SRR1766464.1447890 chr11 134738880 N chr11 134739013 N DEL 24
SRR1766442.44233628 chr11 134738880 N chr11 134739013 N DEL 14
SRR1766466.97568 chr11 134738880 N chr11 134739013 N DEL 24
SRR1766472.7390616 chr11 134738880 N chr11 134739013 N DEL 24
SRR1766460.1648769 chr11 134738880 N chr11 134739013 N DEL 24
SRR1766455.618696 chr11 134738883 N chr11 134739042 N DUP 5
SRR1766467.10867589 chr11 134738883 N chr11 134739042 N DUP 5
SRR1766481.8157875 chr11 134738883 N chr11 134739106 N DUP 10
SRR1766461.9897859 chr11 134738891 N chr11 134739050 N DUP 5
SRR1766481.9584675 chr11 134738883 N chr11 134739042 N DUP 5
SRR1766484.9684471 chr11 134738928 N chr11 134738991 N DUP 5
SRR1766443.4839167 chr11 134738883 N chr11 134739042 N DUP 5
SRR1766484.8876146 chr11 134738891 N chr11 134739050 N DUP 8
SRR1766475.10531837 chr11 134738864 N chr11 134738961 N DEL 5
SRR1766460.1937249 chr11 134738950 N chr11 134739045 N DUP 5
SRR1766478.3014565 chr11 134738869 N chr11 134739062 N DEL 3
SRR1766455.7001159 chr11 134738847 N chr11 134739040 N DEL 5
SRR1766486.875628 chr11 134738867 N chr11 134739060 N DEL 15
SRR1766443.2758932 chr11 134738982 N chr11 134739079 N DEL 5
SRR1766475.1287883 chr11 134738982 N chr11 134739079 N DEL 5
SRR1766482.11377240 chr11 134738918 N chr11 134739079 N DEL 5
SRR1766474.3194954 chr11 134738974 N chr11 134739103 N DEL 4
SRR1766478.4865254 chr11 134738858 N chr11 134739115 N DEL 5
SRR1766452.1673892 chr11 134738864 N chr11 134739121 N DEL 2
SRR1766469.265821 chr11 134738835 N chr11 134739186 N DEL 1
SRR1766477.4881521 chr20 24730148 N chr20 24730206 N DUP 5
SRR1766449.8696161 chr20 24730209 N chr20 24730393 N DUP 5
SRR1766484.4750501 chr20 24730213 N chr20 24730338 N DUP 5
SRR1766442.16093572 chr20 24730131 N chr20 24730305 N DEL 2
SRR1766455.7065965 chr18 76896197 N chr18 76896365 N DEL 3
SRR1766466.9068340 chr18 76896348 N chr18 76896411 N DEL 1
SRR1766478.10230582 chr18 76896488 N chr18 76896537 N DUP 10
SRR1766442.18384499 chr18 76896107 N chr18 76896442 N DEL 2
SRR1766469.8108530 chr18 76896486 N chr18 76896672 N DUP 5
SRR1766484.10596280 chr20 56761545 N chr20 56761745 N DUP 4
SRR1766449.4017162 chr20 56761743 N chr20 56761876 N DEL 5
SRR1766484.5506905 chr20 56761639 N chr20 56761979 N DEL 5
SRR1766451.9729379 chr4 2856748 N chr4 2857073 N DEL 10
SRR1766478.2437952 chr4 2856812 N chr4 2857134 N DEL 12
SRR1766479.4303626 chr4 2856796 N chr4 2857118 N DEL 10
SRR1766450.10254967 chr1 45782324 N chr1 45782638 N DEL 2
SRR1766445.10420309 chrX 142126002 N chrX 142126061 N DUP 8
SRR1766442.11037812 chrX 142126082 N chrX 142126142 N DEL 4
SRR1766467.4065500 chrX 142126033 N chrX 142126097 N DEL 10
SRR1766469.5630912 chrX 142126115 N chrX 142126198 N DEL 12
SRR1766459.7612526 chrX 142126115 N chrX 142126198 N DEL 12
SRR1766475.8832170 chrX 142126133 N chrX 142126203 N DEL 4
SRR1766451.2760684 chrX 142126133 N chrX 142126203 N DEL 9
SRR1766479.13050065 chrX 142126133 N chrX 142126203 N DEL 9
SRR1766476.6471060 chrX 142126133 N chrX 142126203 N DEL 11
SRR1766463.5107930 chrX 142126133 N chrX 142126203 N DEL 14
SRR1766485.412779 chrX 142126133 N chrX 142126203 N DEL 23
SRR1766452.7510255 chrX 142126133 N chrX 142126203 N DEL 15
SRR1766482.4570856 chrX 142126145 N chrX 142126215 N DEL 1
SRR1766479.3154712 chr21 42591832 N chr21 42591903 N DEL 5
SRR1766471.2454953 chr21 42591832 N chr21 42591903 N DEL 10
SRR1766452.8095714 chr21 42591742 N chr21 42591931 N DEL 1
SRR1766469.9196717 chr21 42591869 N chr21 42591926 N DEL 6
SRR1766451.3282733 chr21 42591870 N chr21 42591949 N DEL 5
SRR1766460.8628722 chr8 57382792 N chr8 57382852 N DUP 6
SRR1766476.7281332 chr8 57382456 N chr8 57382895 N DEL 6
SRR1766446.4597257 chr8 57382459 N chr8 57382898 N DEL 3
SRR1766456.6140935 chr14 67193288 N chr14 67193341 N DEL 2
SRR1766442.15357695 chr14 67193288 N chr14 67193341 N DEL 4
SRR1766448.5628682 chr14 67193288 N chr14 67193341 N DEL 4
SRR1766466.11219754 chr14 67193291 N chr14 67193344 N DEL 9
SRR1766466.2206216 chr14 67193293 N chr14 67193346 N DEL 9
SRR1766446.3689052 chr10 122470729 N chr10 122470806 N DEL 5
SRR1766466.4308920 chr10 122470656 N chr10 122470731 N DUP 5
SRR1766483.4071832 chr10 122470656 N chr10 122470731 N DUP 5
SRR1766483.359313 chr10 122470656 N chr10 122470731 N DUP 5
SRR1766473.1352488 chr10 122470656 N chr10 122470731 N DUP 5
SRR1766469.2226416 chr10 122470656 N chr10 122470731 N DUP 5
SRR1766477.5526182 chr10 122470672 N chr10 122470749 N DEL 5
SRR1766444.296411 chr10 122470676 N chr10 122470753 N DEL 2
SRR1766475.10750330 chr14 90528757 N chr14 90528893 N DUP 5
SRR1766462.5943113 chr14 90528799 N chr14 90529096 N DUP 5
SRR1766452.5480858 chr14 90528799 N chr14 90529096 N DUP 5
SRR1766472.9284792 chr14 90528799 N chr14 90529096 N DUP 5
SRR1766442.8181176 chr14 90528807 N chr14 90529104 N DUP 5
SRR1766444.2581949 chr14 90528807 N chr14 90529104 N DUP 5
SRR1766445.8953653 chr14 90528717 N chr14 90528892 N DEL 1
SRR1766454.10706367 chr14 90528771 N chr14 90529068 N DUP 5
SRR1766458.4935064 chr14 90528818 N chr14 90528993 N DEL 5
SRR1766458.7434075 chr14 90528837 N chr14 90529097 N DUP 7
SRR1766474.8045795 chr18 41349885 N chr18 41349953 N DUP 4
SRR1766449.330591 chr18 41349899 N chr18 41349967 N DUP 13
SRR1766442.22059425 chr18 41349926 N chr18 41350003 N DUP 22
SRR1766485.9523507 chr18 41349926 N chr18 41350003 N DUP 22
SRR1766480.2338625 chr18 41349886 N chr18 41349996 N DUP 8
SRR1766484.11242492 chr18 41349885 N chr18 41349953 N DUP 24
SRR1766463.9726641 chr18 41349886 N chr18 41349996 N DUP 9
SRR1766451.4955734 chr18 41349886 N chr18 41349996 N DUP 12
SRR1766448.8984370 chr18 41349886 N chr18 41349996 N DUP 13
SRR1766451.6414193 chr18 41349886 N chr18 41349996 N DUP 14
SRR1766460.3994208 chr18 41349886 N chr18 41349996 N DUP 16
SRR1766485.4573420 chr18 41349886 N chr18 41349996 N DUP 16
SRR1766482.3731191 chr18 41349926 N chr18 41350003 N DUP 21
SRR1766450.1825494 chr18 41349886 N chr18 41349996 N DUP 28
SRR1766467.5983629 chr18 41349886 N chr18 41349996 N DUP 28
SRR1766453.2523118 chr18 41349926 N chr18 41350003 N DUP 18
SRR1766454.6080382 chr18 41349893 N chr18 41349961 N DUP 7
SRR1766442.7309810 chr18 41349926 N chr18 41350003 N DUP 20
SRR1766460.5261827 chr18 41349899 N chr18 41349967 N DUP 1
SRR1766446.2070074 chr18 41349926 N chr18 41350003 N DUP 29
SRR1766442.1331155 chr18 41349926 N chr18 41350003 N DUP 30
SRR1766470.9433185 chr18 41349926 N chr18 41350003 N DUP 32
SRR1766471.8057925 chr5 173128934 N chr5 173129271 N DEL 30
SRR1766454.3227865 chr5 173129051 N chr5 173129388 N DEL 5
SRR1766445.9769098 chr5 173129150 N chr5 173129487 N DEL 5
SRR1766485.12036142 chr5 173129190 N chr5 173129527 N DEL 10
SRR1766442.40572898 chr5 173129047 N chr5 173129384 N DEL 1
SRR1766452.3217424 chr5 173129124 N chr5 173129461 N DEL 5
SRR1766461.10990412 chr5 173129209 N chr5 173129546 N DEL 20
SRR1766445.895049 chr9 40590175 N chr9 40590342 N DEL 13
SRR1766475.9732305 chr6 94711526 N chr6 94711888 N DUP 14
SRR1766442.30049145 chr6 94711526 N chr6 94711888 N DUP 14
SRR1766442.26998185 chr6 94711670 N chr6 94711854 N DUP 10
SRR1766454.8228689 chr6 94711525 N chr6 94711761 N DEL 11
SRR1766475.9732305 chr6 94711511 N chr6 94711888 N DUP 14
SRR1766449.6667992 chr3 163618630 N chr3 163618735 N DEL 7
SRR1766466.9728593 chr5 162906168 N chr5 162906219 N DEL 14
SRR1766457.772081 chr5 162906168 N chr5 162906219 N DEL 42
SRR1766447.6415499 chr13 63111392 N chr13 63111465 N DUP 5
SRR1766472.140325 chr10 73262122 N chr10 73262217 N DUP 12
SRR1766478.1726151 chr10 73262122 N chr10 73262217 N DUP 12
SRR1766484.9450932 chr10 73262122 N chr10 73262217 N DUP 12
SRR1766449.984472 chr10 73262172 N chr10 73262231 N DEL 10
SRR1766454.10509117 chr10 73262145 N chr10 73262240 N DEL 1
SRR1766473.11785463 chr9 69340761 N chr9 69340856 N DEL 4
SRR1766470.723184 chr9 69340774 N chr9 69340841 N DEL 10
SRR1766473.7764161 chr9 69340761 N chr9 69340856 N DEL 12
SRR1766474.3914949 chr9 69340785 N chr9 69340946 N DEL 5
SRR1766485.6642500 chr9 69340794 N chr9 69340951 N DEL 7
SRR1766475.2695665 chr9 69340785 N chr9 69340934 N DEL 10
SRR1766486.7830327 chr9 69340745 N chr9 69340824 N DUP 9
SRR1766477.4935965 chr9 69340830 N chr9 69340951 N DEL 11
SRR1766480.8708878 chr9 69340818 N chr9 69340885 N DEL 16
SRR1766453.10133426 chr9 69340816 N chr9 69340939 N DUP 24
SRR1766484.5103234 chr9 69340817 N chr9 69340886 N DUP 10
SRR1766460.3848292 chr9 69340870 N chr9 69340939 N DEL 23
SRR1766442.36868283 chr9 69340892 N chr9 69340977 N DUP 5
SRR1766467.324415 chr9 69340843 N chr9 69340950 N DEL 38
SRR1766445.6515273 chr9 69340897 N chr9 69340976 N DUP 10
SRR1766458.7064041 chr9 69340860 N chr9 69340913 N DEL 17
SRR1766476.10601518 chr9 69340928 N chr9 69340977 N DUP 5
SRR1766476.10594913 chr9 69340870 N chr9 69340939 N DEL 19
SRR1766482.2451125 chr9 69340870 N chr9 69340939 N DEL 15
SRR1766442.32359574 chr9 69340870 N chr9 69340939 N DEL 9
SRR1766484.1704866 chr9 69340870 N chr9 69340939 N DEL 9
SRR1766463.10093242 chr9 69340767 N chr9 69340942 N DEL 9
SRR1766476.8840086 chr9 69340844 N chr9 69340965 N DEL 7
SRR1766463.9860548 chr9 69340774 N chr9 69340965 N DEL 12
SRR1766449.636547 chr9 69340850 N chr9 69340971 N DEL 7
SRR1766459.3000442 chr9 69340853 N chr9 69340974 N DEL 6
SRR1766447.3101985 chr4 157544042 N chr4 157544095 N DEL 57
SRR1766485.6648189 chr3 73738838 N chr3 73738953 N DEL 5
SRR1766454.8628093 chr18 72675618 N chr18 72675709 N DEL 3
SRR1766449.3755098 chr18 72675618 N chr18 72675709 N DEL 5
SRR1766459.11320707 chr18 72675642 N chr18 72675778 N DEL 5
SRR1766469.3552383 chr18 72675642 N chr18 72675778 N DEL 5
SRR1766472.3524687 chr18 72675722 N chr18 72675858 N DEL 5
SRR1766449.70100 chr18 72675722 N chr18 72675858 N DEL 5
SRR1766482.3985323 chr18 72675722 N chr18 72675858 N DEL 5
SRR1766442.8114676 chr18 72675635 N chr18 72675724 N DUP 5
SRR1766484.8751317 chr18 72675635 N chr18 72675724 N DUP 5
SRR1766474.7739364 chr18 72675641 N chr18 72675730 N DUP 5
SRR1766471.4633476 chr18 72675687 N chr18 72675778 N DEL 15
SRR1766481.11282398 chr18 72675797 N chr18 72675888 N DEL 10
SRR1766479.3512450 chr18 72675708 N chr18 72675797 N DUP 8
SRR1766468.6753293 chr18 72675619 N chr18 72675843 N DUP 1
SRR1766480.3650182 chr18 72675663 N chr18 72675754 N DEL 3
SRR1766479.2750750 chr18 72675816 N chr18 72675907 N DEL 15
SRR1766479.3512450 chr18 72675811 N chr18 72675902 N DEL 10
SRR1766446.1541378 chr18 72675737 N chr18 72675918 N DEL 4
SRR1766484.8751317 chr18 72675767 N chr18 72675948 N DEL 5
SRR1766465.3572067 chr18 72675633 N chr18 72675949 N DEL 5
SRR1766452.1874782 chrX 131135822 N chrX 131135930 N DUP 2
SRR1766455.3019197 chr5 1081135 N chr5 1081216 N DUP 7
SRR1766456.102739 chr5 1081135 N chr5 1081216 N DUP 7
SRR1766478.3639108 chr5 1081135 N chr5 1081214 N DUP 5
SRR1766481.11205265 chr5 1081135 N chr5 1081216 N DUP 7
SRR1766451.3483997 chr2 168631704 N chr2 168631765 N DUP 10
SRR1766457.4946375 chr2 168631704 N chr2 168631765 N DUP 11
SRR1766451.720893 chr21 20587258 N chr21 20587370 N DEL 5
SRR1766463.1316277 chr21 20587256 N chr21 20587370 N DEL 5
SRR1766474.3916281 chr21 20587256 N chr21 20587370 N DEL 5
SRR1766473.3526707 chr21 20587300 N chr21 20587434 N DEL 5
SRR1766442.25455395 chr21 20587300 N chr21 20587434 N DEL 5
SRR1766473.5150155 chr9 10323351 N chr9 10323437 N DEL 8
SRR1766446.9720002 chr17 28810524 N chr17 28810613 N DEL 5
SRR1766468.406534 chr22 16387036 N chr22 16387186 N DUP 5
SRR1766456.4861695 chr3 122747602 N chr3 122747700 N DEL 9
SRR1766473.5390991 chr3 122747620 N chr3 122747716 N DUP 5
SRR1766469.7731842 chr3 122747698 N chr3 122747872 N DUP 5
SRR1766486.4559536 chr3 122747698 N chr3 122747872 N DUP 5
SRR1766478.1554901 chr3 122747769 N chr3 122747895 N DUP 5
SRR1766463.5216538 chr3 122747685 N chr3 122747908 N DUP 5
SRR1766447.7001743 chr3 122747769 N chr3 122747895 N DUP 5
SRR1766468.4852233 chr3 122747685 N chr3 122747908 N DUP 5
SRR1766472.6674727 chr21 40498777 N chr21 40498881 N DEL 5
SRR1766444.7206059 chr21 40498801 N chr21 40498908 N DEL 5
SRR1766482.6869986 chr21 40498824 N chr21 40498885 N DEL 1
SRR1766463.7757231 chr21 40498824 N chr21 40498885 N DEL 2
SRR1766460.4694396 chr21 40498824 N chr21 40498885 N DEL 3
SRR1766444.4806079 chr21 40498824 N chr21 40498885 N DEL 4
SRR1766473.2361610 chr21 40498824 N chr21 40498885 N DEL 4
SRR1766473.6866406 chr21 40498824 N chr21 40498885 N DEL 4
SRR1766458.4550563 chr21 40498824 N chr21 40498885 N DEL 5
SRR1766462.2182359 chr21 40498824 N chr21 40498885 N DEL 7
SRR1766454.8056275 chr21 40498824 N chr21 40498885 N DEL 8
SRR1766461.5970728 chr21 40498824 N chr21 40498885 N DEL 11
SRR1766448.702158 chr21 40498824 N chr21 40498885 N DEL 9
SRR1766469.10376467 chr21 40498826 N chr21 40498885 N DEL 4
SRR1766471.11049906 chr21 40498824 N chr21 40498885 N DEL 7
SRR1766484.6832801 chr21 40498824 N chr21 40498885 N DEL 17
SRR1766479.10786416 chr21 40498741 N chr21 40498791 N DUP 9
SRR1766480.589887 chr21 40498824 N chr21 40498885 N DEL 13
SRR1766459.7914985 chr21 40498824 N chr21 40498885 N DEL 13
SRR1766471.9171108 chr21 40498824 N chr21 40498885 N DEL 16
SRR1766452.9452455 chr21 40498824 N chr21 40498885 N DEL 16
SRR1766442.6581226 chr21 40498864 N chr21 40498955 N DEL 6
SRR1766460.8572665 chr21 40498864 N chr21 40498955 N DEL 10
SRR1766451.8221494 chr21 40498828 N chr21 40498889 N DEL 11
SRR1766454.8056275 chr21 40498795 N chr21 40498895 N DEL 5
SRR1766462.3425978 chr21 40498864 N chr21 40498955 N DEL 15
SRR1766475.609192 chr21 40498792 N chr21 40498966 N DEL 2
SRR1766446.6537908 chr21 40498793 N chr21 40498967 N DEL 1
SRR1766448.6504242 chr21 40498873 N chr21 40498962 N DEL 6
SRR1766450.9251218 chr21 40498870 N chr21 40498959 N DEL 9
SRR1766476.8874557 chr21 40498875 N chr21 40498964 N DEL 4
SRR1766458.9182075 chr21 40498793 N chr21 40498969 N DEL 1
SRR1766460.3089862 chr21 40498869 N chr21 40498960 N DEL 10
SRR1766476.4488547 chr21 40498873 N chr21 40498964 N DEL 6
SRR1766447.1562684 chr12 121750661 N chr12 121751045 N DEL 11
SRR1766469.2479386 chr12 121750803 N chr12 121751030 N DEL 12
SRR1766477.5187207 chr12 121750823 N chr12 121751156 N DEL 5
SRR1766452.801941 chr12 121750646 N chr12 121750990 N DUP 9
SRR1766466.7603159 chr12 121751018 N chr12 121751116 N DEL 1
SRR1766463.6787856 chr12 121751023 N chr12 121751493 N DEL 11
SRR1766447.10334534 chr12 121751029 N chr12 121751474 N DEL 1
SRR1766448.6665453 chr12 121751019 N chr12 121751507 N DUP 5
SRR1766468.1780920 chr12 121750947 N chr12 121751177 N DEL 12
SRR1766467.8598657 chr12 121750655 N chr12 121751247 N DEL 5
SRR1766480.7317745 chr12 121751272 N chr12 121751513 N DUP 11
SRR1766462.9683539 chr12 121750655 N chr12 121751279 N DEL 5
SRR1766459.7797481 chr8 46062699 N chr8 46062872 N DEL 5
SRR1766476.9853407 chr17 8829586 N chr17 8829693 N DUP 9
SRR1766448.1816541 chr17 8829691 N chr17 8829742 N DUP 17
SRR1766474.9694965 chr17 8829560 N chr17 8829703 N DEL 5
SRR1766471.5853055 chr17 8829514 N chr17 8829751 N DEL 15
SRR1766478.3000287 chr16 34599865 N chr16 34600107 N DUP 5
SRR1766471.4697917 chr11 89112662 N chr11 89112823 N DEL 11
SRR1766460.3574579 chr17 22722933 N chr17 22723103 N DUP 5
SRR1766471.1186612 chr17 22722303 N chr17 22723117 N DUP 5
SRR1766450.9221364 chr5 180707399 N chr5 180707706 N DEL 5
SRR1766473.2225107 chr1 144542193 N chr1 144542336 N DEL 6
SRR1766479.7530684 chr6 168257712 N chr6 168257801 N DEL 10
SRR1766445.5859122 chr6 168257676 N chr6 168257745 N DEL 13
SRR1766444.1677376 chr6 168257476 N chr6 168257672 N DEL 7
SRR1766478.7114344 chr6 168257644 N chr6 168257705 N DEL 3
SRR1766442.5103920 chr6 168257746 N chr6 168257795 N DUP 4
SRR1766472.751564 chr6 168257765 N chr6 168257814 N DUP 5
SRR1766442.796572 chr20 64017353 N chr20 64017530 N DEL 5
SRR1766460.172122 chr20 64017433 N chr20 64017564 N DUP 5
SRR1766485.2355786 chr20 64017383 N chr20 64017602 N DUP 5
SRR1766449.2217343 chr20 64017515 N chr20 64017602 N DUP 5
SRR1766478.5479094 chr20 64017515 N chr20 64017602 N DUP 5
SRR1766442.39577855 chr20 64017515 N chr20 64017602 N DUP 5
SRR1766481.10455399 chr20 64017515 N chr20 64017602 N DUP 5
SRR1766476.11182595 chr20 64017515 N chr20 64017602 N DUP 5
SRR1766468.5107672 chr20 64017531 N chr20 64017706 N DUP 5
SRR1766462.1887528 chr20 64017573 N chr20 64017706 N DEL 5
SRR1766448.5931310 chr20 64017397 N chr20 64017750 N DEL 5
SRR1766462.3731772 chr20 64017391 N chr20 64017788 N DEL 16
SRR1766444.2643093 chr20 64017416 N chr20 64017769 N DEL 11
SRR1766458.2376493 chr20 41556394 N chr20 41556459 N DUP 5
SRR1766451.7814960 chr20 41556394 N chr20 41556459 N DUP 6
SRR1766446.5347632 chr22 49476931 N chr22 49477066 N DEL 7
SRR1766465.2597196 chr22 49476992 N chr22 49477381 N DEL 5
SRR1766452.9215856 chr22 49477096 N chr22 49477261 N DEL 6
SRR1766465.3457480 chr22 49477091 N chr22 49477256 N DEL 10
SRR1766458.769346 chr22 49477127 N chr22 49477243 N DEL 5
SRR1766464.10713482 chr22 49476903 N chr22 49477018 N DEL 8
SRR1766481.10478203 chr22 49477091 N chr22 49477948 N DEL 15
SRR1766481.1653144 chr22 49477151 N chr22 49477576 N DEL 4
SRR1766462.10591002 chr22 49476997 N chr22 49477289 N DUP 5
SRR1766467.8368136 chr22 49477282 N chr22 49477895 N DEL 3
SRR1766442.18966119 chr22 49477331 N chr22 49477814 N DEL 2
SRR1766471.11555581 chr22 49477267 N chr22 49477376 N DUP 9
SRR1766467.7030489 chr22 49477091 N chr22 49477313 N DEL 12
SRR1766454.7558473 chr22 49477333 N chr22 49478005 N DUP 6
SRR1766452.131257 chr22 49477031 N chr22 49477417 N DUP 2
SRR1766465.3457480 chr22 49477012 N chr22 49477325 N DEL 11
SRR1766448.10595125 chr22 49477081 N chr22 49477333 N DEL 10
SRR1766442.10179735 chr22 49477534 N chr22 49477671 N DEL 5
SRR1766485.5525528 chr22 49477528 N chr22 49477623 N DEL 10
SRR1766481.2790040 chr22 49477587 N chr22 49477645 N DEL 5
SRR1766468.3263652 chr22 49476991 N chr22 49477599 N DUP 5
SRR1766467.2267873 chr22 49477610 N chr22 49477766 N DEL 14
SRR1766467.9754977 chr22 49477364 N chr22 49477508 N DEL 8
SRR1766461.8752569 chr22 49477347 N chr22 49477616 N DUP 4
SRR1766451.1196526 chr22 49477600 N chr22 49477958 N DEL 5
SRR1766466.5081350 chr22 49476992 N chr22 49477661 N DUP 14
SRR1766465.10122247 chr22 49476922 N chr22 49477571 N DEL 4
SRR1766462.11123785 chr22 49477070 N chr22 49477868 N DUP 10
SRR1766457.3349760 chr22 49477354 N chr22 49477892 N DUP 10
SRR1766477.3135440 chr22 49477052 N chr22 49477906 N DUP 3
SRR1766446.6093525 chr22 49477080 N chr22 49477940 N DEL 5
SRR1766467.8418238 chr22 49477006 N chr22 49477954 N DEL 1
SRR1766481.12591158 chr22 49477502 N chr22 49477953 N DEL 11
SRR1766469.1434362 chr22 49477362 N chr22 49477967 N DEL 5
SRR1766465.2272352 chr22 49477598 N chr22 49477971 N DEL 9
SRR1766467.6876468 chr22 49477092 N chr22 49477979 N DEL 11
SRR1766472.6834379 chr22 49477094 N chr22 49477985 N DEL 1
SRR1766469.3603474 chr22 49477661 N chr22 49477989 N DEL 1
SRR1766447.3220964 chr22 49477908 N chr22 49478019 N DEL 7
SRR1766458.267417 chr22 49477661 N chr22 49478019 N DEL 5
SRR1766450.10933809 chr22 49477661 N chr22 49478019 N DEL 5
SRR1766453.8621767 chr22 49477377 N chr22 49478024 N DEL 5
SRR1766468.4118076 chr10 97193373 N chr10 97193440 N DUP 5
SRR1766460.8446611 chr18 9887642 N chr18 9887823 N DEL 17
SRR1766442.21531532 chr18 9887525 N chr18 9887749 N DUP 14
SRR1766479.13488027 chr18 9887721 N chr18 9887857 N DEL 5
SRR1766442.11268621 chr18 9887555 N chr18 9887646 N DEL 5
SRR1766466.3085849 chr18 9887555 N chr18 9887646 N DEL 5
SRR1766444.1091324 chr18 9887766 N chr18 9887857 N DEL 5
SRR1766456.3273218 chr18 9887604 N chr18 9887695 N DEL 10
SRR1766449.2121950 chr18 9887604 N chr18 9887695 N DEL 5
SRR1766442.30092733 chr18 9887604 N chr18 9887695 N DEL 5
SRR1766477.6360351 chr18 9887565 N chr18 9887701 N DEL 5
SRR1766470.11000406 chr18 9887569 N chr18 9887705 N DEL 5
SRR1766458.9550686 chr18 9887615 N chr18 9887751 N DEL 5
SRR1766459.1308588 chr18 9887585 N chr18 9887766 N DEL 5
SRR1766468.3608113 chr20 4089507 N chr20 4089663 N DEL 5
SRR1766473.575046 chr20 4089507 N chr20 4089663 N DEL 5
SRR1766479.13247960 chr20 4089507 N chr20 4089663 N DEL 5
SRR1766484.1826323 chr20 4089507 N chr20 4089663 N DEL 5
SRR1766453.3606973 chr20 4089507 N chr20 4089663 N DEL 5
SRR1766459.383987 chr7 73137945 N chr7 73138034 N DEL 4
SRR1766448.8387519 chr6 157283053 N chr6 157283466 N DUP 10
SRR1766463.1957723 chr6 157283353 N chr6 157283467 N DUP 5
SRR1766484.7663916 chr6 157283077 N chr6 157283354 N DEL 5
SRR1766485.2498221 chr6 157283078 N chr6 157283401 N DEL 5
SRR1766442.7102652 chr6 157283076 N chr6 157283445 N DEL 5
SRR1766468.1556016 chr6 157283078 N chr6 157283447 N DEL 5
SRR1766469.9135501 chr6 157283063 N chr6 157283455 N DEL 1
SRR1766462.6662113 chr10 67727924 N chr10 67728021 N DUP 5
SRR1766464.5530242 chr10 67727926 N chr10 67728056 N DUP 5
SRR1766450.3033374 chr4 46273632 N chr4 46273689 N DEL 7
SRR1766486.6267016 chr10 123572702 N chr10 123572872 N DEL 3
SRR1766446.2256505 chr1 3834406 N chr1 3834566 N DEL 7
SRR1766455.2723821 chr1 228631236 N chr1 228631289 N DUP 3
SRR1766475.4072308 chr1 228631236 N chr1 228631289 N DUP 4
SRR1766486.1596459 chr1 228631234 N chr1 228631293 N DUP 12
SRR1766478.9047626 chr1 228631236 N chr1 228631289 N DUP 7
SRR1766444.4096235 chr2 118305297 N chr2 118305361 N DEL 12
SRR1766484.11681189 chr2 118305360 N chr2 118305519 N DEL 2
SRR1766465.5107044 chr2 118305257 N chr2 118305316 N DUP 4
SRR1766465.11120104 chr2 118305296 N chr2 118305358 N DUP 10
SRR1766458.7036061 chr2 118305264 N chr2 118305323 N DUP 4
SRR1766442.11735860 chr2 118305297 N chr2 118305361 N DEL 22
SRR1766461.5992344 chr2 118305297 N chr2 118305361 N DEL 19
SRR1766446.7225883 chr2 118305292 N chr2 118305375 N DEL 1
SRR1766459.4666186 chr2 118305162 N chr2 118305372 N DEL 4
SRR1766484.8129889 chr2 118305576 N chr2 118305673 N DEL 1
SRR1766456.2100271 chr2 118305576 N chr2 118305673 N DEL 5
SRR1766473.5963425 chr2 118305590 N chr2 118305663 N DEL 5
SRR1766460.7695086 chr2 118305590 N chr2 118305663 N DEL 5
SRR1766469.10578912 chr2 118305590 N chr2 118305663 N DEL 5
SRR1766463.4270180 chr2 118305590 N chr2 118305663 N DEL 5
SRR1766452.1583991 chr2 118305590 N chr2 118305663 N DEL 6
SRR1766467.6332427 chr2 118305590 N chr2 118305663 N DEL 7
SRR1766485.1656465 chr2 118305590 N chr2 118305663 N DEL 7
SRR1766459.2004797 chr2 118305590 N chr2 118305663 N DEL 9
SRR1766448.9427886 chr2 118305486 N chr2 118305654 N DUP 1
SRR1766450.9287962 chr2 118305695 N chr2 118305758 N DUP 21
SRR1766448.6374881 chr2 118305687 N chr2 118305766 N DUP 15
SRR1766464.10849360 chr2 118305687 N chr2 118305766 N DUP 15
SRR1766445.2480899 chr2 118305687 N chr2 118305766 N DUP 15
SRR1766474.9841002 chr2 118305398 N chr2 118305803 N DEL 5
SRR1766449.4069206 chr2 118305400 N chr2 118305805 N DEL 5
SRR1766461.4805174 chr2 118305590 N chr2 118305809 N DEL 5
SRR1766473.2909757 chr2 118305317 N chr2 118305813 N DEL 4
SRR1766474.11649540 chr2 118305498 N chr2 118305816 N DEL 1
SRR1766444.1566573 chr1 248522890 N chr1 248522991 N DEL 25
SRR1766485.7484538 chr16 48932387 N chr16 48932500 N DUP 16
SRR1766449.6517976 chr1 87636067 N chr1 87636229 N DEL 6
SRR1766465.7601568 chr2 105210573 N chr2 105211248 N DEL 7
SRR1766485.6766333 chr2 105210653 N chr2 105211248 N DEL 5
SRR1766465.10610913 chr2 105210596 N chr2 105210995 N DEL 5
SRR1766449.8992807 chr2 105210575 N chr2 105211118 N DUP 6
SRR1766454.2122006 chr2 105210575 N chr2 105211118 N DUP 6
SRR1766455.3653124 chr2 105210436 N chr2 105211011 N DEL 1
SRR1766446.7067725 chr2 105210750 N chr2 105211118 N DUP 6
SRR1766443.1631790 chr2 105210750 N chr2 105211118 N DUP 6
SRR1766459.9185262 chr2 105210750 N chr2 105211118 N DUP 6
SRR1766447.9766573 chr2 105210449 N chr2 105211025 N DEL 6
SRR1766443.3131790 chr2 105210750 N chr2 105211118 N DUP 6
SRR1766450.7761712 chr2 105210494 N chr2 105211164 N DUP 6
SRR1766471.10349905 chr2 105211081 N chr2 105211207 N DUP 5
SRR1766455.3653124 chr2 105210478 N chr2 105211118 N DEL 10
SRR1766483.12190389 chr2 105211082 N chr2 105211208 N DUP 2
SRR1766478.877785 chr18 79236864 N chr18 79236916 N DEL 5
SRR1766476.4894098 chr18 79236837 N chr18 79237427 N DEL 25
SRR1766464.8327636 chr18 79236985 N chr18 79237044 N DEL 5
SRR1766444.934745 chr18 79236997 N chr18 79237047 N DUP 5
SRR1766468.3782951 chr18 79236901 N chr18 79237004 N DEL 9
SRR1766472.297509 chr18 79237117 N chr18 79237276 N DUP 5
SRR1766452.4880890 chr18 79237117 N chr18 79237276 N DUP 5
SRR1766478.10596275 chr18 79237033 N chr18 79237468 N DUP 5
SRR1766455.4447275 chr18 79237067 N chr18 79237393 N DUP 5
SRR1766481.7362363 chr18 79237007 N chr18 79237117 N DEL 10
SRR1766464.1524448 chr18 79236956 N chr18 79237117 N DEL 10
SRR1766442.2983741 chr18 79236916 N chr18 79237126 N DUP 5
SRR1766479.4990994 chr18 79237167 N chr18 79237335 N DEL 5
SRR1766453.1871095 chr18 79236902 N chr18 79237061 N DUP 5
SRR1766451.4901703 chr18 79236959 N chr18 79237338 N DEL 5
SRR1766471.4802654 chr18 79236902 N chr18 79237061 N DUP 10
SRR1766442.7734551 chr18 79237498 N chr18 79237550 N DEL 5
SRR1766479.456604 chr18 79236885 N chr18 79237475 N DEL 7
SRR1766453.4199231 chr18 79237129 N chr18 79237508 N DEL 30
SRR1766446.4013180 chr18 79236953 N chr18 79237492 N DEL 5
SRR1766474.2101939 chr18 79237069 N chr18 79237499 N DEL 10
SRR1766453.9563237 chr6 108989656 N chr6 108989727 N DEL 5
SRR1766482.6670008 chr6 108989656 N chr6 108989727 N DEL 5
SRR1766474.7149651 chr6 108989675 N chr6 108989744 N DUP 5
SRR1766483.6421710 chr6 30475035 N chr6 30475349 N DEL 1
SRR1766442.37981808 chr6 30475058 N chr6 30475175 N DEL 5
SRR1766472.8521073 chr6 30475237 N chr6 30475312 N DUP 5
SRR1766448.6385855 chr9 65432754 N chr9 65432879 N DEL 5
SRR1766464.8183306 chr3 127154827 N chr3 127154916 N DEL 5
SRR1766476.9625697 chr3 127154836 N chr3 127155123 N DEL 7
SRR1766470.9526081 chr3 127154843 N chr3 127155086 N DEL 11
SRR1766458.5314047 chr3 127154874 N chr3 127155426 N DEL 5
SRR1766484.3576095 chr3 127154928 N chr3 127155029 N DEL 5
SRR1766459.6905542 chr3 127154840 N chr3 127154929 N DUP 8
SRR1766456.3210256 chr3 127154860 N chr3 127155071 N DEL 33
SRR1766485.253810 chr3 127154896 N chr3 127155032 N DUP 1
SRR1766452.3597420 chr3 127155024 N chr3 127155190 N DUP 9
SRR1766481.9682978 chr3 127155110 N chr3 127155184 N DUP 5
SRR1766479.6358088 chr3 127155110 N chr3 127155184 N DUP 7
SRR1766478.6919107 chr3 127155114 N chr3 127155216 N DUP 2
SRR1766485.3178873 chr3 127154835 N chr3 127155197 N DEL 9
SRR1766446.3799978 chr3 127155125 N chr3 127155199 N DEL 9
SRR1766451.3826749 chr3 127154832 N chr3 127155202 N DEL 6
SRR1766453.9507247 chr3 127154832 N chr3 127155202 N DEL 6
SRR1766457.4042045 chr19 8530055 N chr19 8530133 N DEL 5
SRR1766457.6321681 chr19 8529959 N chr19 8530112 N DUP 8
SRR1766476.6071675 chr19 8529971 N chr19 8530049 N DEL 5
SRR1766444.1405123 chr19 8530035 N chr19 8530113 N DEL 5
SRR1766472.9246500 chr19 8530218 N chr19 8530294 N DUP 1
SRR1766472.1171945 chr1 232368459 N chr1 232368722 N DUP 4
SRR1766446.7547004 chr1 232368459 N chr1 232368722 N DUP 15
SRR1766442.26787874 chr19 53990572 N chr19 53990683 N DEL 13
SRR1766466.4360062 chr19 53990662 N chr19 53991210 N DUP 5
SRR1766464.8380183 chr19 53990587 N chr19 53990661 N DEL 9
SRR1766478.7522360 chr19 53990761 N chr19 53991019 N DEL 4
SRR1766479.2543895 chr19 53990717 N chr19 53991050 N DEL 8
SRR1766470.10505792 chr19 53990620 N chr19 53990838 N DUP 21
SRR1766461.10652840 chr19 53990712 N chr19 53990934 N DEL 5
SRR1766448.684865 chr19 53990799 N chr19 53991094 N DEL 2
SRR1766471.6330094 chr19 53991104 N chr19 53991210 N DUP 22
SRR1766442.39206125 chr19 53991199 N chr19 53991271 N DUP 11
SRR1766454.2721593 chr19 53990751 N chr19 53991263 N DEL 17
SRR1766448.9487496 chr19 53990753 N chr19 53991265 N DEL 17
SRR1766455.4415555 chr19 53990716 N chr19 53991265 N DEL 17
SRR1766466.1766866 chr19 53990713 N chr19 53991262 N DEL 13
SRR1766474.6535639 chr19 53990713 N chr19 53991262 N DEL 10
SRR1766445.2330495 chr19 53990713 N chr19 53991262 N DEL 10
SRR1766461.6559010 chr19 53990677 N chr19 53991263 N DEL 10
SRR1766481.4076187 chr19 53990677 N chr19 53991263 N DEL 10
SRR1766447.10637151 chr19 53990944 N chr19 53991273 N DEL 2
SRR1766484.7382337 chr19 53990684 N chr19 53991270 N DEL 7
SRR1766456.5150522 chrX 23523187 N chrX 23523448 N DEL 1
SRR1766486.968210 chrX 23523206 N chrX 23523426 N DUP 5
SRR1766472.9282592 chrX 23523206 N chrX 23523426 N DUP 5
SRR1766484.6688805 chrX 23523206 N chrX 23523426 N DUP 5
SRR1766455.4497613 chrX 23523224 N chrX 23523446 N DEL 5
SRR1766460.6968870 chrX 23523013 N chrX 23523458 N DEL 3
SRR1766442.11489316 chrX 23523383 N chrX 23523497 N DEL 15
SRR1766485.8395553 chrX 23523101 N chrX 23523628 N DEL 5
SRR1766451.6004862 chrX 23523366 N chrX 23523635 N DEL 5
SRR1766446.10628040 chr1 4544775 N chr1 4545055 N DEL 5
SRR1766451.10697768 chr7 145271697 N chr7 145271813 N DUP 4
SRR1766470.4234979 chr7 145271808 N chr7 145271861 N DEL 6
SRR1766474.6870307 chr22 41643842 N chr22 41644169 N DEL 35
SRR1766486.4187846 chr22 41643924 N chr22 41644251 N DEL 4
SRR1766442.27301401 chr22 41643885 N chr22 41644050 N DEL 1
SRR1766459.5029076 chr22 41643971 N chr22 41644134 N DEL 1
SRR1766457.1493023 chr22 41643969 N chr22 41644135 N DEL 6
SRR1766471.7861820 chr3 81229093 N chr3 81229142 N DUP 3
SRR1766471.1800015 chr3 81229093 N chr3 81229142 N DUP 3
SRR1766465.4626733 chr3 81229095 N chr3 81229144 N DUP 1
SRR1766486.4843313 chr3 81229095 N chr3 81229144 N DUP 1
SRR1766473.8342092 chr4 32832214 N chr4 32833166 N DEL 6
SRR1766480.6056627 chr4 32832219 N chr4 32833166 N DEL 7
SRR1766470.2528414 chr4 32832225 N chr4 32833165 N DEL 6
SRR1766442.6552877 chr4 32832228 N chr4 32833166 N DEL 6
SRR1766486.5199326 chr4 32832247 N chr4 32833166 N DEL 5
SRR1766442.11606445 chr4 32832252 N chr4 32833165 N DEL 3
SRR1766442.5389982 chr4 32832260 N chr4 32833166 N DEL 6
SRR1766466.3217265 chr4 32832269 N chr4 32833166 N DEL 5
SRR1766483.7219585 chr4 32832274 N chr4 32833166 N DEL 6
SRR1766484.3123492 chr4 32832240 N chr4 32833166 N DEL 6
SRR1766442.26231870 chr4 32832304 N chr4 32833166 N DEL 4
SRR1766446.7163736 chr4 32832304 N chr4 32833166 N DEL 4
SRR1766443.8547467 chr4 32832309 N chr4 32833165 N DEL 5
SRR1766486.9769863 chr4 32832315 N chr4 32833166 N DEL 5
SRR1766485.3574501 chr4 32832325 N chr4 32833165 N DEL 6
SRR1766473.10152984 chr4 32832329 N chr4 32833165 N DEL 7
SRR1766465.1582654 chr4 32832349 N chr4 32833165 N DEL 5
SRR1766474.4394482 chr4 32832359 N chr4 32833164 N DEL 5
SRR1766442.23934358 chr4 32832367 N chr4 32833166 N DEL 2
SRR1766469.778657 chr4 32832379 N chr4 32833165 N DEL 5
SRR1766442.6552877 chr4 32832393 N chr4 32833165 N DEL 5
SRR1766451.1962529 chr4 32832396 N chr4 32833166 N DEL 5
SRR1766442.2499078 chr4 32832397 N chr4 32833165 N DEL 4
SRR1766452.10655315 chr4 32832402 N chr4 32833166 N DEL 3
SRR1766473.7892062 chr4 32832403 N chr4 32833165 N DEL 4
SRR1766473.10359285 chr4 32832407 N chr4 32833166 N DEL 6
SRR1766465.6103417 chr4 32832419 N chr4 32833163 N DEL 5
SRR1766480.5503759 chr4 32832424 N chr4 32833163 N DEL 2
SRR1766443.8823819 chr4 32832762 N chr4 32833166 N DEL 6
SRR1766483.7219585 chr4 32832575 N chr4 32833179 N DUP 2
SRR1766462.10472022 chr4 32832400 N chr4 32833164 N DEL 2
SRR1766449.4268372 chr4 32832627 N chr4 32833163 N DEL 4
SRR1766442.11606445 chr4 32832676 N chr4 32833165 N DEL 5
SRR1766443.8547467 chr4 32832703 N chr4 32833166 N DEL 6
SRR1766447.2209434 chr4 32832735 N chr4 32833166 N DEL 2
SRR1766471.932094 chr4 32832901 N chr4 32833166 N DEL 2
SRR1766445.8629386 chr4 168793270 N chr4 168793463 N DEL 4
SRR1766469.2643177 chr4 168793270 N chr4 168793463 N DEL 4
SRR1766466.8157034 chr4 168793270 N chr4 168793415 N DEL 1
SRR1766446.6379945 chr4 168793274 N chr4 168793513 N DUP 2
SRR1766445.7249306 chr4 168793274 N chr4 168793511 N DUP 6
SRR1766465.10783745 chr4 168793335 N chr4 168793434 N DEL 11
SRR1766480.4593468 chr4 168793274 N chr4 168793511 N DUP 6
SRR1766486.7550105 chr4 168793290 N chr4 168793359 N DUP 7
SRR1766476.10937606 chr4 168793290 N chr4 168793383 N DUP 7
SRR1766478.11261213 chr4 168793271 N chr4 168793531 N DUP 8
SRR1766475.6601955 chr4 168793271 N chr4 168793531 N DUP 8
SRR1766442.28912190 chr4 168793275 N chr4 168793512 N DUP 6
SRR1766449.4489166 chr4 168793278 N chr4 168793515 N DUP 3
SRR1766480.7373929 chr4 168793278 N chr4 168793515 N DUP 3
SRR1766459.9267253 chr4 168793271 N chr4 168793531 N DUP 8
SRR1766450.6691221 chr4 168793284 N chr4 168793405 N DUP 3
SRR1766454.4535107 chr4 168793277 N chr4 168793514 N DUP 4
SRR1766444.833047 chr4 168793276 N chr4 168793513 N DUP 5
SRR1766464.368907 chr4 168793280 N chr4 168793517 N DUP 1
SRR1766472.1979346 chr4 168793280 N chr4 168793517 N DUP 1
SRR1766442.19867146 chr4 168793271 N chr4 168793531 N DUP 8
SRR1766481.9659482 chr4 168793271 N chr4 168793531 N DUP 8
SRR1766483.11265334 chr4 168793311 N chr4 168793410 N DEL 12
SRR1766472.232346 chr4 168793359 N chr4 168793458 N DEL 11
SRR1766474.2549351 chr4 168793311 N chr4 168793410 N DEL 11
SRR1766474.27397 chr4 168793284 N chr4 168793381 N DEL 1
SRR1766483.1384191 chr4 168793271 N chr4 168793531 N DUP 2
SRR1766466.881151 chr4 168793271 N chr4 168793531 N DUP 3
SRR1766456.2609589 chr4 168793271 N chr4 168793531 N DUP 2
SRR1766463.6135632 chr4 168793391 N chr4 168793510 N DUP 5
SRR1766483.3609025 chr4 168793391 N chr4 168793510 N DUP 5
SRR1766464.3227612 chr4 168793271 N chr4 168793531 N DUP 7
SRR1766459.9212335 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766476.2342203 chr4 168793439 N chr4 168793531 N DUP 8
SRR1766481.2024056 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766442.29952833 chr4 168793271 N chr4 168793531 N DUP 6
SRR1766455.1325294 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766442.8588090 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766467.11788071 chr4 168793418 N chr4 168793516 N DEL 11
SRR1766444.833047 chr4 168793418 N chr4 168793516 N DEL 11
SRR1766463.8305745 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766459.9267253 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766459.9982881 chr4 168793284 N chr4 168793532 N DUP 10
SRR1766445.2189057 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766443.2235559 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766479.2134224 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766486.82444 chr4 168793394 N chr4 168793516 N DEL 11
SRR1766453.8348741 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766481.3212651 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766443.904725 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766466.881151 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766447.598630 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766460.10706412 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766442.19349917 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766443.6213861 chr4 168793370 N chr4 168793516 N DEL 11
SRR1766471.2318564 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766458.2755623 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766449.9613880 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766477.399156 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766454.4999230 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766479.13870801 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766458.2553896 chr4 168793346 N chr4 168793516 N DEL 11
SRR1766450.189355 chr4 168793322 N chr4 168793516 N DEL 11
SRR1766453.6179082 chr4 168793323 N chr4 168793517 N DEL 16
SRR1766479.9068621 chr4 168793322 N chr4 168793516 N DEL 11
SRR1766456.2709829 chr4 168793322 N chr4 168793516 N DEL 11
SRR1766449.5797437 chr4 168793322 N chr4 168793516 N DEL 11
SRR1766442.32762427 chr4 168793298 N chr4 168793516 N DEL 11
SRR1766460.3374870 chr4 168793298 N chr4 168793516 N DEL 11
SRR1766452.3058440 chr4 168793298 N chr4 168793516 N DEL 11
SRR1766479.5943555 chr4 168793298 N chr4 168793516 N DEL 11
SRR1766444.337386 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766445.2863050 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766449.9940941 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766476.11122362 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766452.3617401 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766459.650723 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766482.5621176 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766453.4114526 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766459.951454 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766448.5103897 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766486.271282 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766453.7299465 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766461.3639402 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766481.11652766 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766466.11151667 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766473.10925460 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766467.10518540 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766454.1695624 chr7 158950530 N chr7 158950836 N DEL 5
SRR1766476.868937 chr7 158950530 N chr7 158950836 N DEL 10
SRR1766454.10692326 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766442.10971825 chr7 158950547 N chr7 158950851 N DUP 4
SRR1766481.12326936 chr7 158950547 N chr7 158950851 N DUP 5
SRR1766472.8614289 chr7 158950548 N chr7 158950852 N DUP 4
SRR1766483.625924 chr7 158950549 N chr7 158950853 N DUP 3
SRR1766474.2355428 chr7 158950551 N chr7 158950611 N DUP 1
SRR1766471.2208138 chr7 158950597 N chr7 158951023 N DUP 5
SRR1766444.6055709 chr7 158950597 N chr7 158951023 N DUP 5
SRR1766481.8964949 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766450.7974480 chr7 158950595 N chr7 158950901 N DEL 5
SRR1766478.9747975 chr7 158950597 N chr7 158951023 N DUP 5
SRR1766484.4311807 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766449.9370257 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766476.8781181 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766480.7922883 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766472.2661281 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766480.6223155 chr7 158950597 N chr7 158950840 N DUP 5
SRR1766466.10032301 chr7 158950596 N chr7 158950963 N DEL 5
SRR1766469.4898300 chr7 158950674 N chr7 158950980 N DEL 5
SRR1766465.10853257 chr7 158950622 N chr7 158950928 N DEL 5
SRR1766466.1228450 chr7 158950598 N chr7 158950841 N DUP 5
SRR1766455.2473682 chr7 158950597 N chr7 158950840 N DUP 5
SRR1766447.9729015 chr7 158950719 N chr7 158950840 N DUP 5
SRR1766483.1888008 chr7 158950719 N chr7 158950840 N DUP 5
SRR1766475.3096953 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766446.3407032 chr7 158950719 N chr7 158950840 N DUP 5
SRR1766485.10559442 chr7 158950719 N chr7 158950840 N DUP 5
SRR1766442.29461411 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766443.2101123 chr7 158950720 N chr7 158950841 N DUP 5
SRR1766466.154508 chr7 158950721 N chr7 158950842 N DUP 5
SRR1766477.9266510 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766478.3586655 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766453.2591929 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766462.9903974 chr7 158950674 N chr7 158950980 N DEL 1
SRR1766466.1228450 chr7 158950678 N chr7 158950984 N DEL 1
SRR1766473.144859 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766479.2106849 chr7 158950678 N chr7 158950984 N DEL 3
SRR1766481.2299530 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766480.2994254 chr7 158950674 N chr7 158950980 N DEL 5
SRR1766472.5450819 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766449.1295870 chr7 158950674 N chr7 158950980 N DEL 5
SRR1766473.2591228 chr7 158950674 N chr7 158950980 N DEL 5
SRR1766476.8540581 chr7 158950674 N chr7 158950980 N DEL 5
SRR1766462.3824676 chr7 158950674 N chr7 158950980 N DEL 5
SRR1766470.3627691 chr7 158950674 N chr7 158950980 N DEL 5
SRR1766447.996196 chr7 158950780 N chr7 158950840 N DUP 5
SRR1766485.10611558 chr7 158950920 N chr7 158951041 N DUP 7
SRR1766444.6055709 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766475.6087177 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766459.9278196 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766442.29821866 chr7 158950797 N chr7 158950857 N DUP 10
SRR1766485.9923337 chr7 158950552 N chr7 158950797 N DEL 5
SRR1766473.728576 chr7 158950555 N chr7 158950800 N DEL 5
SRR1766463.7566270 chr7 158950557 N chr7 158950802 N DEL 5
SRR1766473.728576 chr7 158950560 N chr7 158950805 N DEL 5
SRR1766446.3363742 chr7 158950563 N chr7 158950808 N DEL 4
SRR1766446.4283791 chr7 158950563 N chr7 158950808 N DEL 4
SRR1766477.2968863 chr7 158950565 N chr7 158950810 N DEL 2
SRR1766462.1409209 chr7 158950596 N chr7 158950841 N DEL 5
SRR1766467.1292247 chr7 158950779 N chr7 158950900 N DUP 5
SRR1766442.23824068 chr7 158950919 N chr7 158950981 N DEL 4
SRR1766454.10692326 chr7 158950919 N chr7 158950981 N DEL 5
SRR1766484.7252231 chr7 158950919 N chr7 158950981 N DEL 5
SRR1766442.29253855 chr7 158950919 N chr7 158950981 N DEL 5
SRR1766458.8055177 chr7 158950919 N chr7 158950981 N DEL 5
SRR1766443.2244463 chr7 158950595 N chr7 158950901 N DEL 5
SRR1766442.5666344 chr7 158950919 N chr7 158950981 N DEL 5
SRR1766480.7922883 chr7 158950595 N chr7 158950901 N DEL 5
SRR1766469.3037349 chr7 158950921 N chr7 158950983 N DEL 5
SRR1766480.5073724 chr7 158950919 N chr7 158950981 N DEL 5
SRR1766478.9747975 chr7 158950737 N chr7 158950919 N DUP 10
SRR1766482.3346353 chr7 158950614 N chr7 158950920 N DEL 6
SRR1766442.27458637 chr7 158950614 N chr7 158950920 N DEL 5
SRR1766470.9993654 chr7 158950615 N chr7 158950921 N DEL 5
SRR1766467.1131528 chr7 158950616 N chr7 158950922 N DEL 5
SRR1766446.145815 chr7 158950617 N chr7 158950923 N DEL 5
SRR1766442.29461411 chr7 158950559 N chr7 158950924 N DUP 5
SRR1766445.3328767 chr7 158950797 N chr7 158950857 N DUP 9
SRR1766449.8907196 chr7 158950623 N chr7 158950929 N DEL 5
SRR1766475.3099024 chr7 158950797 N chr7 158950857 N DUP 7
SRR1766473.5765480 chr7 158950797 N chr7 158950857 N DUP 6
SRR1766471.11872906 chr7 158950596 N chr7 158950963 N DEL 6
SRR1766485.5853260 chr7 158950797 N chr7 158950857 N DUP 5
SRR1766459.8669783 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766477.8427437 chr7 158950797 N chr7 158950857 N DUP 5
SRR1766476.6112682 chr7 158950797 N chr7 158950857 N DUP 5
SRR1766457.1439474 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766466.11151667 chr7 158950596 N chr7 158950963 N DEL 5
SRR1766483.2640804 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766483.5318081 chr7 158950597 N chr7 158951023 N DUP 5
SRR1766467.4728417 chr7 158950920 N chr7 158951041 N DUP 10
SRR1766473.5765480 chr7 158950605 N chr7 158950972 N DEL 5
SRR1766473.2869778 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766443.680067 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766480.6223155 chr7 158950984 N chr7 158951044 N DUP 5
SRR1766450.7984806 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766474.2949210 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766442.13626128 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766451.763235 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766449.9869448 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766442.13805056 chr7 158950980 N chr7 158951040 N DUP 5
SRR1766464.1044974 chr7 158950613 N chr7 158950980 N DEL 5
SRR1766474.2949210 chr7 158950605 N chr7 158951033 N DEL 5
SRR1766455.3053842 chr7 158950596 N chr7 158951024 N DEL 5
SRR1766482.6796751 chr7 158950596 N chr7 158951024 N DEL 5
SRR1766442.26883389 chr7 158950596 N chr7 158951085 N DEL 5
SRR1766462.7581550 chr17 82009748 N chr17 82009920 N DEL 11
SRR1766457.1322557 chr17 82009753 N chr17 82009807 N DUP 10
SRR1766464.6445769 chr17 82009753 N chr17 82009807 N DUP 26
SRR1766451.650599 chr17 82009740 N chr17 82009910 N DUP 7
SRR1766473.8684139 chr17 82009740 N chr17 82009910 N DUP 5
SRR1766484.3220993 chr17 82009783 N chr17 82009897 N DEL 1
SRR1766465.8748957 chr17 82009759 N chr17 82009931 N DEL 4
SRR1766484.5828129 chr3 26615388 N chr3 26615473 N DUP 2
SRR1766452.9992565 chr19 54770302 N chr19 54770417 N DUP 5
SRR1766455.5388063 chr19 54770300 N chr19 54770415 N DUP 5
SRR1766464.8002664 chr19 54770300 N chr19 54770415 N DUP 6
SRR1766479.12058537 chr19 54770438 N chr19 54770782 N DUP 5
SRR1766473.1521708 chr19 54770317 N chr19 54770453 N DEL 5
SRR1766474.2617036 chr19 54770324 N chr19 54770460 N DEL 5
SRR1766459.8869696 chr19 54770329 N chr19 54770465 N DEL 10
SRR1766469.8213701 chr19 54770300 N chr19 54770608 N DUP 11
SRR1766483.6642310 chr19 54770137 N chr19 54770506 N DEL 5
SRR1766477.8981579 chr19 54770299 N chr19 54770645 N DUP 1
SRR1766479.10274469 chr19 54770331 N chr19 54770563 N DEL 14
SRR1766466.8709599 chr19 54770459 N chr19 54770691 N DEL 15
SRR1766467.1381089 chr19 54770300 N chr19 54770760 N DUP 5
SRR1766442.28179874 chr19 54770684 N chr19 54770742 N DEL 5
SRR1766446.2241319 chr19 54770744 N chr19 54770800 N DUP 5
SRR1766469.8099906 chr19 54770339 N chr19 54770781 N DEL 1
SRR1766479.2018240 chr6 1260975 N chr6 1261191 N DEL 5
SRR1766471.4051835 chr6 1261095 N chr6 1261182 N DEL 5
SRR1766476.2580141 chr6 1261095 N chr6 1261182 N DEL 5
SRR1766468.127886 chr6 1261052 N chr6 1261182 N DEL 5
SRR1766463.7143417 chr17 44984368 N chr17 44984639 N DEL 1
SRR1766485.7290112 chr17 44984359 N chr17 44984657 N DEL 26
SRR1766442.1847651 chr17 44984377 N chr17 44985186 N DUP 5
SRR1766450.9543883 chr17 44984425 N chr17 44985186 N DUP 13
SRR1766442.17220758 chr17 44984407 N chr17 44985189 N DUP 4
SRR1766442.47037598 chr17 44984511 N chr17 44984944 N DEL 5
SRR1766457.66159 chr17 44984539 N chr17 44985186 N DUP 5
SRR1766456.2297768 chr17 44984562 N chr17 44985182 N DUP 5
SRR1766486.1201177 chr17 44984576 N chr17 44984629 N DUP 5
SRR1766444.361851 chr17 44984558 N chr17 44985178 N DUP 5
SRR1766478.2121904 chr17 44984590 N chr17 44985327 N DUP 14
SRR1766452.10612735 chr17 44984661 N chr17 44984905 N DEL 5
SRR1766480.7793587 chr17 44984600 N chr17 44985229 N DUP 10
SRR1766451.10557192 chr17 44984600 N chr17 44985166 N DUP 5
SRR1766469.695442 chr17 44984652 N chr17 44985281 N DUP 1
SRR1766475.6886038 chr17 44984627 N chr17 44984680 N DUP 5
SRR1766466.4008558 chr17 44984603 N chr17 44984656 N DUP 5
SRR1766469.2935742 chr17 44984707 N chr17 44985140 N DEL 15
SRR1766463.7427346 chr17 44984359 N chr17 44984630 N DEL 11
SRR1766485.4748013 chr17 44984616 N chr17 44984693 N DUP 8
SRR1766452.4228250 chr17 44984429 N chr17 44984646 N DEL 5
SRR1766462.9127446 chr17 44984706 N chr17 44985200 N DUP 2
SRR1766464.4736827 chr17 44984390 N chr17 44984607 N DEL 5
SRR1766466.10414297 chr17 44984668 N chr17 44985020 N DEL 5
SRR1766447.7352218 chr17 44984749 N chr17 44985270 N DUP 16
SRR1766482.4546937 chr17 44984644 N chr17 44985156 N DUP 10
SRR1766466.2394144 chr17 44984909 N chr17 44985268 N DUP 10
SRR1766457.914526 chr17 44984774 N chr17 44985178 N DUP 10
SRR1766479.5121013 chr17 44984670 N chr17 44984806 N DEL 5
SRR1766450.5937451 chr17 44984585 N chr17 44985178 N DUP 11
SRR1766482.11531981 chr17 44984782 N chr17 44985186 N DUP 5
SRR1766450.9361324 chr17 44984668 N chr17 44985020 N DEL 5
SRR1766465.2637815 chr17 44984689 N chr17 44985212 N DEL 5
SRR1766443.6165460 chr17 44985267 N chr17 44985370 N DEL 9
SRR1766442.10596442 chr17 44984692 N chr17 44985242 N DEL 13
SRR1766456.1143039 chr17 44984734 N chr17 44985257 N DEL 30
SRR1766478.6794463 chr17 44984680 N chr17 44985284 N DEL 10
SRR1766464.8921506 chr17 44984653 N chr17 44985257 N DEL 18
SRR1766442.41162515 chr17 44984689 N chr17 44985266 N DEL 1
SRR1766479.1288029 chr17 44985188 N chr17 44985282 N DEL 8
SRR1766477.3929566 chr17 44985184 N chr17 44985302 N DEL 10
SRR1766464.6843622 chrY 10646342 N chrY 10646672 N DEL 10
SRR1766463.7510430 chr10 102637739 N chr10 102637791 N DUP 20
SRR1766471.4373513 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766442.33495784 chr10 102637463 N chr10 102637662 N DEL 7
SRR1766463.4328658 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766465.9847987 chr10 102637416 N chr10 102637532 N DUP 12
SRR1766442.1763377 chr10 102637718 N chr10 102637807 N DUP 11
SRR1766474.9837836 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766453.3178474 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766466.5791553 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766463.1209469 chr10 102637560 N chr10 102638339 N DEL 3
SRR1766483.11979038 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766486.1512701 chr10 102637463 N chr10 102637662 N DEL 7
SRR1766464.960101 chr10 102637701 N chr10 102637823 N DUP 14
SRR1766477.7700857 chr10 102637701 N chr10 102637790 N DUP 35
SRR1766442.11737665 chr10 102637509 N chr10 102637970 N DUP 6
SRR1766476.2983707 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766458.4327978 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766455.8706349 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766442.33831480 chr10 102637543 N chr10 102638046 N DEL 5
SRR1766442.7307863 chr10 102637739 N chr10 102637791 N DUP 23
SRR1766449.10509094 chr10 102637739 N chr10 102637833 N DUP 21
SRR1766442.33601028 chr10 102637739 N chr10 102637833 N DUP 16
SRR1766472.8515428 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766482.743722 chr10 102637538 N chr10 102637783 N DUP 3
SRR1766472.4239913 chr10 102637740 N chr10 102637797 N DUP 14
SRR1766465.7725181 chr10 102637718 N chr10 102637807 N DUP 11
SRR1766480.8729074 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766461.2338778 chr10 102637739 N chr10 102637791 N DUP 31
SRR1766447.535015 chr10 102637532 N chr10 102637807 N DUP 8
SRR1766442.39982411 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766471.7997679 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766459.7466408 chr10 102637739 N chr10 102637833 N DUP 19
SRR1766452.4617588 chr10 102637420 N chr10 102637535 N DUP 8
SRR1766477.2807594 chr10 102637756 N chr10 102637820 N DEL 1
SRR1766442.45623447 chr10 102637740 N chr10 102637834 N DUP 6
SRR1766484.6987771 chr10 102637408 N chr10 102637487 N DUP 7
SRR1766453.9605507 chr20 63466387 N chr20 63466437 N DUP 5
SRR1766447.10854112 chrX 35600780 N chrX 35600893 N DEL 5
SRR1766459.1232431 chrX 35600780 N chrX 35600893 N DEL 7
SRR1766473.714143 chrX 35600821 N chrX 35601037 N DUP 9
SRR1766445.3651237 chrX 35600911 N chrX 35601011 N DUP 14
SRR1766450.4639613 chrX 35600886 N chrX 35601030 N DUP 10
SRR1766454.1716095 chrX 35600965 N chrX 35601054 N DUP 7
SRR1766470.5548123 chrX 35600889 N chrX 35601037 N DUP 14
SRR1766474.11734541 chrX 35600965 N chrX 35601054 N DUP 6
SRR1766473.714143 chrX 35600898 N chrX 35601070 N DUP 14
SRR1766458.1716387 chrX 35600936 N chrX 35601011 N DUP 17
SRR1766465.2637436 chrX 35600939 N chrX 35601007 N DUP 12
SRR1766480.1051086 chrX 35600939 N chrX 35601007 N DUP 11
SRR1766442.17847578 chrX 35600949 N chrX 35601017 N DUP 19
SRR1766453.4492762 chrX 35600785 N chrX 35601017 N DUP 3
SRR1766463.7851643 chrX 35600765 N chrX 35601007 N DUP 6
SRR1766452.10449664 chrX 35600972 N chrX 35601077 N DUP 18
SRR1766481.13043448 chrX 35600897 N chrX 35601030 N DUP 9
SRR1766456.1325496 chrX 35600897 N chrX 35601030 N DUP 9
SRR1766442.11179291 chrX 35600897 N chrX 35601030 N DUP 10
SRR1766459.4268173 chrX 35600887 N chrX 35601054 N DUP 13
SRR1766449.2498364 chrX 35600910 N chrX 35600987 N DUP 5
SRR1766465.4433618 chrX 35600886 N chrX 35600940 N DUP 5
SRR1766442.30999057 chrX 35600949 N chrX 35601006 N DUP 16
SRR1766449.7845810 chrX 35600780 N chrX 35600948 N DEL 2
SRR1766484.415740 chrX 35600949 N chrX 35601006 N DUP 16
SRR1766451.4261790 chrX 35600981 N chrX 35601095 N DUP 17
SRR1766469.8810954 chrX 35600974 N chrX 35601135 N DUP 10
SRR1766446.1977179 chrX 35600927 N chrX 35600986 N DUP 11
SRR1766446.3687907 chrX 35600927 N chrX 35600986 N DUP 11
SRR1766473.9910788 chrX 35600914 N chrX 35600969 N DUP 17
SRR1766474.7604554 chrX 35600949 N chrX 35601010 N DUP 16
SRR1766462.4034393 chrX 35600925 N chrX 35601009 N DUP 11
SRR1766451.9365831 chrX 35600749 N chrX 35601086 N DUP 9
SRR1766483.7203161 chrX 35600821 N chrX 35601085 N DUP 8
SRR1766466.4113245 chrX 35600889 N chrX 35601079 N DUP 7
SRR1766443.6370100 chrX 35600785 N chrX 35600944 N DEL 9
SRR1766444.4355655 chrX 35600992 N chrX 35601085 N DUP 7
SRR1766457.4979407 chrX 35600873 N chrX 35600944 N DEL 13
SRR1766472.10109703 chrX 35600785 N chrX 35600944 N DEL 9
SRR1766452.2239816 chrX 35600789 N chrX 35600928 N DEL 16
SRR1766449.8215278 chrX 35600913 N chrX 35601041 N DUP 10
SRR1766442.36879467 chrX 35600888 N chrX 35601021 N DUP 19
SRR1766443.7143205 chrX 35600919 N chrX 35601063 N DUP 5
SRR1766465.3701226 chrX 35600919 N chrX 35601063 N DUP 7
SRR1766463.4124714 chrX 35600919 N chrX 35601063 N DUP 12
SRR1766475.8228710 chrX 35600919 N chrX 35601063 N DUP 18
SRR1766485.3403172 chrX 35600919 N chrX 35601063 N DUP 19
SRR1766474.6117537 chrX 35600765 N chrX 35601085 N DUP 15
SRR1766442.3020537 chrX 35600936 N chrX 35601025 N DEL 9
SRR1766486.1973818 chrX 35600936 N chrX 35601025 N DEL 9
SRR1766452.7849988 chrX 35600936 N chrX 35601025 N DEL 9
SRR1766461.355423 chrX 35600936 N chrX 35601025 N DEL 9
SRR1766477.5700268 chrX 35600936 N chrX 35601034 N DEL 6
SRR1766476.93414 chrX 35600938 N chrX 35601036 N DEL 4
SRR1766455.779315 chr16 17167631 N chr16 17167787 N DEL 5
SRR1766465.1754152 chr16 17167628 N chr16 17167753 N DEL 10
SRR1766452.42900 chr16 17167570 N chr16 17167662 N DUP 5
SRR1766478.1056753 chr16 17167662 N chr16 17167725 N DEL 5
SRR1766485.2798648 chr16 17167662 N chr16 17167725 N DEL 5
SRR1766483.1193136 chr16 17167662 N chr16 17167725 N DEL 10
SRR1766465.8383353 chr16 17167662 N chr16 17167725 N DEL 10
SRR1766455.9858731 chr16 17167562 N chr16 17167685 N DUP 15
SRR1766446.2438935 chr16 17167662 N chr16 17167725 N DEL 10
SRR1766455.9858804 chr16 17167562 N chr16 17167716 N DUP 10
SRR1766478.5075514 chr16 17167567 N chr16 17167721 N DUP 5
SRR1766451.1366538 chr16 17167722 N chr16 17167783 N DUP 5
SRR1766479.6327442 chr16 17167753 N chr16 17167814 N DUP 10
SRR1766442.3797846 chr16 17167722 N chr16 17167783 N DUP 5
SRR1766458.9053629 chr16 17167628 N chr16 17167753 N DEL 13
SRR1766469.1850529 chr16 17167597 N chr16 17167722 N DEL 5
SRR1766444.3103207 chr16 17167799 N chr16 17167862 N DEL 15
SRR1766454.9187347 chr16 17167605 N chr16 17167730 N DEL 5
SRR1766472.3250424 chr16 17167843 N chr16 17167999 N DEL 19
SRR1766470.3765744 chr16 17167862 N chr16 17168018 N DEL 5
SRR1766447.5680734 chr16 17167772 N chr16 17167926 N DUP 5
SRR1766454.9788577 chr16 17167887 N chr16 17167981 N DEL 5
SRR1766471.3883007 chr16 17167631 N chr16 17167818 N DEL 5
SRR1766455.779315 chr16 17167613 N chr16 17167862 N DEL 10
SRR1766477.485333 chr16 17167582 N chr16 17167862 N DEL 8
SRR1766448.5117871 chr16 17167583 N chr16 17167863 N DEL 5
SRR1766454.796036 chr16 17167588 N chr16 17167868 N DEL 5
SRR1766447.3031845 chr16 17167588 N chr16 17167992 N DEL 4
SRR1766472.7347093 chr7 105433769 N chr7 105433905 N DEL 19
SRR1766471.1720986 chr7 105434345 N chr7 105434508 N DUP 5
SRR1766446.3426805 chr18 13946676 N chr18 13946857 N DEL 7
SRR1766457.6445179 chr18 13946676 N chr18 13946857 N DEL 7
SRR1766477.4480609 chr11 101629020 N chr11 101629084 N DUP 22
SRR1766445.1717709 chr11 101629020 N chr11 101629084 N DUP 19
SRR1766480.6373995 chr5 43136625 N chr5 43136798 N DUP 2
SRR1766480.118460 chr5 43136640 N chr5 43136801 N DEL 11
SRR1766446.1718874 chr5 43136644 N chr5 43136806 N DEL 7
SRR1766478.10581363 chr5 43136640 N chr5 43136808 N DEL 6
SRR1766472.1542771 chr7 57182354 N chr7 57182459 N DUP 5
SRR1766460.493980 chr7 57182354 N chr7 57182459 N DUP 5
SRR1766475.756274 chr2 152590090 N chr2 152590157 N DUP 22
SRR1766448.8068102 chr11 71362100 N chr11 71362485 N DEL 13
SRR1766442.17665723 chr11 71362165 N chr11 71363037 N DEL 15
SRR1766451.6611787 chr11 71362191 N chr11 71363167 N DEL 3
SRR1766473.5157919 chr11 71362222 N chr11 71362671 N DEL 14
SRR1766442.18334665 chr11 71362239 N chr11 71362959 N DEL 5
SRR1766483.7914222 chr11 71362227 N chr11 71363171 N DEL 5
SRR1766447.5894118 chr11 71362257 N chr11 71362658 N DEL 16
SRR1766449.4645274 chr11 71362227 N chr11 71362939 N DEL 10
SRR1766461.2314969 chr11 71362243 N chr11 71362931 N DEL 5
SRR1766478.3681812 chr11 71362293 N chr11 71362933 N DEL 4
SRR1766451.8700734 chr11 71362293 N chr11 71362933 N DEL 5
SRR1766457.2548201 chr11 71362305 N chr11 71362658 N DEL 5
SRR1766465.10284368 chr11 71362305 N chr11 71362658 N DEL 5
SRR1766454.4259208 chr11 71362305 N chr11 71362658 N DEL 5
SRR1766442.24254785 chr11 71362305 N chr11 71362658 N DEL 5
SRR1766465.11210800 chr11 71362307 N chr11 71362995 N DEL 15
SRR1766475.8749751 chr11 71362308 N chr11 71362365 N DEL 5
SRR1766476.3235695 chr11 71362311 N chr11 71362408 N DEL 5
SRR1766466.5005942 chr11 71362305 N chr11 71362658 N DEL 10
SRR1766449.10492512 chr11 71362309 N chr11 71362574 N DEL 4
SRR1766471.9152596 chr11 71362311 N chr11 71362408 N DEL 14
SRR1766442.27533844 chr11 71362343 N chr11 71363366 N DEL 20
SRR1766453.2986693 chr11 71362343 N chr11 71363159 N DEL 25
SRR1766464.7570945 chr11 71362327 N chr11 71362807 N DEL 13
SRR1766446.4475112 chr11 71362188 N chr11 71362411 N DUP 5
SRR1766478.3259748 chr11 71362316 N chr11 71362954 N DUP 5
SRR1766442.28290113 chr11 71362197 N chr11 71362326 N DEL 5
SRR1766447.11179387 chr11 71362198 N chr11 71362327 N DEL 4
SRR1766454.9971722 chr11 71362200 N chr11 71362329 N DEL 2
SRR1766456.861808 chr11 71362439 N chr11 71363109 N DUP 45
SRR1766470.1359243 chr11 71362415 N chr11 71363374 N DEL 5
SRR1766449.2647419 chr11 71362461 N chr11 71363356 N DEL 11
SRR1766448.2289497 chr11 71362471 N chr11 71362919 N DEL 9
SRR1766461.9928101 chr11 71362487 N chr11 71363358 N DEL 7
SRR1766478.3458102 chr11 71362495 N chr11 71362871 N DEL 5
SRR1766470.3575750 chr11 71362509 N chr11 71362965 N DEL 15
SRR1766460.1980267 chr11 71362515 N chr11 71362851 N DEL 14
SRR1766473.1606098 chr11 71362495 N chr11 71362871 N DEL 5
SRR1766471.850228 chr11 71362495 N chr11 71363151 N DEL 1
SRR1766471.2296894 chr11 71362497 N chr11 71363321 N DEL 7
SRR1766460.5861818 chr11 71362497 N chr11 71363321 N DEL 18
SRR1766467.5103498 chr11 71362164 N chr11 71362429 N DEL 5
SRR1766458.1408391 chr11 71362378 N chr11 71362443 N DEL 7
SRR1766472.10784921 chr11 71362464 N chr11 71362886 N DUP 11
SRR1766482.10824207 chr11 71362446 N chr11 71362565 N DUP 5
SRR1766445.727329 chr11 71362549 N chr11 71362662 N DEL 10
SRR1766443.2128645 chr11 71362211 N chr11 71362452 N DEL 2
SRR1766449.5479671 chr11 71362472 N chr11 71362870 N DUP 13
SRR1766482.7754462 chr11 71362559 N chr11 71363374 N DEL 5
SRR1766475.10654974 chr11 71362198 N chr11 71362471 N DEL 5
SRR1766456.4229224 chr11 71362543 N chr11 71362823 N DEL 15
SRR1766460.3720636 chr11 71362567 N chr11 71362815 N DEL 6
SRR1766467.7172944 chr11 71362569 N chr11 71362658 N DEL 15
SRR1766446.5774531 chr11 71362569 N chr11 71362658 N DEL 16
SRR1766455.8453985 chr11 71362551 N chr11 71363366 N DEL 8
SRR1766464.9570163 chr11 71362513 N chr11 71362991 N DUP 15
SRR1766450.9876851 chr11 71362496 N chr11 71362894 N DUP 9
SRR1766485.5978334 chr11 71362190 N chr11 71362597 N DUP 10
SRR1766466.7963314 chr11 71362490 N chr11 71362673 N DUP 3
SRR1766459.9383911 chr11 71362527 N chr11 71363436 N DUP 22
SRR1766474.6302661 chr11 71362527 N chr11 71363436 N DUP 22
SRR1766442.33072783 chr11 71362583 N chr11 71363167 N DEL 14
SRR1766469.2613072 chr11 71362214 N chr11 71362511 N DEL 15
SRR1766468.5177052 chr11 71362524 N chr11 71362834 N DUP 15
SRR1766465.5169907 chr11 71362591 N chr11 71362871 N DEL 12
SRR1766478.4976335 chr11 71362342 N chr11 71362511 N DEL 10
SRR1766484.9064412 chr11 71362529 N chr11 71363207 N DUP 24
SRR1766445.8402921 chr11 71362529 N chr11 71362903 N DUP 12
SRR1766446.4771634 chr11 71362526 N chr11 71362836 N DUP 20
SRR1766466.2328616 chr11 71362524 N chr11 71362834 N DUP 15
SRR1766448.9344259 chr11 71362621 N chr11 71362853 N DEL 5
SRR1766450.8117858 chr11 71362621 N chr11 71363388 N DEL 5
SRR1766460.7385137 chr11 71362605 N chr11 71362965 N DEL 10
SRR1766480.2108999 chr11 71362560 N chr11 71362687 N DUP 23
SRR1766481.5419689 chr11 71362205 N chr11 71362550 N DEL 10
SRR1766485.9379500 chr11 71362560 N chr11 71362695 N DUP 10
SRR1766482.10144820 chr11 71362202 N chr11 71362571 N DEL 3
SRR1766450.9315424 chr11 71362685 N chr11 71363356 N DEL 15
SRR1766479.12672498 chr11 71362236 N chr11 71362613 N DEL 17
SRR1766442.12162768 chr11 71362365 N chr11 71362700 N DUP 15
SRR1766485.7538658 chr11 71362652 N chr11 71363058 N DUP 25
SRR1766478.3558518 chr11 71362679 N chr11 71363159 N DEL 15
SRR1766472.5416717 chr11 71362636 N chr11 71362890 N DUP 15
SRR1766469.1259714 chr11 71362639 N chr11 71362893 N DUP 20
SRR1766449.6633775 chr11 71362636 N chr11 71362890 N DUP 15
SRR1766446.7138424 chr11 71362212 N chr11 71362621 N DEL 5
SRR1766479.13270635 chr11 71362639 N chr11 71362893 N DUP 9
SRR1766473.5110401 chr11 71362326 N chr11 71362639 N DEL 10
SRR1766470.4431211 chr11 71362756 N chr11 71362917 N DEL 5
SRR1766474.4577651 chr11 71362641 N chr11 71363079 N DUP 10
SRR1766486.4408733 chr11 71362652 N chr11 71362882 N DUP 5
SRR1766486.917352 chr11 71362652 N chr11 71362986 N DUP 10
SRR1766482.12080067 chr11 71362454 N chr11 71362647 N DEL 7
SRR1766484.4953417 chr11 71362214 N chr11 71362655 N DEL 10
SRR1766472.10343707 chr11 71362287 N chr11 71362664 N DEL 3
SRR1766479.5114827 chr11 71362802 N chr11 71363442 N DEL 5
SRR1766485.9033971 chr11 71362658 N chr11 71362824 N DUP 10
SRR1766444.1552354 chr11 71362192 N chr11 71362854 N DUP 5
SRR1766485.8281298 chr11 71362868 N chr11 71363157 N DEL 5
SRR1766447.11179387 chr11 71362587 N chr11 71362779 N DEL 10
SRR1766459.10823652 chr11 71362335 N chr11 71362767 N DEL 5
SRR1766470.5845601 chr11 71362878 N chr11 71362967 N DEL 9
SRR1766471.10629522 chr11 71362807 N chr11 71362870 N DUP 4
SRR1766477.11320401 chr11 71362459 N chr11 71362795 N DEL 22
SRR1766481.5258286 chr11 71362868 N chr11 71363157 N DEL 13
SRR1766466.1682812 chr11 71362862 N chr11 71362975 N DEL 20
SRR1766482.6952144 chr11 71362559 N chr11 71362861 N DUP 10
SRR1766446.4475112 chr11 71362619 N chr11 71362787 N DEL 10
SRR1766466.6559651 chr11 71362897 N chr11 71363186 N DEL 13
SRR1766473.1464989 chr11 71362894 N chr11 71363175 N DEL 15
SRR1766446.7945186 chr11 71362571 N chr11 71362897 N DUP 2
SRR1766445.6337357 chr11 71362897 N chr11 71363385 N DEL 5
SRR1766453.2445991 chr11 71362659 N chr11 71362897 N DUP 10
SRR1766466.10304556 chr11 71362406 N chr11 71362916 N DUP 5
SRR1766461.8189875 chr11 71362205 N chr11 71362813 N DEL 13
SRR1766452.7927641 chr11 71362213 N chr11 71362813 N DEL 15
SRR1766469.10943672 chr11 71362460 N chr11 71362796 N DEL 9
SRR1766472.7236773 chr11 71362210 N chr11 71362818 N DEL 5
SRR1766457.2138614 chr11 71362813 N chr11 71362988 N DUP 11
SRR1766452.2485757 chr11 71362184 N chr11 71362926 N DUP 5
SRR1766470.6829964 chr11 71362664 N chr11 71362926 N DUP 5
SRR1766485.6125841 chr11 71362942 N chr11 71363159 N DEL 4
SRR1766471.850228 chr11 71362845 N chr11 71363403 N DUP 5
SRR1766470.1359243 chr11 71362855 N chr11 71363166 N DUP 10
SRR1766470.4415029 chr11 71362972 N chr11 71363157 N DEL 2
SRR1766484.8698302 chr11 71362863 N chr11 71363206 N DUP 15
SRR1766461.2314969 chr11 71362199 N chr11 71362871 N DEL 5
SRR1766446.3196653 chr11 71362184 N chr11 71362990 N DUP 11
SRR1766456.1307408 chr11 71362901 N chr11 71363188 N DUP 15
SRR1766473.1332290 chr11 71362201 N chr11 71362897 N DEL 5
SRR1766459.10587405 chr11 71362455 N chr11 71362903 N DEL 5
SRR1766477.10958934 chr11 71362918 N chr11 71363181 N DUP 11
SRR1766442.32474973 chr11 71362494 N chr11 71362918 N DEL 5
SRR1766465.11210800 chr11 71362207 N chr11 71362927 N DEL 15
SRR1766473.1606098 chr11 71362200 N chr11 71362920 N DEL 5
SRR1766466.5005942 chr11 71362698 N chr11 71362938 N DEL 20
SRR1766460.5861818 chr11 71362848 N chr11 71362929 N DEL 4
SRR1766459.5240387 chr11 71362200 N chr11 71363046 N DUP 1
SRR1766467.5595986 chr11 71362426 N chr11 71362938 N DEL 10
SRR1766443.8525842 chr11 71362304 N chr11 71363054 N DUP 5
SRR1766442.12162768 chr11 71362939 N chr11 71363010 N DUP 1
SRR1766471.2296894 chr11 71362674 N chr11 71362938 N DEL 10
SRR1766442.4336325 chr11 71362215 N chr11 71362959 N DEL 10
SRR1766459.5943714 chr11 71363061 N chr11 71363501 N DEL 5
SRR1766451.5112281 chr11 71362202 N chr11 71362946 N DEL 5
SRR1766456.4229224 chr11 71362214 N chr11 71362950 N DEL 8
SRR1766448.9344259 chr11 71362965 N chr11 71363188 N DUP 12
SRR1766472.6742305 chr11 71362215 N chr11 71362959 N DEL 5
SRR1766442.29131103 chr11 71363010 N chr11 71363081 N DUP 10
SRR1766470.4099495 chr11 71362938 N chr11 71363065 N DUP 5
SRR1766442.25539265 chr11 71362658 N chr11 71363072 N DUP 8
SRR1766448.2289497 chr11 71363031 N chr11 71363110 N DUP 17
SRR1766455.8415563 chr11 71363010 N chr11 71363081 N DUP 10
SRR1766475.4023532 chr11 71362842 N chr11 71362995 N DEL 11
SRR1766474.6510952 chr11 71362938 N chr11 71363065 N DUP 5
SRR1766474.6981653 chr11 71362699 N chr11 71362995 N DEL 8
SRR1766457.4792320 chr11 71363086 N chr11 71363167 N DEL 7
SRR1766453.7954749 chr11 71362698 N chr11 71363010 N DEL 15
SRR1766461.3964281 chr11 71363010 N chr11 71363065 N DUP 5
SRR1766484.9911170 chr11 71362330 N chr11 71363010 N DEL 5
SRR1766459.916242 chr11 71363010 N chr11 71363345 N DUP 10
SRR1766483.7914222 chr11 71362203 N chr11 71363011 N DEL 5
SRR1766442.27533844 chr11 71362213 N chr11 71363013 N DEL 10
SRR1766452.10412259 chr11 71363118 N chr11 71363374 N DEL 11
SRR1766458.7519955 chr11 71362658 N chr11 71363128 N DUP 5
SRR1766450.8117858 chr11 71362677 N chr11 71363037 N DEL 5
SRR1766463.5234507 chr11 71362886 N chr11 71363047 N DEL 20
SRR1766445.3357383 chr11 71363067 N chr11 71363385 N DUP 15
SRR1766482.6952144 chr11 71362205 N chr11 71363045 N DEL 5
SRR1766475.4358429 chr11 71362664 N chr11 71363142 N DUP 15
SRR1766472.9810353 chr11 71363148 N chr11 71363253 N DEL 3
SRR1766481.6645569 chr11 71363148 N chr11 71363253 N DEL 5
SRR1766465.499719 chr11 71362478 N chr11 71363164 N DUP 5
SRR1766482.7754462 chr11 71362198 N chr11 71363070 N DEL 5
SRR1766447.10981121 chr11 71363093 N chr11 71363403 N DUP 9
SRR1766484.3690769 chr11 71363151 N chr11 71363296 N DEL 15
SRR1766480.3540835 chr11 71363166 N chr11 71363436 N DUP 18
SRR1766445.7582500 chr11 71363097 N chr11 71363154 N DEL 10
SRR1766460.7385137 chr11 71363085 N chr11 71363204 N DUP 1
SRR1766485.1435462 chr11 71362185 N chr11 71363183 N DUP 12
SRR1766479.4077893 chr11 71363200 N chr11 71363265 N DEL 5
SRR1766442.34935350 chr11 71363196 N chr11 71363261 N DEL 5
SRR1766454.4259208 chr11 71362990 N chr11 71363167 N DEL 31
SRR1766471.10629522 chr11 71362988 N chr11 71363149 N DEL 16
SRR1766471.7148702 chr11 71362986 N chr11 71363163 N DEL 18
SRR1766478.3655375 chr11 71362938 N chr11 71363209 N DUP 12
SRR1766486.1892815 chr11 71363159 N chr11 71363214 N DUP 26
SRR1766442.33072783 chr11 71362866 N chr11 71363163 N DEL 26
SRR1766473.3677126 chr11 71363095 N chr11 71363152 N DEL 10
SRR1766453.7352481 chr11 71362996 N chr11 71363235 N DUP 2
SRR1766477.6075709 chr11 71362814 N chr11 71363181 N DUP 22
SRR1766444.1552354 chr11 71362843 N chr11 71363148 N DEL 10
SRR1766442.25317029 chr11 71362965 N chr11 71363252 N DUP 7
SRR1766442.13375828 chr11 71362858 N chr11 71363249 N DUP 5
SRR1766470.6829964 chr11 71362204 N chr11 71363164 N DEL 10
SRR1766446.7945186 chr11 71362988 N chr11 71363157 N DEL 16
SRR1766457.5192195 chr11 71362197 N chr11 71363165 N DEL 9
SRR1766466.1682812 chr11 71363191 N chr11 71363397 N DUP 5
SRR1766467.2515553 chr11 71363159 N chr11 71363278 N DUP 12
SRR1766476.10202326 chr11 71362672 N chr11 71363192 N DEL 5
SRR1766447.1172997 chr11 71362893 N chr11 71363222 N DEL 10
SRR1766453.2384033 chr11 71363149 N chr11 71363292 N DUP 5
SRR1766455.4595522 chr11 71362090 N chr11 71363202 N DEL 4
SRR1766466.6559651 chr11 71363261 N chr11 71363427 N DUP 15
SRR1766476.9714925 chr11 71363222 N chr11 71363285 N DUP 5
SRR1766467.1238712 chr11 71362382 N chr11 71363222 N DEL 10
SRR1766478.3558518 chr11 71362690 N chr11 71363250 N DEL 12
SRR1766468.1656437 chr11 71362205 N chr11 71363245 N DEL 5
SRR1766470.4099495 chr11 71363202 N chr11 71363283 N DEL 5
SRR1766444.5716179 chr11 71362965 N chr11 71363332 N DUP 32
SRR1766450.8030381 chr11 71363185 N chr11 71363282 N DEL 12
SRR1766484.11211100 chr11 71363203 N chr11 71363284 N DEL 10
SRR1766469.9045967 chr11 71362992 N chr11 71363281 N DEL 9
SRR1766455.8453985 chr11 71362215 N chr11 71363295 N DEL 10
SRR1766443.8525842 chr11 71363086 N chr11 71363366 N DEL 17
SRR1766449.2647419 chr11 71363197 N chr11 71363365 N DEL 6
SRR1766470.4431211 chr11 71362382 N chr11 71363405 N DEL 5
SRR1766445.2362630 chr11 71362204 N chr11 71363411 N DEL 5
SRR1766446.3196653 chr11 71362337 N chr11 71363416 N DEL 4
SRR1766468.7089761 chr11 71362378 N chr11 71363425 N DEL 2
SRR1766486.1591932 chr11 71362483 N chr11 71363458 N DEL 5
SRR1766484.4001374 chr19 55530605 N chr19 55530942 N DEL 3
SRR1766445.3103884 chr19 55530597 N chr19 55530934 N DEL 11
SRR1766443.10812473 chr6 95502056 N chr6 95502163 N DUP 18
SRR1766473.6699064 chr6 95502056 N chr6 95502163 N DUP 19
SRR1766442.21787624 chr6 95502075 N chr6 95502146 N DUP 18
SRR1766442.2535608 chr6 95502075 N chr6 95502146 N DUP 20
SRR1766445.7045337 chr6 95502145 N chr6 95502198 N DEL 34
SRR1766477.2963336 chr6 95502145 N chr6 95502198 N DEL 34
SRR1766463.1810392 chr6 95502102 N chr6 95502247 N DEL 12
SRR1766454.2697701 chr6 95502109 N chr6 95502198 N DEL 34
SRR1766461.9654485 chr6 95502237 N chr6 95502350 N DEL 5
SRR1766475.1562888 chr6 95502237 N chr6 95502350 N DEL 6
SRR1766477.7491277 chr6 95502321 N chr6 95502407 N DEL 6
SRR1766469.10892917 chr6 95502060 N chr6 95502332 N DUP 16
SRR1766452.3848279 chr6 95502225 N chr6 95502310 N DUP 18
SRR1766450.6146715 chr6 95502108 N chr6 95502329 N DUP 4
SRR1766465.812864 chr6 95502326 N chr6 95502414 N DEL 16
SRR1766443.9439229 chr6 95502263 N chr6 95502324 N DUP 17
SRR1766473.4780268 chr6 95502356 N chr6 95502417 N DEL 21
SRR1766455.9427814 chr6 95502060 N chr6 95502129 N DUP 25
SRR1766478.5601427 chr6 95502040 N chr6 95502569 N DUP 26
SRR1766445.325905 chr6 95502263 N chr6 95502324 N DUP 17
SRR1766460.9195407 chr6 95502087 N chr6 95502413 N DEL 8
SRR1766455.9427814 chr6 95502522 N chr6 95503045 N DEL 15
SRR1766484.6430850 chr6 95502504 N chr6 95503162 N DUP 8
SRR1766463.4611848 chr6 95502629 N chr6 95503099 N DEL 24
SRR1766450.10426355 chr6 95502562 N chr6 95503099 N DEL 14
SRR1766450.98598 chr6 95502562 N chr6 95503099 N DEL 14
SRR1766464.9675500 chr6 95502629 N chr6 95503099 N DEL 21
SRR1766468.5301496 chr6 95502629 N chr6 95503099 N DEL 21
SRR1766449.4949800 chr6 95502629 N chr6 95503099 N DEL 21
SRR1766454.9052230 chr6 95502629 N chr6 95503099 N DEL 21
SRR1766473.8081173 chr6 95502536 N chr6 95503107 N DEL 7
SRR1766467.8252274 chr6 95502602 N chr6 95503237 N DUP 3
SRR1766486.4975504 chr6 95502569 N chr6 95503129 N DEL 7
SRR1766443.8918103 chr6 95503164 N chr6 95503230 N DUP 21
SRR1766451.8225970 chr6 95502531 N chr6 95503132 N DEL 10
SRR1766477.1828385 chr6 95503106 N chr6 95503175 N DUP 7
SRR1766472.6222309 chr6 95502538 N chr6 95503132 N DEL 5
SRR1766442.7162371 chr6 95503164 N chr6 95503230 N DUP 26
SRR1766477.10290181 chr6 95502629 N chr6 95503099 N DEL 25
SRR1766464.6484272 chr6 95502534 N chr6 95503135 N DEL 7
SRR1766483.10054416 chr6 95503164 N chr6 95503267 N DUP 25
SRR1766483.8520803 chr6 95502603 N chr6 95503268 N DUP 11
SRR1766475.7525721 chr6 95502621 N chr6 95503147 N DEL 9
SRR1766471.1031726 chr6 95502603 N chr6 95503268 N DUP 8
SRR1766469.6912328 chr6 95502603 N chr6 95503268 N DUP 9
SRR1766470.7324205 chr6 95502622 N chr6 95503148 N DEL 9
SRR1766474.3642564 chr6 95502603 N chr6 95503268 N DUP 10
SRR1766459.2158058 chr6 95502537 N chr6 95503173 N DEL 6
SRR1766451.5596099 chr6 95502538 N chr6 95503174 N DEL 5
SRR1766443.4658238 chr6 95502532 N chr6 95503205 N DEL 11
SRR1766463.5637768 chr6 95502614 N chr6 95503214 N DEL 2
SRR1766481.10835673 chr6 95502614 N chr6 95503214 N DEL 2
SRR1766478.5601427 chr6 95502533 N chr6 95503243 N DEL 10
SRR1766478.7658322 chr6 95502534 N chr6 95503244 N DEL 9
SRR1766485.11254779 chr6 95502536 N chr6 95503246 N DEL 7
SRR1766456.2893237 chr15 28371637 N chr15 28371691 N DEL 4
SRR1766452.1068694 chr1 109654236 N chr1 109654340 N DEL 10
SRR1766464.9546549 chr1 109654236 N chr1 109654340 N DEL 10
SRR1766481.1909562 chr1 109654236 N chr1 109654340 N DEL 10
SRR1766467.2741961 chr1 109654236 N chr1 109654340 N DEL 18
SRR1766483.5445389 chr1 109654307 N chr1 109654383 N DEL 7
SRR1766481.797284 chr1 109654236 N chr1 109654340 N DEL 7
SRR1766446.405548 chr1 109654253 N chr1 109654378 N DEL 4
SRR1766479.8252656 chr1 109654254 N chr1 109654379 N DEL 3
SRR1766448.2381653 chr5 181437379 N chr5 181437446 N DUP 5
SRR1766482.26435 chr5 181437394 N chr5 181437597 N DUP 5
SRR1766462.2076577 chr5 181437394 N chr5 181437529 N DUP 5
SRR1766442.15867481 chr5 181437461 N chr5 181437598 N DEL 5
SRR1766447.3866896 chr5 181437420 N chr5 181437555 N DUP 5
SRR1766462.1217967 chr3 9639315 N chr3 9639364 N DUP 13
SRR1766471.1235813 chr3 9639281 N chr3 9639334 N DEL 2
SRR1766442.47143513 chr7 60919983 N chr7 60920129 N DUP 5
SRR1766479.3973489 chr7 60920027 N chr7 60920320 N DUP 5
SRR1766442.1060365 chr7 60919991 N chr7 60920137 N DUP 5
SRR1766475.6671660 chr7 60919976 N chr7 60920122 N DUP 1
SRR1766476.6111175 chr7 60919991 N chr7 60920137 N DUP 10
SRR1766468.4353498 chr7 60919976 N chr7 60920122 N DUP 10
SRR1766442.27133974 chr7 60920011 N chr7 60920157 N DUP 5
SRR1766455.9808171 chr7 60919991 N chr7 60920137 N DUP 15
SRR1766478.11977666 chr7 60920011 N chr7 60920157 N DUP 5
SRR1766479.6682525 chr7 60920030 N chr7 60920178 N DEL 5
SRR1766448.2413914 chr15 63547907 N chr15 63548006 N DUP 11
SRR1766465.3421185 chr15 63547920 N chr15 63548015 N DUP 6
SRR1766444.666408 chr15 63547886 N chr15 63547979 N DEL 2
SRR1766468.3452328 chr15 63547953 N chr15 63548038 N DEL 15
SRR1766475.6928772 chr15 63547953 N chr15 63548038 N DEL 15
SRR1766461.1328256 chr15 63547956 N chr15 63548041 N DEL 12
SRR1766458.5317367 chr1 24907798 N chr1 24908349 N DEL 5
SRR1766452.9406567 chr1 24907858 N chr1 24908259 N DEL 4
SRR1766442.35488036 chr1 24907789 N chr1 24907863 N DUP 5
SRR1766470.7748660 chr1 24907789 N chr1 24907863 N DUP 12
SRR1766468.2921351 chr1 24907863 N chr1 24907964 N DEL 9
SRR1766442.28055915 chr1 24907838 N chr1 24908214 N DEL 46
SRR1766462.9549874 chr1 24907853 N chr1 24907904 N DEL 19
SRR1766449.25683 chr1 24907798 N chr1 24907847 N DUP 15
SRR1766463.6255815 chr1 24907772 N chr1 24907896 N DUP 5
SRR1766461.6646043 chr1 24907814 N chr1 24907888 N DUP 10
SRR1766442.37972525 chr1 24907797 N chr1 24907896 N DUP 5
SRR1766473.8145816 chr1 24907838 N chr1 24907964 N DEL 5
SRR1766448.4688978 chr1 24907883 N chr1 24908259 N DEL 15
SRR1766442.13855244 chr1 24907846 N chr1 24907897 N DEL 5
SRR1766463.5124091 chr1 24907779 N chr1 24907928 N DUP 4
SRR1766476.4593966 chr1 24907958 N chr1 24908384 N DEL 17
SRR1766445.1939040 chr1 24907914 N chr1 24907963 N DUP 3
SRR1766446.1414159 chr1 24907814 N chr1 24907963 N DUP 5
SRR1766464.1279360 chr1 24907843 N chr1 24907894 N DEL 5
SRR1766457.5101521 chr1 24907814 N chr1 24907988 N DUP 3
SRR1766474.6169101 chr1 24907964 N chr1 24908440 N DEL 5
SRR1766485.3604234 chr1 24907769 N chr1 24907993 N DUP 5
SRR1766442.28107993 chr1 24907797 N chr1 24907923 N DEL 5
SRR1766465.7677414 chr1 24907797 N chr1 24908021 N DUP 5
SRR1766475.2026128 chr1 24907778 N chr1 24908002 N DUP 5
SRR1766447.1626678 chr1 24907797 N chr1 24908021 N DUP 5
SRR1766442.24885332 chr1 24907864 N chr1 24907988 N DUP 2
SRR1766463.9151774 chr1 24907839 N chr1 24908013 N DUP 10
SRR1766471.10855959 chr1 24908063 N chr1 24908139 N DEL 10
SRR1766475.5398998 chr1 24907940 N chr1 24908016 N DEL 5
SRR1766459.7712357 chr1 24907789 N chr1 24908113 N DUP 5
SRR1766460.10188705 chr1 24908133 N chr1 24908259 N DEL 2
SRR1766461.1487471 chr1 24907797 N chr1 24908071 N DUP 15
SRR1766444.3779310 chr1 24907789 N chr1 24908138 N DUP 5
SRR1766442.16443552 chr1 24907789 N chr1 24908138 N DUP 5
SRR1766485.10646826 chr1 24907789 N chr1 24908138 N DUP 5
SRR1766464.5546754 chr1 24908123 N chr1 24908224 N DEL 10
SRR1766477.191771 chr1 24908158 N chr1 24908259 N DEL 2
SRR1766442.45998972 chr1 24908113 N chr1 24908214 N DEL 12
SRR1766442.33929118 chr1 24908098 N chr1 24908172 N DUP 5
SRR1766478.1764817 chr1 24907789 N chr1 24908138 N DUP 5
SRR1766484.10456616 chr1 24907790 N chr1 24908066 N DEL 5
SRR1766486.2662318 chr1 24907883 N chr1 24908334 N DEL 29
SRR1766450.9369944 chr1 24907883 N chr1 24908384 N DEL 24
SRR1766452.8642710 chr1 24907830 N chr1 24908106 N DEL 8
SRR1766462.7209640 chr1 24908198 N chr1 24908449 N DEL 5
SRR1766479.9220674 chr1 24908123 N chr1 24908172 N DUP 11
SRR1766484.8920565 chr1 24907977 N chr1 24908128 N DEL 1
SRR1766449.10873285 chr1 24907958 N chr1 24908184 N DEL 15
SRR1766442.29140521 chr1 24907783 N chr1 24908184 N DEL 15
SRR1766442.35488036 chr1 24908123 N chr1 24908172 N DUP 5
SRR1766456.2379281 chr1 24908214 N chr1 24908263 N DUP 10
SRR1766442.28055915 chr1 24908214 N chr1 24908263 N DUP 15
SRR1766446.1414159 chr1 24908285 N chr1 24908336 N DEL 9
SRR1766477.5304532 chr1 24908214 N chr1 24908263 N DUP 15
SRR1766452.9406567 chr1 24908214 N chr1 24908263 N DUP 10
SRR1766485.3604234 chr1 24908282 N chr1 24908333 N DEL 10
SRR1766447.6754007 chr1 24908199 N chr1 24908273 N DUP 10
SRR1766478.5748053 chr1 24907807 N chr1 24908258 N DEL 5
SRR1766464.7141671 chr1 24908214 N chr1 24908263 N DUP 14
SRR1766469.4339725 chr1 24908251 N chr1 24908327 N DEL 15
SRR1766475.2712178 chr1 24908282 N chr1 24908333 N DEL 15
SRR1766477.6135919 chr1 24908208 N chr1 24908284 N DEL 10
SRR1766484.1858938 chr1 24908208 N chr1 24908284 N DEL 10
SRR1766442.24885332 chr1 24908282 N chr1 24908333 N DEL 11
SRR1766483.4939124 chr1 24908251 N chr1 24908327 N DEL 5
SRR1766444.3894676 chr1 24908251 N chr1 24908327 N DEL 5
SRR1766443.6686168 chr1 24908251 N chr1 24908327 N DEL 5
SRR1766465.7020159 chr1 24908267 N chr1 24908343 N DEL 5
SRR1766448.4688978 chr1 24908251 N chr1 24908327 N DEL 5
SRR1766479.13071233 chr1 24908273 N chr1 24908349 N DEL 10
SRR1766478.8958767 chr1 24908212 N chr1 24908338 N DEL 5
SRR1766482.7191304 chr1 24907807 N chr1 24908333 N DEL 9
SRR1766457.5101521 chr1 24908258 N chr1 24908359 N DEL 5
SRR1766464.5546754 chr1 24908288 N chr1 24908339 N DEL 8
SRR1766451.8353345 chr1 24908294 N chr1 24908345 N DEL 3
SRR1766457.5759551 chr1 24907808 N chr1 24908359 N DEL 10
SRR1766460.115271 chr1 24907883 N chr1 24908409 N DEL 26
SRR1766471.10855959 chr1 24907858 N chr1 24908409 N DEL 25
SRR1766477.1740154 chr1 24907864 N chr1 24908440 N DEL 10
SRR1766470.7748660 chr1 24907864 N chr1 24908440 N DEL 20
SRR1766445.7170298 chr1 24907819 N chr1 24908420 N DEL 4
SRR1766449.6903238 chr1 24907820 N chr1 24908421 N DEL 3
SRR1766450.3484013 chr1 24908266 N chr1 24908442 N DEL 5
SRR1766460.10188705 chr1 24908241 N chr1 24908442 N DEL 10
SRR1766456.2379281 chr1 24907803 N chr1 24908454 N DEL 1
SRR1766443.3928177 chr9 80740993 N chr9 80741074 N DEL 4
SRR1766442.26659058 chr9 80741006 N chr9 80741070 N DEL 3
SRR1766485.4198702 chr9 80740993 N chr9 80741074 N DEL 3
SRR1766469.543586 chr9 80741011 N chr9 80741073 N DEL 6
SRR1766449.9247023 chr7 205394 N chr7 205485 N DUP 5
SRR1766445.9655537 chr7 205405 N chr7 205496 N DUP 14
SRR1766476.2639533 chr7 205405 N chr7 205496 N DUP 27
SRR1766466.11305139 chr7 205394 N chr7 205485 N DUP 22
SRR1766483.9406399 chr7 205408 N chr7 205499 N DUP 6
SRR1766447.6251263 chr7 205394 N chr7 205485 N DUP 27
SRR1766482.7684917 chr2 202215769 N chr2 202216113 N DEL 5
SRR1766442.21365535 chr2 202215769 N chr2 202216113 N DEL 5
SRR1766449.5296168 chr2 202215769 N chr2 202216113 N DEL 5
SRR1766447.1871558 chr2 202215769 N chr2 202216113 N DEL 5
SRR1766481.3136639 chr2 202215769 N chr2 202216113 N DEL 5
SRR1766458.8365830 chr2 202215769 N chr2 202216113 N DEL 5
SRR1766446.3980025 chr2 202215769 N chr2 202216113 N DEL 5
SRR1766466.10469718 chr1 125179251 N chr1 125179397 N DUP 5
SRR1766445.929483 chr1 125179329 N chr1 125179449 N DUP 2
SRR1766444.4740112 chr1 125179395 N chr1 125179492 N DUP 3
SRR1766478.4488520 chr1 125179352 N chr1 125179428 N DEL 20
SRR1766451.5194082 chr1 125179352 N chr1 125179428 N DEL 12
SRR1766470.6503590 chr1 125179251 N chr1 125179469 N DUP 2
SRR1766459.4039858 chr1 125179296 N chr1 125179465 N DUP 5
SRR1766466.4273055 chr1 125179358 N chr1 125179434 N DEL 5
SRR1766481.10385244 chr1 125179351 N chr1 125179404 N DEL 57
SRR1766445.6516164 chr1 125179352 N chr1 125179428 N DEL 32
SRR1766442.33367673 chr1 125179358 N chr1 125179434 N DEL 10
SRR1766486.2919519 chr1 125179293 N chr1 125179413 N DUP 5
SRR1766467.2287342 chr1 125179358 N chr1 125179434 N DEL 23
SRR1766454.10731734 chr1 125179309 N chr1 125179431 N DEL 5
SRR1766444.2249590 chr9 80232120 N chr9 80232234 N DEL 29
SRR1766482.9769953 chr17 44590233 N chr17 44591084 N DEL 5
SRR1766450.8761951 chr17 44590290 N chr17 44590385 N DEL 5
SRR1766459.8859478 chr17 44590321 N chr17 44590820 N DEL 5
SRR1766454.578896 chr17 44590321 N chr17 44590820 N DEL 5
SRR1766442.35238573 chr17 44590324 N chr17 44590761 N DEL 6
SRR1766468.1723132 chr17 44590290 N chr17 44590385 N DEL 5
SRR1766479.8177296 chr17 44590321 N chr17 44590820 N DEL 5
SRR1766482.11466502 chr17 44590291 N chr17 44590384 N DUP 4
SRR1766469.2496600 chr17 44590386 N chr17 44591083 N DEL 10
SRR1766464.9138537 chr17 44590415 N chr17 44590930 N DEL 10
SRR1766479.3020842 chr17 44590349 N chr17 44591074 N DUP 5
SRR1766462.4211385 chr17 44590248 N chr17 44590343 N DEL 1
SRR1766449.3016692 chr17 44590271 N chr17 44590366 N DEL 5
SRR1766463.7386450 chr17 44590388 N chr17 44590543 N DUP 1
SRR1766485.8032887 chr17 44590412 N chr17 44591203 N DUP 5
SRR1766451.2180247 chr17 44590193 N chr17 44590532 N DUP 1
SRR1766482.6468820 chr17 44590539 N chr17 44590930 N DEL 5
SRR1766483.3552551 chr17 44590539 N chr17 44590930 N DEL 5
SRR1766462.9241409 chr17 44590489 N chr17 44590548 N DUP 9
SRR1766443.7114113 chr17 44590539 N chr17 44590930 N DEL 5
SRR1766484.2797225 chr17 44590240 N chr17 44590551 N DUP 5
SRR1766462.4873983 chr17 44590539 N chr17 44590930 N DEL 5
SRR1766446.3778975 chr17 44590492 N chr17 44590551 N DUP 1
SRR1766445.2617548 chr17 44590583 N chr17 44591092 N DEL 8
SRR1766454.1684115 chr17 44590385 N chr17 44590606 N DUP 15
SRR1766477.2070612 chr17 44590252 N chr17 44590565 N DEL 3
SRR1766485.7384872 chr17 44590242 N chr17 44590677 N DUP 1
SRR1766483.10037354 chr17 44590677 N chr17 44591092 N DEL 10
SRR1766445.3499027 chr17 44590620 N chr17 44591127 N DUP 14
SRR1766450.5753278 chr17 44590689 N chr17 44591104 N DEL 6
SRR1766448.439448 chr17 44590241 N chr17 44590740 N DUP 1
SRR1766450.10727211 chr17 44590395 N chr17 44590740 N DUP 3
SRR1766464.3403357 chr17 44590395 N chr17 44590740 N DUP 3
SRR1766486.55062 chr17 44590395 N chr17 44590740 N DUP 4
SRR1766442.15969032 chr17 44590395 N chr17 44590740 N DUP 12
SRR1766443.8243244 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766473.2822904 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766484.3240924 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766475.9173113 chr17 44590740 N chr17 44591091 N DEL 13
SRR1766463.6044678 chr17 44590740 N chr17 44591091 N DEL 13
SRR1766449.7492892 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766471.6130177 chr17 44590761 N chr17 44590930 N DEL 18
SRR1766442.10353299 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766475.5759455 chr17 44590253 N chr17 44590660 N DEL 3
SRR1766450.8761951 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766477.2407161 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766479.13315133 chr17 44590395 N chr17 44590740 N DUP 13
SRR1766455.947410 chr17 44590389 N chr17 44590734 N DUP 11
SRR1766485.9632066 chr17 44590306 N chr17 44590717 N DEL 8
SRR1766446.3261484 chr17 44590807 N chr17 44591100 N DEL 1
SRR1766455.8843831 chr17 44590443 N chr17 44590786 N DEL 8
SRR1766478.11726904 chr17 44590422 N chr17 44590765 N DEL 13
SRR1766455.7350953 chr17 44590337 N chr17 44590774 N DEL 6
SRR1766459.8859478 chr17 44590799 N chr17 44590860 N DUP 9
SRR1766442.24034544 chr17 44590254 N chr17 44590785 N DEL 5
SRR1766466.2844710 chr17 44590823 N chr17 44591022 N DUP 5
SRR1766483.3552551 chr17 44590512 N chr17 44590853 N DEL 2
SRR1766477.11942491 chr17 44590924 N chr17 44591001 N DUP 5
SRR1766483.10037354 chr17 44590408 N chr17 44591041 N DEL 8
SRR1766476.9104055 chr17 44590524 N chr17 44591125 N DUP 5
SRR1766483.2086671 chr17 44590408 N chr17 44591041 N DEL 6
SRR1766481.12704635 chr17 44590970 N chr17 44591055 N DEL 6
SRR1766443.8442555 chr17 44590816 N chr17 44591139 N DUP 5
SRR1766467.4290667 chr17 44590261 N chr17 44591048 N DEL 5
SRR1766471.213104 chr17 44590270 N chr17 44591057 N DEL 10
SRR1766455.8223330 chr17 44590422 N chr17 44591055 N DEL 1
SRR1766457.7947741 chr17 44590265 N chr17 44591052 N DEL 2
SRR1766478.4840639 chr17 44590484 N chr17 44591085 N DEL 4
SRR1766457.3267102 chr17 44591076 N chr17 44591201 N DUP 5
SRR1766471.6130177 chr17 44591076 N chr17 44591201 N DUP 5
SRR1766475.7695180 chr17 44591076 N chr17 44591201 N DUP 9
SRR1766454.1684115 chr17 44590262 N chr17 44591083 N DEL 5
SRR1766447.3709357 chr17 44590391 N chr17 44591114 N DEL 3
SRR1766478.4333706 chr17 44591106 N chr17 44591201 N DUP 5
SRR1766455.7350953 chr17 44590262 N chr17 44591147 N DEL 5
SRR1766479.8310289 chr17 44590249 N chr17 44591306 N DUP 2
SRR1766485.4094960 chr17 44590249 N chr17 44591306 N DUP 5
SRR1766465.4341180 chr17 44590305 N chr17 44591192 N DEL 4
SRR1766442.46023542 chr17 44590249 N chr17 44591306 N DUP 8
SRR1766463.3603547 chr17 44590249 N chr17 44591306 N DUP 9
SRR1766476.8203177 chr17 44591099 N chr17 44591306 N DUP 9
SRR1766445.8982419 chr17 44590808 N chr17 44591307 N DUP 9
SRR1766442.31747534 chr17 44590808 N chr17 44591307 N DUP 9
SRR1766445.9900784 chr17 44590808 N chr17 44591307 N DUP 9
SRR1766480.623884 chr17 44590808 N chr17 44591307 N DUP 9
SRR1766479.7322480 chr17 44590267 N chr17 44591230 N DEL 2
SRR1766463.4457992 chr17 44590808 N chr17 44591307 N DUP 9
SRR1766484.12105646 chr17 44590812 N chr17 44591311 N DUP 9
SRR1766457.8828096 chr17 44590274 N chr17 44591299 N DEL 5
SRR1766443.10678939 chr17 44590271 N chr17 44591328 N DEL 2
SRR1766450.1105841 chr16 88470628 N chr16 88470679 N DEL 10
SRR1766485.5672307 chr16 88470679 N chr16 88471028 N DUP 5
SRR1766442.217937 chr16 88470713 N chr16 88470914 N DEL 5
SRR1766469.10831011 chr16 88470714 N chr16 88470915 N DEL 5
SRR1766486.11340589 chr16 88470674 N chr16 88470925 N DEL 4
SRR1766461.9353432 chr9 37752584 N chr9 37752745 N DEL 1
SRR1766460.10825514 chr2 3170747 N chr2 3171169 N DEL 4
SRR1766464.9334641 chr2 3170747 N chr2 3171169 N DEL 4
SRR1766451.5444657 chr2 3170747 N chr2 3171169 N DEL 5
SRR1766464.1048660 chr2 3170747 N chr2 3171169 N DEL 6
SRR1766465.3958736 chr2 3170751 N chr2 3170808 N DUP 5
SRR1766470.5210468 chr2 3170850 N chr2 3171046 N DEL 5
SRR1766443.8514314 chr2 3170899 N chr2 3170954 N DUP 7
SRR1766447.10208748 chr2 3171063 N chr2 3171180 N DEL 23
SRR1766450.8204601 chr2 3170874 N chr2 3171014 N DEL 5
SRR1766458.5734426 chr2 3170772 N chr2 3171109 N DEL 1
SRR1766486.3159767 chr2 3171071 N chr2 3171241 N DUP 5
SRR1766465.6468038 chr2 3171071 N chr2 3171241 N DUP 5
SRR1766478.479485 chr2 3171190 N chr2 3171244 N DUP 6
SRR1766479.11691689 chr2 3171190 N chr2 3171244 N DUP 18
SRR1766479.11281910 chr2 3171196 N chr2 3171250 N DUP 8
SRR1766451.4716138 chr2 3171196 N chr2 3171250 N DUP 8
SRR1766466.10352372 chr2 3171086 N chr2 3171203 N DEL 2
SRR1766460.3353206 chr2 3170821 N chr2 3171216 N DEL 10
SRR1766481.9609543 chr11 134759990 N chr11 134760197 N DUP 15
SRR1766462.8992315 chr11 134760064 N chr11 134760197 N DUP 24
SRR1766463.7812259 chr11 134760031 N chr11 134760178 N DUP 5
SRR1766443.5917413 chr11 134760031 N chr11 134760104 N DUP 18
SRR1766463.3743914 chr11 134760031 N chr11 134760178 N DUP 5
SRR1766456.3078444 chr11 134760031 N chr11 134760104 N DUP 15
SRR1766457.6354110 chr11 134760031 N chr11 134760178 N DUP 5
SRR1766466.10149980 chr11 134760067 N chr11 134760200 N DUP 24
SRR1766466.4152538 chr11 134760031 N chr11 134760104 N DUP 14
SRR1766467.3018696 chr11 134760067 N chr11 134760200 N DUP 24
SRR1766442.21274371 chr11 134760031 N chr11 134760178 N DUP 5
SRR1766478.4044906 chr11 134760031 N chr11 134760178 N DUP 5
SRR1766459.10183360 chr11 134760033 N chr11 134760106 N DUP 7
SRR1766443.9572108 chr11 134760034 N chr11 134760107 N DUP 6
SRR1766483.3873771 chr11 134760031 N chr11 134760104 N DUP 10
SRR1766485.517087 chr11 134760040 N chr11 134760395 N DUP 10
SRR1766474.7113443 chr11 134760041 N chr11 134760114 N DUP 5
SRR1766485.8543405 chr11 134760042 N chr11 134760115 N DUP 4
SRR1766472.11564031 chr11 134760042 N chr11 134760397 N DUP 9
SRR1766442.11731002 chr11 134760045 N chr11 134760118 N DUP 1
SRR1766455.3245018 chr11 134760071 N chr11 134760278 N DUP 5
SRR1766455.6454893 chr11 134760061 N chr11 134760268 N DUP 7
SRR1766458.4850667 chr11 134760054 N chr11 134760261 N DUP 1
SRR1766442.7435638 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766482.6260456 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766474.9422298 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766457.7477206 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766442.2689425 chr11 134760069 N chr11 134760276 N DUP 5
SRR1766443.35058 chr11 134760069 N chr11 134760276 N DUP 10
SRR1766461.8531692 chr11 134760069 N chr11 134760276 N DUP 7
SRR1766443.10428085 chr11 134760094 N chr11 134760301 N DUP 16
SRR1766483.8493958 chr11 134760069 N chr11 134760276 N DUP 6
SRR1766463.3696355 chr11 134760075 N chr11 134760208 N DUP 4
SRR1766446.10520792 chr11 134759990 N chr11 134760197 N DUP 8
SRR1766462.1531734 chr11 134760143 N chr11 134760202 N DUP 11
SRR1766459.1477109 chr11 134760211 N chr11 134760360 N DEL 1
SRR1766456.3047089 chr11 134759990 N chr11 134760197 N DUP 31
SRR1766474.6168090 chr11 134760117 N chr11 134760190 N DUP 4
SRR1766474.3903465 chr11 134760118 N chr11 134760191 N DUP 3
SRR1766482.887027 chr11 134760119 N chr11 134760192 N DUP 2
SRR1766446.9018027 chr11 134760211 N chr11 134760286 N DEL 15
SRR1766447.10436602 chr11 134760143 N chr11 134760202 N DUP 11
SRR1766442.10088735 chr11 134760143 N chr11 134760202 N DUP 18
SRR1766465.10897309 chr11 134760143 N chr11 134760202 N DUP 20
SRR1766475.6873438 chr11 134760144 N chr11 134760351 N DUP 10
SRR1766467.3838176 chr11 134760143 N chr11 134760202 N DUP 37
SRR1766478.6104799 chr11 134760113 N chr11 134760188 N DEL 4
SRR1766456.3047089 chr11 134760004 N chr11 134760285 N DUP 14
SRR1766483.458014 chr11 134760240 N chr11 134760313 N DUP 5
SRR1766468.7882697 chr11 134760104 N chr11 134760239 N DEL 10
SRR1766454.5165818 chr11 134760239 N chr11 134760386 N DUP 5
SRR1766465.4675722 chr11 134760239 N chr11 134760386 N DUP 5
SRR1766469.7363042 chr11 134760239 N chr11 134760386 N DUP 5
SRR1766444.1231017 chr11 134760239 N chr11 134760386 N DUP 5
SRR1766453.7656884 chr11 134760239 N chr11 134760386 N DUP 5
SRR1766442.15336647 chr11 134760239 N chr11 134760386 N DUP 5
SRR1766460.10223199 chr11 134760239 N chr11 134760386 N DUP 5
SRR1766472.11752423 chr11 134760239 N chr11 134760386 N DUP 5
SRR1766471.10661128 chr11 134760063 N chr11 134760344 N DUP 3
SRR1766473.10258808 chr11 134760063 N chr11 134760344 N DUP 6
SRR1766451.5231405 chr11 134760063 N chr11 134760344 N DUP 7
SRR1766462.5882867 chr11 134760063 N chr11 134760344 N DUP 10
SRR1766456.737250 chr3 197518859 N chr3 197519217 N DEL 2
SRR1766450.8769198 chr3 197518828 N chr3 197519239 N DEL 5
SRR1766478.4310245 chr3 197518840 N chr3 197519251 N DEL 28
SRR1766454.2434953 chr3 197519106 N chr3 197519245 N DEL 5
SRR1766445.8997835 chr1 241713498 N chr1 241713566 N DEL 14
SRR1766486.1390320 chr20 38284610 N chr20 38284916 N DEL 6
SRR1766481.2768284 chr1 22227678 N chr1 22227733 N DUP 16
SRR1766481.723426 chr11 105491340 N chr11 105491393 N DEL 9
SRR1766472.7448157 chr22 18418040 N chr22 18418094 N DEL 1
SRR1766457.1937608 chr22 18418066 N chr22 18418235 N DEL 9
SRR1766469.9191209 chr22 18418066 N chr22 18418235 N DEL 13
SRR1766466.9481213 chr22 18418066 N chr22 18418235 N DEL 15
SRR1766442.23128855 chr22 18418152 N chr22 18418273 N DUP 28
SRR1766448.5933464 chr22 18418152 N chr22 18418273 N DUP 27
SRR1766450.1178376 chr22 18418212 N chr22 18418294 N DUP 17
SRR1766472.9672541 chr22 18418214 N chr22 18418326 N DUP 20
SRR1766465.3728799 chr22 18418189 N chr22 18418266 N DUP 39
SRR1766465.4943142 chr22 18418212 N chr22 18418294 N DUP 18
SRR1766464.5510248 chr22 18418189 N chr22 18418266 N DUP 32
SRR1766485.10781574 chr22 18418212 N chr22 18418294 N DUP 19
SRR1766462.8834263 chr22 18418127 N chr22 18418260 N DUP 2
SRR1766471.11937713 chr22 18418189 N chr22 18418266 N DUP 32
SRR1766477.3328323 chr22 18418212 N chr22 18418294 N DUP 17
SRR1766447.7280118 chr22 18418189 N chr22 18418266 N DUP 26
SRR1766442.37538566 chr22 18418189 N chr22 18418266 N DUP 26
SRR1766476.9848852 chr22 18418189 N chr22 18418266 N DUP 21
SRR1766466.6327549 chr22 18418189 N chr22 18418266 N DUP 26
SRR1766458.9247823 chr22 18418189 N chr22 18418266 N DUP 22
SRR1766442.11164701 chr22 18418189 N chr22 18418266 N DUP 27
SRR1766465.5426755 chr22 18418189 N chr22 18418266 N DUP 15
SRR1766470.5908973 chr22 18418152 N chr22 18418273 N DUP 25
SRR1766449.8824936 chr22 18418145 N chr22 18418209 N DEL 14
SRR1766459.10890299 chr22 18418060 N chr22 18418211 N DEL 10
SRR1766471.1389166 chr22 18418086 N chr22 18418214 N DEL 9
SRR1766484.3202362 chr22 18418059 N chr22 18418217 N DEL 6
SRR1766455.8370433 chr22 18418153 N chr22 18418251 N DEL 7
SRR1766459.9571510 chr22 18418143 N chr22 18418391 N DUP 10
SRR1766442.17251044 chr22 18418145 N chr22 18418280 N DEL 5
SRR1766442.3053089 chr22 18418145 N chr22 18418280 N DEL 5
SRR1766481.3639483 chr22 18418392 N chr22 18418611 N DUP 8
SRR1766442.22207367 chr22 18418140 N chr22 18418410 N DEL 19
SRR1766476.5808589 chr22 18418140 N chr22 18418410 N DEL 19
SRR1766452.6905395 chr22 18418228 N chr22 18418418 N DEL 7
SRR1766457.4857609 chr22 18418144 N chr22 18418416 N DEL 10
SRR1766484.2964924 chr22 18418208 N chr22 18418658 N DUP 7
SRR1766446.6669165 chr22 18417990 N chr22 18418587 N DEL 5
SRR1766461.8860696 chr22 18418058 N chr22 18418588 N DEL 5
SRR1766475.499825 chr22 18418243 N chr22 18418711 N DUP 2
SRR1766442.11542737 chr22 18418547 N chr22 18418729 N DUP 11
SRR1766478.10964601 chr22 18418547 N chr22 18418729 N DUP 14
SRR1766460.758014 chr1 225833945 N chr1 225834247 N DUP 5
SRR1766468.3139261 chr1 225833959 N chr1 225834264 N DEL 5
SRR1766483.6169853 chr1 225833959 N chr1 225834268 N DEL 5
SRR1766465.9486362 chr1 225833959 N chr1 225834272 N DEL 5
SRR1766442.44751700 chr1 225833959 N chr1 225834275 N DEL 2
SRR1766442.30975724 chr1 225834055 N chr1 225834365 N DEL 5
SRR1766442.31499190 chr1 225833808 N chr1 225834419 N DEL 12
SRR1766442.4852873 chr1 225834117 N chr1 225834425 N DEL 5
SRR1766482.1056390 chr1 225834129 N chr1 225834437 N DEL 7
SRR1766486.7534306 chr11 73935624 N chr11 73935750 N DUP 8
SRR1766442.2578512 chr18 2222995 N chr18 2223048 N DEL 57
SRR1766483.6667452 chr2 108937648 N chr2 108937836 N DEL 6
SRR1766485.3985534 chr18 59233821 N chr18 59234102 N DEL 7
SRR1766474.8333605 chr18 59233821 N chr18 59234102 N DEL 8
SRR1766452.1750196 chr18 59233861 N chr18 59234146 N DEL 3
SRR1766459.9796378 chr18 59233861 N chr18 59234146 N DEL 5
SRR1766461.6452719 chr18 59233861 N chr18 59234146 N DEL 6
SRR1766472.2942756 chr18 59233868 N chr18 59233988 N DEL 8
SRR1766471.9015319 chr18 59233864 N chr18 59234137 N DEL 6
SRR1766479.295951 chr18 59233868 N chr18 59233988 N DEL 12
SRR1766483.3881660 chr18 59233868 N chr18 59233988 N DEL 12
SRR1766478.8731711 chr18 59233835 N chr18 59233932 N DUP 11
SRR1766475.9609132 chr18 59233810 N chr18 59233931 N DUP 15
SRR1766446.3165791 chr18 59233835 N chr18 59233932 N DUP 13
SRR1766443.729958 chr18 59233850 N chr18 59233913 N DEL 7
SRR1766463.259549 chr18 59233851 N chr18 59233900 N DUP 25
SRR1766442.45297134 chr18 59233810 N chr18 59233931 N DUP 22
SRR1766466.3317853 chr18 59233852 N chr18 59233901 N DUP 14
SRR1766442.9341603 chr18 59233751 N chr18 59234005 N DUP 14
SRR1766461.10760957 chr18 59233823 N chr18 59234088 N DUP 12
SRR1766442.22999578 chr18 59234185 N chr18 59234258 N DEL 1
SRR1766458.5704118 chr18 59234185 N chr18 59234258 N DEL 11
SRR1766448.6989772 chr18 59234185 N chr18 59234258 N DEL 13
SRR1766461.10703115 chr18 59234185 N chr18 59234258 N DEL 24
SRR1766469.7383809 chr18 59234187 N chr18 59234260 N DEL 10
SRR1766472.5458148 chr18 59234185 N chr18 59234258 N DEL 20
SRR1766481.1496601 chr18 59234187 N chr18 59234260 N DEL 10
SRR1766454.1764960 chr9 35460529 N chr9 35460617 N DUP 5
SRR1766448.2097785 chr9 35460531 N chr9 35460619 N DUP 3
SRR1766457.3040827 chr1 55664221 N chr1 55664478 N DUP 4
SRR1766481.7195825 chr1 55664307 N chr1 55664540 N DUP 6
SRR1766472.7285134 chr1 55664570 N chr1 55664624 N DEL 5
SRR1766469.7717429 chr1 188210807 N chr1 188210903 N DEL 2
SRR1766442.23626244 chr1 188210807 N chr1 188210907 N DEL 3
SRR1766481.804726 chr1 188210807 N chr1 188210907 N DEL 4
SRR1766468.1096737 chr1 188210807 N chr1 188210907 N DEL 8
SRR1766442.20799439 chr1 188210807 N chr1 188210907 N DEL 9
SRR1766474.1320832 chr1 188210856 N chr1 188210909 N DUP 9
SRR1766467.4865326 chr10 69792040 N chr10 69792132 N DUP 5
SRR1766470.7982521 chrX 140768792 N chrX 140768849 N DEL 12
SRR1766481.10174862 chrX 140768792 N chrX 140768849 N DEL 13
SRR1766442.43291554 chr8 18489112 N chr8 18489248 N DUP 1
SRR1766445.3644902 chr8 18489241 N chr8 18489302 N DUP 3
SRR1766467.10878909 chr8 18489081 N chr8 18489304 N DEL 3
SRR1766442.20578156 chr12 5928554 N chr12 5928618 N DEL 13
SRR1766442.20617090 chr12 5928554 N chr12 5928618 N DEL 13
SRR1766442.25710574 chr12 5928554 N chr12 5928618 N DEL 13
SRR1766452.7158607 chr12 5928554 N chr12 5928618 N DEL 18
SRR1766457.8394693 chr12 5928691 N chr12 5929724 N DEL 8
SRR1766468.5479529 chr12 5928691 N chr12 5929724 N DEL 10
SRR1766461.10704418 chr12 5928691 N chr12 5929724 N DEL 15
SRR1766470.6906476 chr12 5928691 N chr12 5929724 N DEL 15
SRR1766442.35696168 chr12 5928691 N chr12 5929724 N DEL 15
SRR1766467.1280076 chr12 5928691 N chr12 5929724 N DEL 15
SRR1766476.10023263 chr12 5928755 N chr12 5929327 N DEL 5
SRR1766472.2551058 chr12 5928755 N chr12 5929327 N DEL 5
SRR1766446.3027580 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766459.2811676 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766477.9709290 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766449.9216613 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766471.12207763 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766452.6820522 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766469.4702599 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766446.7427157 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766459.898553 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766446.10526081 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766459.3715909 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766477.10938337 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766481.7981316 chr12 5928687 N chr12 5929792 N DUP 6
SRR1766460.7652011 chr12 5928899 N chr12 5929782 N DUP 7
SRR1766467.2562635 chr12 5928687 N chr12 5929792 N DUP 7
SRR1766467.11511842 chr12 5928673 N chr12 5929338 N DUP 5
SRR1766470.6387460 chr12 5928899 N chr12 5929782 N DUP 7
SRR1766476.8843704 chr12 5928899 N chr12 5929782 N DUP 7
SRR1766445.2056253 chr12 5928678 N chr12 5928901 N DEL 5
SRR1766469.3814881 chr12 5929797 N chr12 5929868 N DEL 10
SRR1766463.3562469 chr12 5928687 N chr12 5929792 N DUP 5
SRR1766475.4266602 chr12 5929797 N chr12 5929868 N DEL 10
SRR1766482.550243 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766456.4130722 chr12 5928687 N chr12 5928739 N DUP 5
SRR1766479.11403056 chr12 5928691 N chr12 5928743 N DUP 5
SRR1766471.34104 chr12 5928692 N chr12 5928744 N DUP 5
SRR1766476.7888934 chr12 5928693 N chr12 5929337 N DUP 5
SRR1766454.5418474 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766484.1866593 chr12 5928696 N chr12 5929340 N DUP 5
SRR1766472.7202458 chr12 5928696 N chr12 5929340 N DUP 5
SRR1766467.11511842 chr12 5929341 N chr12 5929729 N DEL 7
SRR1766470.1420152 chr12 5928765 N chr12 5929428 N DEL 4
SRR1766475.5056492 chr12 5928663 N chr12 5928810 N DUP 10
SRR1766482.3930703 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766442.34141561 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766443.6187103 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766453.1126053 chr12 5928744 N chr12 5929263 N DEL 10
SRR1766485.7276342 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766470.6387460 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766486.11566260 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766477.4216808 chr12 5929337 N chr12 5929630 N DEL 9
SRR1766467.8152235 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766470.3645154 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766470.3952904 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766456.2132819 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766463.1491058 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766458.2751128 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766477.4216808 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766478.1657900 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766464.8127649 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766477.4271506 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766470.3952904 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766450.6808582 chr12 5928688 N chr12 5928909 N DUP 1
SRR1766469.10298811 chr12 5928775 N chr12 5929804 N DEL 5
SRR1766442.29850140 chr12 5928746 N chr12 5929703 N DUP 5
SRR1766484.809816 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766446.6596242 chr12 5928746 N chr12 5929703 N DUP 5
SRR1766442.13385760 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766472.8895753 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766475.536178 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766444.5430644 chr12 5928820 N chr12 5929337 N DUP 5
SRR1766469.6666315 chr12 5928777 N chr12 5929222 N DEL 1
SRR1766482.7241224 chr12 5928777 N chr12 5929222 N DEL 1
SRR1766486.2556641 chr12 5928777 N chr12 5929222 N DEL 3
SRR1766459.3614255 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766449.907380 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766442.38968041 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766479.4768605 chr12 5928663 N chr12 5928810 N DUP 5
SRR1766442.16581484 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766475.961206 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766464.2967461 chr12 5928663 N chr12 5929328 N DUP 8
SRR1766484.7848537 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766442.40349687 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766469.10298811 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766457.309465 chr12 5928672 N chr12 5928745 N DUP 5
SRR1766458.2911336 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766460.8653614 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766482.3930703 chr12 5928894 N chr12 5929337 N DUP 10
SRR1766456.2132819 chr12 5929511 N chr12 5929804 N DEL 15
SRR1766462.8068802 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766447.6487537 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766463.1491058 chr12 5928923 N chr12 5929804 N DEL 5
SRR1766450.8794248 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766465.2393348 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766481.424250 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766481.6765539 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766471.3674475 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766481.7697176 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766484.9151315 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766474.7186199 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766442.13385760 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766455.9250164 chr12 5928894 N chr12 5929337 N DUP 10
SRR1766463.3562469 chr12 5929804 N chr12 5929877 N DUP 10
SRR1766459.4505908 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766473.3316822 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766446.6596242 chr12 5928894 N chr12 5929337 N DUP 10
SRR1766453.11133758 chr12 5928663 N chr12 5929472 N DUP 5
SRR1766481.8082011 chr12 5928967 N chr12 5930144 N DEL 6
SRR1766469.2484114 chr12 5928764 N chr12 5930089 N DEL 3
SRR1766482.6561632 chr12 5928663 N chr12 5928958 N DUP 10
SRR1766442.16581484 chr12 5928893 N chr12 5928966 N DUP 5
SRR1766463.2108008 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766442.34598884 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766452.2226149 chr12 5928754 N chr12 5930153 N DEL 5
SRR1766481.7981316 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766476.7888934 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766446.1555345 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766474.10714393 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766442.1020869 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766463.5892525 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766443.8598106 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766446.3027580 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766457.8394693 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766459.3715909 chr12 5928777 N chr12 5929222 N DEL 5
SRR1766464.8127649 chr12 5928769 N chr12 5929728 N DEL 2
SRR1766460.9120995 chr12 5928769 N chr12 5929728 N DEL 4
SRR1766484.3367451 chr12 5928703 N chr12 5929222 N DEL 5
SRR1766454.2961043 chr12 5928904 N chr12 5929715 N DEL 9
SRR1766461.9288666 chr12 5928904 N chr12 5929715 N DEL 9
SRR1766442.13764130 chr12 5928892 N chr12 5929629 N DEL 10
SRR1766442.41978246 chr12 5929269 N chr12 5929782 N DUP 10
SRR1766454.5418474 chr12 5928744 N chr12 5929263 N DEL 10
SRR1766468.2956101 chr12 5928892 N chr12 5929629 N DEL 9
SRR1766444.5430644 chr12 5928744 N chr12 5929263 N DEL 9
SRR1766442.15119110 chr12 5928744 N chr12 5929263 N DEL 8
SRR1766482.2985557 chr12 5928892 N chr12 5929629 N DEL 7
SRR1766478.2533654 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766484.5530922 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766473.2157837 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766442.26905964 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766470.1420152 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766460.2502789 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766483.3214319 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766442.26905964 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766459.4629066 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766456.3939774 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766443.10316276 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766452.7956447 chr12 5928746 N chr12 5929703 N DUP 5
SRR1766475.5056492 chr12 5929424 N chr12 5930087 N DEL 14
SRR1766473.529077 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766455.7828540 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766445.124014 chr12 5928745 N chr12 5930144 N DEL 5
SRR1766475.9371722 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766469.3814881 chr12 5929264 N chr12 5929337 N DUP 5
SRR1766456.4130722 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766465.9405178 chr12 5929269 N chr12 5929782 N DUP 8
SRR1766457.8425680 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766459.4629066 chr12 5929789 N chr12 5930082 N DEL 10
SRR1766442.30776721 chr12 5928898 N chr12 5930149 N DEL 5
SRR1766471.7865627 chr12 5928663 N chr12 5929328 N DUP 10
SRR1766465.9807133 chr12 5928663 N chr12 5929328 N DUP 9
SRR1766447.5098379 chr12 5928770 N chr12 5930095 N DEL 2
SRR1766477.4899102 chr12 5928663 N chr12 5928736 N DUP 10
SRR1766461.10704418 chr12 5928696 N chr12 5929289 N DEL 3
SRR1766453.4061447 chr12 5929358 N chr12 5929723 N DUP 5
SRR1766485.1973263 chr12 5929342 N chr12 5929999 N DUP 1
SRR1766442.43340493 chr12 5928913 N chr12 5929284 N DEL 5
SRR1766454.4674653 chr12 5928681 N chr12 5929274 N DEL 10
SRR1766459.898553 chr12 5928683 N chr12 5929276 N DEL 8
SRR1766479.7657679 chr12 5928918 N chr12 5929289 N DEL 5
SRR1766442.44138396 chr12 5928919 N chr12 5929290 N DEL 5
SRR1766485.7276342 chr12 5928919 N chr12 5929290 N DEL 5
SRR1766442.35696168 chr12 5928925 N chr12 5929296 N DEL 3
SRR1766476.8843704 chr12 5928927 N chr12 5929298 N DEL 1
SRR1766466.4717076 chr12 5928889 N chr12 5929402 N DUP 5
SRR1766469.1265258 chr12 5929367 N chr12 5929804 N DEL 13
SRR1766479.11887998 chr12 5929367 N chr12 5929804 N DEL 1
SRR1766479.12148770 chr12 5929433 N chr12 5929800 N DEL 5
SRR1766454.6793110 chr12 5929418 N chr12 5929493 N DEL 5
SRR1766455.408025 chr12 5929287 N chr12 5929430 N DUP 5
SRR1766477.4271506 chr12 5929422 N chr12 5930011 N DEL 5
SRR1766451.6226572 chr12 5929433 N chr12 5929800 N DEL 6
SRR1766460.9137463 chr12 5929403 N chr12 5930208 N DUP 5
SRR1766442.14279952 chr12 5929422 N chr12 5930085 N DEL 10
SRR1766460.9137463 chr12 5929481 N chr12 5930070 N DEL 5
SRR1766442.11314633 chr12 5929422 N chr12 5930085 N DEL 10
SRR1766459.10593179 chr12 5929422 N chr12 5930085 N DEL 11
SRR1766453.1126053 chr12 5929481 N chr12 5929704 N DEL 4
SRR1766442.40349687 chr12 5929481 N chr12 5929704 N DEL 2
SRR1766472.8895753 chr12 5929419 N chr12 5930082 N DEL 15
SRR1766452.3700988 chr12 5929422 N chr12 5930085 N DEL 15
SRR1766473.529077 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766465.6848241 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766481.4209435 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766474.9457543 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766485.11783333 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766443.1801683 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766469.1366437 chr12 5929481 N chr12 5929704 N DEL 5
SRR1766448.8597871 chr12 5928760 N chr12 5930085 N DEL 10
SRR1766481.7697176 chr12 5928905 N chr12 5929492 N DUP 5
SRR1766458.7161007 chr12 5929487 N chr12 5929782 N DUP 10
SRR1766454.7436758 chr12 5928967 N chr12 5930144 N DEL 5
SRR1766442.6809372 chr12 5928905 N chr12 5929492 N DUP 10
SRR1766477.2409670 chr12 5928905 N chr12 5929492 N DUP 10
SRR1766464.5984668 chr12 5929493 N chr12 5930082 N DEL 10
SRR1766447.8588736 chr12 5929511 N chr12 5929804 N DEL 11
SRR1766442.38379008 chr12 5929074 N chr12 5929513 N DUP 5
SRR1766443.286116 chr12 5928905 N chr12 5929126 N DUP 5
SRR1766443.2697334 chr12 5929511 N chr12 5929804 N DEL 15
SRR1766464.1168502 chr12 5929511 N chr12 5929804 N DEL 6
SRR1766485.6063647 chr12 5929511 N chr12 5929804 N DEL 7
SRR1766476.2299154 chr12 5928714 N chr12 5929599 N DEL 1
SRR1766477.11226155 chr12 5928700 N chr12 5929344 N DUP 2
SRR1766477.11129207 chr12 5928892 N chr12 5929629 N DEL 8
SRR1766442.10393556 chr12 5928744 N chr12 5929263 N DEL 9
SRR1766478.2533654 chr12 5928744 N chr12 5929263 N DEL 10
SRR1766483.11302872 chr12 5928720 N chr12 5929605 N DEL 5
SRR1766442.23668787 chr12 5929650 N chr12 5929867 N DUP 10
SRR1766465.696922 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766442.36054067 chr12 5929337 N chr12 5929630 N DEL 5
SRR1766469.6104689 chr12 5929402 N chr12 5929621 N DEL 5
SRR1766466.2117814 chr12 5929337 N chr12 5929630 N DEL 5
SRR1766442.42200809 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766465.3969839 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766467.692760 chr12 5929126 N chr12 5929641 N DEL 5
SRR1766448.6711066 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766469.9006952 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766460.2502789 chr12 5928744 N chr12 5929263 N DEL 5
SRR1766445.4204844 chr12 5929126 N chr12 5929641 N DEL 5
SRR1766456.3939774 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766463.5892525 chr12 5928663 N chr12 5928810 N DUP 5
SRR1766448.8184556 chr12 5929126 N chr12 5929641 N DEL 5
SRR1766470.250806 chr12 5929126 N chr12 5929641 N DEL 5
SRR1766474.9591594 chr12 5929126 N chr12 5929641 N DEL 5
SRR1766443.1801683 chr12 5929429 N chr12 5929652 N DEL 10
SRR1766482.6561632 chr12 5929337 N chr12 5929630 N DEL 5
SRR1766445.8424435 chr12 5929126 N chr12 5929641 N DEL 5
SRR1766476.6140423 chr12 5928746 N chr12 5929703 N DUP 5
SRR1766466.621726 chr12 5929491 N chr12 5929786 N DUP 10
SRR1766482.2985557 chr12 5928845 N chr12 5929140 N DUP 5
SRR1766446.1555345 chr12 5928663 N chr12 5928810 N DUP 5
SRR1766449.1295593 chr12 5929147 N chr12 5929641 N DEL 5
SRR1766466.10933280 chr12 5929126 N chr12 5929641 N DEL 5
SRR1766469.6428948 chr12 5929132 N chr12 5929647 N DEL 5
SRR1766464.694524 chr12 5929427 N chr12 5929650 N DEL 5
SRR1766477.9709290 chr12 5929357 N chr12 5929724 N DEL 5
SRR1766442.46155632 chr12 5929357 N chr12 5929724 N DEL 5
SRR1766448.6711066 chr12 5929337 N chr12 5929848 N DEL 10
SRR1766442.36126599 chr12 5928978 N chr12 5929715 N DEL 15
SRR1766469.9544908 chr12 5929357 N chr12 5929724 N DEL 5
SRR1766442.17094521 chr12 5928663 N chr12 5930282 N DUP 6
SRR1766456.2078241 chr12 5928905 N chr12 5929492 N DUP 10
SRR1766482.612998 chr12 5928663 N chr12 5930282 N DUP 10
SRR1766469.2484114 chr12 5928978 N chr12 5929715 N DEL 11
SRR1766448.10418503 chr12 5928756 N chr12 5929715 N DEL 10
SRR1766470.10141030 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766481.11343330 chr12 5928756 N chr12 5929715 N DEL 10
SRR1766442.46155632 chr12 5928756 N chr12 5929715 N DEL 10
SRR1766482.10295176 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766442.29850140 chr12 5928756 N chr12 5929715 N DEL 10
SRR1766478.1657900 chr12 5928663 N chr12 5930208 N DUP 9
SRR1766482.11883983 chr12 5928715 N chr12 5929818 N DEL 1
SRR1766473.4342316 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766454.2961043 chr12 5929642 N chr12 5930081 N DUP 10
SRR1766473.3316822 chr12 5928663 N chr12 5928958 N DUP 9
SRR1766465.696922 chr12 5928687 N chr12 5929792 N DUP 13
SRR1766446.9972609 chr12 5928687 N chr12 5929792 N DUP 13
SRR1766459.7056156 chr12 5928687 N chr12 5929792 N DUP 8
SRR1766479.10974705 chr12 5928687 N chr12 5929792 N DUP 15
SRR1766477.2540560 chr12 5928687 N chr12 5929792 N DUP 8
SRR1766459.8171267 chr12 5928687 N chr12 5929792 N DUP 8
SRR1766451.970503 chr12 5928687 N chr12 5929792 N DUP 8
SRR1766466.8360635 chr12 5928687 N chr12 5929792 N DUP 8
SRR1766452.10252382 chr12 5928687 N chr12 5929792 N DUP 8
SRR1766460.6908919 chr12 5928687 N chr12 5929792 N DUP 8
SRR1766454.9626175 chr12 5928687 N chr12 5929792 N DUP 8
SRR1766474.2704687 chr12 5928687 N chr12 5929792 N DUP 14
SRR1766474.7186199 chr12 5928697 N chr12 5929802 N DUP 8
SRR1766466.5373344 chr12 5928687 N chr12 5929792 N DUP 7
SRR1766482.9271944 chr12 5928703 N chr12 5929806 N DEL 5
SRR1766474.2550569 chr12 5928687 N chr12 5929792 N DUP 5
SRR1766445.10593613 chr12 5928704 N chr12 5929807 N DEL 8
SRR1766486.2490837 chr12 5929346 N chr12 5929804 N DEL 13
SRR1766453.7185109 chr12 5929346 N chr12 5929804 N DEL 13
SRR1766462.2937861 chr12 5928703 N chr12 5929806 N DEL 13
SRR1766442.32418744 chr12 5928927 N chr12 5929808 N DEL 10
SRR1766450.3381668 chr12 5928711 N chr12 5929814 N DEL 5
SRR1766467.4086271 chr12 5928663 N chr12 5929912 N DUP 5
SRR1766477.10533136 chr12 5929317 N chr12 5929921 N DUP 5
SRR1766484.7486370 chr12 5929337 N chr12 5929848 N DEL 5
SRR1766454.6337178 chr12 5928663 N chr12 5929912 N DUP 5
SRR1766478.3802562 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766469.4581404 chr12 5928663 N chr12 5929912 N DUP 5
SRR1766468.4458431 chr12 5928663 N chr12 5929912 N DUP 5
SRR1766483.6825840 chr12 5928663 N chr12 5929912 N DUP 5
SRR1766477.2540560 chr12 5928663 N chr12 5929912 N DUP 5
SRR1766466.7490940 chr12 5929354 N chr12 5929865 N DEL 10
SRR1766473.2157837 chr12 5928663 N chr12 5928810 N DUP 5
SRR1766472.7826794 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766485.9868488 chr12 5928663 N chr12 5928958 N DUP 7
SRR1766447.8588736 chr12 5929941 N chr12 5930016 N DEL 3
SRR1766455.408025 chr12 5928899 N chr12 5929782 N DUP 15
SRR1766463.2108008 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766443.9452570 chr12 5928738 N chr12 5929915 N DEL 6
SRR1766444.4841162 chr12 5929789 N chr12 5930082 N DEL 12
SRR1766442.35893354 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766444.5034183 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766479.47885 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766453.1258125 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766463.1949630 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766481.6765539 chr12 5928738 N chr12 5929915 N DEL 5
SRR1766469.9544908 chr12 5928668 N chr12 5928741 N DUP 10
SRR1766483.11302872 chr12 5928738 N chr12 5929915 N DEL 5
SRR1766484.5530922 chr12 5928741 N chr12 5929918 N DEL 5
SRR1766460.700694 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766453.2158332 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766443.6694150 chr12 5929645 N chr12 5929792 N DUP 10
SRR1766465.9789340 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766485.11783333 chr12 5929932 N chr12 5930007 N DEL 10
SRR1766442.30731671 chr12 5929789 N chr12 5930082 N DEL 15
SRR1766469.1101461 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766475.9748323 chr12 5928739 N chr12 5929916 N DEL 5
SRR1766465.11237196 chr12 5929941 N chr12 5930016 N DEL 5
SRR1766477.8070258 chr12 5928691 N chr12 5930016 N DEL 5
SRR1766482.11883983 chr12 5928691 N chr12 5930016 N DEL 5
SRR1766443.9452570 chr12 5928684 N chr12 5930009 N DEL 10
SRR1766459.7056156 chr12 5928691 N chr12 5930016 N DEL 5
SRR1766473.4342316 chr12 5929337 N chr12 5929848 N DEL 10
SRR1766466.621726 chr12 5929622 N chr12 5929989 N DEL 7
SRR1766474.10714393 chr12 5928894 N chr12 5929337 N DUP 10
SRR1766445.8424435 chr12 5928745 N chr12 5929996 N DEL 5
SRR1766477.8896701 chr12 5929348 N chr12 5929419 N DEL 2
SRR1766470.8846594 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766455.7006375 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766485.4395842 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766457.9159348 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766469.8222562 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766464.7176388 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766469.4581404 chr12 5929337 N chr12 5929408 N DEL 5
SRR1766459.9871686 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766442.43671427 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766477.7193919 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766454.6793110 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766464.5984668 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766452.3497594 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766464.10305591 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766454.9626175 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766466.8360635 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766478.5441170 chr12 5929525 N chr12 5929746 N DUP 10
SRR1766481.4209435 chr12 5929501 N chr12 5929650 N DEL 10
SRR1766485.9868488 chr12 5929337 N chr12 5929408 N DEL 5
SRR1766483.11606358 chr12 5930008 N chr12 5930081 N DUP 5
SRR1766446.379038 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766457.5649116 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766466.1999136 chr12 5929777 N chr12 5930292 N DEL 10
SRR1766442.6809372 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766466.5373344 chr12 5929777 N chr12 5930292 N DEL 12
SRR1766469.6573479 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766453.4612066 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766461.6745378 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766442.42200809 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766457.6410389 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766447.1963712 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766486.7747891 chr12 5929650 N chr12 5929723 N DUP 5
SRR1766469.1366437 chr12 5928685 N chr12 5930010 N DEL 1
SRR1766485.6063647 chr12 5928686 N chr12 5930011 N DEL 10
SRR1766464.4366081 chr12 5929511 N chr12 5929804 N DEL 10
SRR1766442.17094521 chr12 5929511 N chr12 5929804 N DEL 10
SRR1766442.35893354 chr12 5929501 N chr12 5929942 N DEL 5
SRR1766448.8184556 chr12 5929276 N chr12 5930081 N DUP 5
SRR1766459.5087434 chr12 5929944 N chr12 5930091 N DUP 5
SRR1766468.6179614 chr12 5929504 N chr12 5929945 N DEL 5
SRR1766443.2697334 chr12 5930082 N chr12 5930155 N DUP 5
SRR1766475.2447978 chr12 5930082 N chr12 5930155 N DUP 5
SRR1766481.380493 chr12 5929650 N chr12 5930089 N DUP 1
SRR1766477.2327514 chr12 5929650 N chr12 5930089 N DUP 2
SRR1766454.3533588 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766455.1715408 chr12 5929650 N chr12 5930089 N DUP 4
SRR1766442.10393556 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766461.7625844 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766469.280951 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766479.13942330 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766467.9779245 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766461.10315855 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766456.2078241 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766485.10841502 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766442.44947228 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766456.2926143 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766460.3972483 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766472.2203981 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766482.612998 chr12 5929402 N chr12 5930061 N DEL 5
SRR1766482.9184375 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766467.8225961 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766452.736183 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766449.1295593 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766458.431038 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766470.397577 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766485.9306232 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766442.1774884 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766460.6908919 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766458.2176834 chr12 5929650 N chr12 5930089 N DUP 5
SRR1766463.4931578 chr12 5928894 N chr12 5929777 N DUP 10
SRR1766443.2920217 chr12 5929148 N chr12 5930082 N DEL 5
SRR1766473.4409993 chr12 5929148 N chr12 5930082 N DEL 5
SRR1766442.36126599 chr12 5929420 N chr12 5930081 N DUP 5
SRR1766464.6713334 chr12 5929148 N chr12 5930082 N DEL 5
SRR1766469.280951 chr12 5929128 N chr12 5930083 N DEL 7
SRR1766482.9718139 chr12 5928762 N chr12 5928911 N DEL 1
SRR1766462.3574483 chr12 5929351 N chr12 5930084 N DEL 5
SRR1766481.10437318 chr12 5929129 N chr12 5930084 N DEL 6
SRR1766446.3914326 chr12 5929130 N chr12 5930085 N DEL 5
SRR1766443.2920217 chr12 5929132 N chr12 5930087 N DEL 5
SRR1766452.736183 chr12 5929133 N chr12 5930088 N DEL 5
SRR1766442.4932921 chr12 5929512 N chr12 5930101 N DEL 5
SRR1766481.3893534 chr12 5928663 N chr12 5930208 N DUP 3
SRR1766469.2360231 chr12 5929504 N chr12 5930093 N DEL 3
SRR1766458.431038 chr12 5929505 N chr12 5930094 N DEL 3
SRR1766458.19027 chr12 5929506 N chr12 5930095 N DEL 1
SRR1766442.11314633 chr12 5928919 N chr12 5929656 N DEL 2
SRR1766451.7079322 chr12 5928688 N chr12 5930087 N DEL 6
SRR1766466.4717076 chr12 5929419 N chr12 5930080 N DUP 5
SRR1766443.10787393 chr12 5930082 N chr12 5930155 N DUP 5
SRR1766468.5407746 chr12 5930082 N chr12 5930155 N DUP 5
SRR1766484.3367451 chr12 5929264 N chr12 5929337 N DUP 5
SRR1766442.38379008 chr12 5928745 N chr12 5930144 N DEL 5
SRR1766442.30731671 chr12 5929548 N chr12 5929915 N DEL 10
SRR1766481.10437318 chr12 5929074 N chr12 5929369 N DUP 5
SRR1766478.5441170 chr12 5929380 N chr12 5929525 N DEL 5
SRR1766452.10233021 chr12 5929380 N chr12 5929525 N DEL 5
SRR1766445.9524992 chr12 5929348 N chr12 5929641 N DEL 5
SRR1766470.8567927 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766458.19027 chr12 5929380 N chr12 5929525 N DEL 5
SRR1766464.6713334 chr12 5929380 N chr12 5929525 N DEL 5
SRR1766480.6408445 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766442.1774884 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766460.7818145 chr12 5929349 N chr12 5930082 N DEL 5
SRR1766482.9718139 chr12 5928903 N chr12 5929786 N DUP 10
SRR1766447.4117854 chr12 5929380 N chr12 5929525 N DEL 5
SRR1766442.14279952 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766466.10933280 chr12 5929348 N chr12 5929641 N DEL 5
SRR1766444.4841162 chr12 5929269 N chr12 5929782 N DUP 10
SRR1766465.9789340 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766459.5087434 chr12 5928663 N chr12 5930208 N DUP 10
SRR1766476.2299154 chr12 5929264 N chr12 5929337 N DUP 5
SRR1766446.7710642 chr12 5929348 N chr12 5929641 N DEL 5
SRR1766479.10974705 chr12 5929269 N chr12 5929782 N DUP 10
SRR1766460.7818145 chr12 5928684 N chr12 5930081 N DUP 5
SRR1766482.11626741 chr12 5928746 N chr12 5930145 N DEL 5
SRR1766445.9524992 chr12 5929147 N chr12 5929641 N DEL 5
SRR1766485.2140434 chr12 5929132 N chr12 5930161 N DEL 5
SRR1766465.8169581 chr12 5929148 N chr12 5930082 N DEL 5
SRR1766454.6337178 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766486.2490837 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766474.9591594 chr12 5929723 N chr12 5930238 N DEL 5
SRR1766464.1168502 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766479.490704 chr12 5929723 N chr12 5930238 N DEL 5
SRR1766465.3724642 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766470.2808913 chr12 5930143 N chr12 5930292 N DEL 15
SRR1766446.9972609 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766474.9457543 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766470.10141030 chr12 5928703 N chr12 5930229 N DEL 6
SRR1766455.5300617 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766455.5652074 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766460.700694 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766456.998954 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766469.9006952 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766453.7185109 chr12 5929777 N chr12 5930292 N DEL 15
SRR1766452.10252382 chr12 5929777 N chr12 5930292 N DEL 11
SRR1766469.1101461 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766477.7193919 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766482.9184375 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766460.2497917 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766467.4086271 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766474.3521928 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766474.2550569 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766465.3807061 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766474.11667806 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766462.3698742 chr12 5929337 N chr12 5930292 N DEL 10
SRR1766460.10344977 chr12 5929341 N chr12 5930296 N DEL 10
SRR1766451.970503 chr12 5929343 N chr12 5930298 N DEL 9
SRR1766443.3802752 chr12 5928702 N chr12 5930302 N DEL 5
SRR1766453.8627402 chr12 5929148 N chr12 5930304 N DEL 3
SRR1766472.9864054 chr12 5929148 N chr12 5930304 N DEL 3
SRR1766475.4296516 chr20 2545990 N chr20 2546056 N DEL 9
SRR1766443.4566253 chr20 2545987 N chr20 2546057 N DEL 8
SRR1766442.46129327 chr3 186874254 N chr3 186874380 N DUP 3
SRR1766482.11871869 chr3 186874222 N chr3 186874348 N DUP 12
SRR1766480.3278339 chr3 186874289 N chr3 186874415 N DUP 3
SRR1766464.6003588 chr3 186874289 N chr3 186874415 N DUP 4
SRR1766446.4443472 chr3 186874308 N chr3 186874436 N DEL 5
SRR1766483.7398782 chr3 186874415 N chr3 186874494 N DEL 18
SRR1766452.3029510 chr3 186874415 N chr3 186874494 N DEL 15
SRR1766476.1240892 chr3 186874415 N chr3 186874494 N DEL 6
SRR1766469.8783793 chr3 186874314 N chr3 186874520 N DEL 5
SRR1766458.5183475 chr3 186874427 N chr3 186874506 N DEL 3
SRR1766442.29156713 chr3 186874259 N chr3 186874639 N DUP 5
SRR1766468.84702 chr19 458138 N chr19 458244 N DEL 10
SRR1766480.1331210 chr19 458207 N chr19 458271 N DEL 4
SRR1766471.6951142 chr19 458083 N chr19 458420 N DUP 3
SRR1766469.3430450 chr19 458293 N chr19 458401 N DEL 1
SRR1766442.11916446 chr19 458096 N chr19 458435 N DEL 1
SRR1766484.3181995 chr19 458444 N chr19 458527 N DUP 5
SRR1766457.3658035 chr19 458118 N chr19 458499 N DEL 9
SRR1766473.6366295 chr19 458643 N chr19 458919 N DEL 7
SRR1766474.5822874 chr19 458133 N chr19 458577 N DEL 7
SRR1766448.5375515 chr19 458594 N chr19 458974 N DUP 5
SRR1766458.1689509 chr19 458138 N chr19 458582 N DEL 5
SRR1766447.1320653 chr19 458137 N chr19 458687 N DEL 13
SRR1766476.5952379 chr19 458094 N chr19 458665 N DEL 3
SRR1766458.1639952 chr19 458758 N chr19 458907 N DEL 10
SRR1766466.7941485 chr19 458294 N chr19 458697 N DEL 10
SRR1766473.11828876 chr19 458118 N chr19 458795 N DEL 5
SRR1766475.7379843 chr19 458437 N chr19 458943 N DUP 5
SRR1766449.8867811 chr19 458708 N chr19 458921 N DEL 8
SRR1766470.8196713 chr7 63204972 N chr7 63205169 N DEL 14
SRR1766471.4577455 chr7 63204931 N chr7 63205024 N DEL 4
SRR1766468.4568942 chr7 63205043 N chr7 63205176 N DUP 1
SRR1766457.342788 chr7 63205043 N chr7 63205176 N DUP 4
SRR1766472.10527916 chr15 71564768 N chr15 71564908 N DEL 2
SRR1766449.7381438 chr15 71564768 N chr15 71564908 N DEL 9
SRR1766456.4752867 chr15 71564768 N chr15 71564908 N DEL 9
SRR1766456.3732264 chr15 71564768 N chr15 71564908 N DEL 9
SRR1766452.6745644 chr15 71564790 N chr15 71564844 N DEL 9
SRR1766461.9163271 chr15 71564790 N chr15 71564844 N DEL 9
SRR1766470.3843351 chr15 71564790 N chr15 71564844 N DEL 9
SRR1766442.6917233 chr15 71564790 N chr15 71564844 N DEL 9
SRR1766478.9800619 chr15 71564790 N chr15 71564844 N DEL 9
SRR1766475.11381165 chr15 71564790 N chr15 71564844 N DEL 9
SRR1766472.1745233 chr15 71564790 N chr15 71564844 N DEL 9
SRR1766459.3512587 chr15 71564843 N chr15 71564930 N DEL 1
SRR1766477.3574256 chr15 71564790 N chr15 71564844 N DEL 10
SRR1766450.7543360 chr15 71564790 N chr15 71564844 N DEL 11
SRR1766449.6751310 chr15 71564790 N chr15 71564844 N DEL 12
SRR1766444.6700862 chr15 71564814 N chr15 71564954 N DUP 9
SRR1766478.4747262 chr15 71564845 N chr15 71564932 N DEL 4
SRR1766451.3683453 chr15 71564845 N chr15 71564932 N DEL 6
SRR1766469.8199101 chr15 71564845 N chr15 71564932 N DEL 7
SRR1766472.4491762 chr15 71564912 N chr15 71565004 N DEL 8
SRR1766470.3843351 chr15 71564853 N chr15 71564940 N DEL 5
SRR1766459.10928820 chr11 119037058 N chr11 119037364 N DUP 4
SRR1766471.7932281 chr19 8706747 N chr19 8706807 N DEL 5
SRR1766478.6594404 chr19 8706747 N chr19 8706807 N DEL 5
SRR1766460.3034318 chr2 239101976 N chr2 239102047 N DUP 5
SRR1766449.4559818 chr2 239102001 N chr2 239102182 N DEL 5
SRR1766480.7910161 chr2 239101994 N chr2 239102247 N DEL 10
SRR1766480.1797953 chr2 239102014 N chr2 239102267 N DEL 3
SRR1766479.13252914 chr2 239102056 N chr2 239102273 N DEL 5
SRR1766463.9401207 chr2 239101938 N chr2 239102299 N DEL 5
SRR1766472.11743302 chr10 128471795 N chr10 128472098 N DUP 5
SRR1766473.7274060 chr19 10187650 N chr19 10187918 N DEL 1
SRR1766456.654239 chr19 10187807 N chr19 10188081 N DEL 10
SRR1766461.11214300 chr19 10187853 N chr19 10188128 N DEL 5
SRR1766475.8093420 chr19 10187539 N chr19 10187807 N DEL 8
SRR1766442.20040263 chr19 10187585 N chr19 10187853 N DEL 5
SRR1766443.8247274 chr19 10187596 N chr19 10187864 N DEL 5
SRR1766442.6530790 chr19 10187577 N chr19 10187978 N DEL 5
SRR1766465.7024414 chr4 49087720 N chr4 49088406 N DUP 2
SRR1766443.7694139 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766472.8841768 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766465.3363995 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766486.4610671 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766485.8831445 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766454.6798768 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766442.45946760 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766445.542444 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766465.8587520 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766466.9789165 chr21 44953585 N chr21 44953635 N DUP 5
SRR1766462.9382248 chr21 44953585 N chr21 44953635 N DUP 7
SRR1766442.12641961 chr21 44953585 N chr21 44953635 N DUP 8
SRR1766466.4287147 chr21 44953585 N chr21 44953635 N DUP 17
SRR1766463.8860220 chr21 44953585 N chr21 44953635 N DUP 17
SRR1766442.29204173 chr21 44953585 N chr21 44953635 N DUP 19
SRR1766450.862540 chr5 181444879 N chr5 181445014 N DEL 1
SRR1766465.6000768 chr8 28882646 N chr8 28882702 N DUP 14
SRR1766485.7409267 chr8 28882640 N chr8 28882696 N DUP 14
SRR1766442.31660393 chr8 28882644 N chr8 28882696 N DUP 15
SRR1766471.6398489 chr13 100986616 N chr13 100986681 N DUP 5
SRR1766484.3553280 chr13 100986616 N chr13 100986681 N DUP 5
SRR1766449.4909111 chr5 142993504 N chr5 142993639 N DEL 5
SRR1766446.5257225 chr12 122093067 N chr12 122093251 N DEL 21
SRR1766486.11178811 chr12 122093068 N chr12 122093269 N DUP 10
SRR1766463.8847399 chr12 122093069 N chr12 122093270 N DUP 10
SRR1766467.9364829 chr12 122093071 N chr12 122093272 N DUP 8
SRR1766486.10501349 chr12 122093073 N chr12 122093274 N DUP 6
SRR1766442.20135552 chr12 122093077 N chr12 122093278 N DUP 4
SRR1766448.8097575 chr12 122093230 N chr12 122093288 N DUP 1
SRR1766479.8152338 chr3 49393906 N chr3 49394068 N DEL 5
SRR1766479.4216713 chr16 13019917 N chr16 13020031 N DUP 5
SRR1766452.1592492 chr16 13019916 N chr16 13020021 N DUP 15
SRR1766460.2282043 chr16 13019916 N chr16 13020021 N DUP 15
SRR1766457.6574383 chr16 13019917 N chr16 13020031 N DUP 5
SRR1766476.2207930 chr16 13019949 N chr16 13020189 N DUP 2
SRR1766442.3573146 chr16 13019917 N chr16 13020031 N DUP 5
SRR1766469.3982793 chr16 13019917 N chr16 13020031 N DUP 5
SRR1766466.8890728 chr16 13019917 N chr16 13020031 N DUP 5
SRR1766455.7956030 chr16 13019931 N chr16 13020047 N DEL 2
SRR1766478.2002723 chr10 668230 N chr10 668382 N DUP 5
SRR1766480.7643360 chr10 668230 N chr10 668382 N DUP 5
SRR1766444.2974746 chr10 668230 N chr10 668382 N DUP 5
SRR1766444.5633944 chr10 668230 N chr10 668382 N DUP 5
SRR1766454.7787447 chr10 668230 N chr10 668382 N DUP 5
SRR1766464.4148186 chr10 668230 N chr10 668382 N DUP 5
SRR1766469.11065821 chr10 668230 N chr10 668382 N DUP 5
SRR1766481.3505041 chr10 668230 N chr10 668382 N DUP 5
SRR1766468.5097600 chr10 668230 N chr10 668382 N DUP 5
SRR1766444.3341258 chr10 668230 N chr10 668382 N DUP 5
SRR1766449.6311578 chr10 668230 N chr10 668382 N DUP 5
SRR1766482.8031130 chr10 668230 N chr10 668382 N DUP 5
SRR1766451.280237 chr10 668230 N chr10 668382 N DUP 5
SRR1766475.6543279 chr10 668230 N chr10 668382 N DUP 5
SRR1766452.1415 chr10 668242 N chr10 668385 N DUP 3
SRR1766467.9968778 chr10 668243 N chr10 668386 N DUP 2
SRR1766460.381290 chr10 668221 N chr10 668376 N DEL 6
SRR1766442.10577646 chr9 65464219 N chr9 65464278 N DEL 5
SRR1766449.1774351 chrX 70371885 N chrX 70372083 N DEL 3
SRR1766468.1999444 chr10 86278044 N chr10 86278115 N DEL 5
SRR1766443.8718823 chr22 37227322 N chr22 37227433 N DEL 5
SRR1766484.3780150 chr16 6773320 N chr16 6773422 N DUP 13
SRR1766457.4703329 chr16 6773320 N chr16 6773424 N DUP 15
SRR1766463.7334598 chr16 6773360 N chr16 6773423 N DUP 5
SRR1766452.9864072 chr21 5329582 N chr21 5329646 N DUP 14
SRR1766474.892858 chr21 5329574 N chr21 5329703 N DUP 21
SRR1766475.2202814 chr21 5329585 N chr21 5329748 N DUP 7
SRR1766475.6352302 chr21 5329585 N chr21 5329748 N DUP 7
SRR1766457.4518083 chr21 5329585 N chr21 5329748 N DUP 7
SRR1766465.3153599 chr21 5329602 N chr21 5329755 N DUP 27
SRR1766453.5341573 chr21 5329659 N chr21 5329791 N DUP 5
SRR1766449.7799874 chr21 5329580 N chr21 5329812 N DUP 10
SRR1766479.7490592 chr21 5329582 N chr21 5329814 N DUP 5
SRR1766480.4383793 chr21 5329567 N chr21 5329799 N DUP 5
SRR1766453.6875770 chr21 5329767 N chr21 5329841 N DUP 15
SRR1766473.3399697 chr10 106130096 N chr10 106130191 N DUP 5
SRR1766481.400046 chr11 473722 N chr11 473791 N DEL 2
SRR1766457.7733511 chr11 473723 N chr11 473858 N DUP 20
SRR1766485.5375791 chr11 473723 N chr11 473858 N DUP 20
SRR1766462.2752522 chr11 473723 N chr11 473858 N DUP 19
SRR1766442.16078834 chr11 473726 N chr11 473861 N DUP 12
SRR1766461.8911752 chr11 473777 N chr11 473844 N DUP 24
SRR1766483.6063020 chr11 473723 N chr11 473858 N DUP 20
SRR1766463.966182 chr11 473723 N chr11 473858 N DUP 22
SRR1766464.10301700 chr11 473788 N chr11 473855 N DUP 6
SRR1766480.5103384 chr11 473788 N chr11 473855 N DUP 7
SRR1766462.1490056 chr11 473788 N chr11 473855 N DUP 12
SRR1766462.209330 chr11 473797 N chr11 473864 N DUP 4
SRR1766444.5233288 chr11 473802 N chr11 473869 N DUP 1
SRR1766459.7007257 chr8 111208388 N chr8 111208439 N DEL 4
SRR1766445.1425739 chr8 3684367 N chr8 3684441 N DUP 1
SRR1766453.4528416 chr8 3684366 N chr8 3684440 N DUP 2
SRR1766473.6994441 chr9 9275208 N chr9 9275278 N DEL 5
SRR1766485.1878805 chr9 9275208 N chr9 9275278 N DEL 6
SRR1766452.4597343 chr9 9275208 N chr9 9275278 N DEL 10
SRR1766462.8462440 chr9 9275257 N chr9 9275359 N DEL 13
SRR1766468.3017360 chr9 9275215 N chr9 9275332 N DUP 1
SRR1766477.8589842 chr9 9275239 N chr9 9275296 N DEL 7
SRR1766446.8531159 chr9 9275243 N chr9 9275349 N DEL 18
SRR1766482.5720344 chr9 9275243 N chr9 9275349 N DEL 18
SRR1766442.35607042 chr9 9275231 N chr9 9275363 N DEL 1
SRR1766449.6263565 chr9 9275249 N chr9 9275355 N DEL 9
SRR1766467.9985835 chr9 9275230 N chr9 9275362 N DEL 2
SRR1766443.8415002 chr9 9275251 N chr9 9275357 N DEL 7
SRR1766461.1201163 chr2 241011217 N chr2 241011416 N DEL 5
SRR1766451.1522215 chr2 241011203 N chr2 241011303 N DEL 9
SRR1766481.12411270 chr2 241011249 N chr2 241011385 N DEL 3
SRR1766446.6455652 chr2 241011227 N chr2 241011291 N DEL 28
SRR1766468.2737368 chr2 241011227 N chr2 241011291 N DEL 28
SRR1766465.9371366 chr2 241011261 N chr2 241011388 N DEL 28
SRR1766460.4052463 chr2 241011233 N chr2 241011396 N DEL 7
SRR1766477.8595857 chr2 241011231 N chr2 241011394 N DEL 9
SRR1766481.1439889 chr2 241011386 N chr2 241011450 N DEL 7
SRR1766461.5205440 chr1 228633475 N chr1 228633534 N DUP 12
SRR1766454.7963000 chr1 228633477 N chr1 228633530 N DUP 11
SRR1766456.5628066 chr1 163552239 N chr1 163552396 N DEL 15
SRR1766462.7106137 chr1 163552239 N chr1 163552357 N DEL 10
SRR1766463.8009831 chr1 163552352 N chr1 163552470 N DEL 3
SRR1766473.2655725 chr1 163552352 N chr1 163552470 N DEL 3
SRR1766442.6191757 chr1 163552352 N chr1 163552470 N DEL 5
SRR1766482.6943266 chr1 163552268 N chr1 163552386 N DEL 1
SRR1766474.847799 chr1 163552352 N chr1 163552470 N DEL 5
SRR1766465.7518315 chr1 163552352 N chr1 163552470 N DEL 5
SRR1766449.7808572 chr1 163552352 N chr1 163552470 N DEL 5
SRR1766442.26073377 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766458.8700375 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766472.11303882 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766462.1368119 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766442.36329790 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766468.4475192 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766471.11604121 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766466.2028982 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766480.514657 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766449.1273778 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766445.1753639 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766451.6358073 chr1 163552313 N chr1 163552470 N DEL 5
SRR1766446.3651710 chr1 163552274 N chr1 163552470 N DEL 5
SRR1766460.5590367 chr1 163552274 N chr1 163552470 N DEL 5
SRR1766473.10855273 chr1 163552277 N chr1 163552473 N DEL 5
SRR1766443.5225866 chr1 163552282 N chr1 163552478 N DEL 5
SRR1766465.8606810 chr2 90382982 N chr2 90383080 N DUP 4
SRR1766442.44251767 chr2 90382996 N chr2 90383045 N DUP 10
SRR1766470.6503296 chr2 90382998 N chr2 90383096 N DUP 10
SRR1766450.4689519 chr2 90382908 N chr2 90383001 N DEL 9
SRR1766473.10885932 chr2 90382908 N chr2 90383001 N DEL 9
SRR1766442.11321687 chr2 90382908 N chr2 90383001 N DEL 9
SRR1766451.1742719 chr2 90382908 N chr2 90383001 N DEL 9
SRR1766468.1435195 chr2 90382908 N chr2 90383001 N DEL 9
SRR1766458.7357316 chr2 90382973 N chr2 90383024 N DEL 1
SRR1766483.6412559 chr2 90382922 N chr2 90383138 N DUP 5
SRR1766442.30844760 chr2 90383099 N chr2 90383170 N DUP 35
SRR1766454.9242232 chr2 90383099 N chr2 90383170 N DUP 35
SRR1766485.2300572 chr2 90383099 N chr2 90383170 N DUP 6
SRR1766460.10535913 chr2 90383099 N chr2 90383170 N DUP 26
SRR1766466.6694867 chr2 90383099 N chr2 90383170 N DUP 26
SRR1766463.10078175 chr2 90383099 N chr2 90383170 N DUP 29
SRR1766484.10631252 chr2 90383099 N chr2 90383170 N DUP 30
SRR1766450.7941652 chr2 90383099 N chr2 90383170 N DUP 24
SRR1766461.3283016 chr2 90383099 N chr2 90383170 N DUP 24
SRR1766475.4116566 chr2 90383068 N chr2 90383214 N DUP 5
SRR1766447.11136813 chr2 90383099 N chr2 90383170 N DUP 23
SRR1766475.459621 chr2 90383099 N chr2 90383170 N DUP 20
SRR1766442.11179299 chr2 90383047 N chr2 90383193 N DUP 2
SRR1766448.7807302 chr2 90383047 N chr2 90383193 N DUP 2
SRR1766449.2141428 chr2 90383047 N chr2 90383193 N DUP 2
SRR1766454.3231859 chr2 90383047 N chr2 90383193 N DUP 2
SRR1766447.7529369 chr2 90383047 N chr2 90383193 N DUP 3
SRR1766461.1492227 chr2 90383047 N chr2 90383193 N DUP 3
SRR1766463.9575886 chr2 90383047 N chr2 90383193 N DUP 3
SRR1766443.9365416 chr2 90383047 N chr2 90383193 N DUP 4
SRR1766451.8996215 chr2 90383047 N chr2 90383193 N DUP 4
SRR1766474.11291487 chr2 90383047 N chr2 90383193 N DUP 4
SRR1766445.2121148 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766445.754935 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766459.5669896 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766472.697615 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766485.461438 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766450.1988474 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766476.7601221 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766448.4489752 chr2 90383062 N chr2 90383135 N DEL 43
SRR1766455.2767355 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766445.8870731 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766458.392582 chr2 90383047 N chr2 90383193 N DUP 5
SRR1766477.5099405 chr2 90383062 N chr2 90383135 N DEL 40
SRR1766485.3592883 chr2 90383062 N chr2 90383135 N DEL 42
SRR1766471.6817426 chr2 90383062 N chr2 90383135 N DEL 40
SRR1766462.8685547 chr2 90383016 N chr2 90383089 N DEL 5
SRR1766477.6899514 chr2 90382907 N chr2 90383099 N DEL 2
SRR1766453.8932800 chr2 90383062 N chr2 90383135 N DEL 35
SRR1766463.7684069 chr2 90383062 N chr2 90383135 N DEL 35
SRR1766445.4784805 chr2 90383109 N chr2 90383206 N DUP 5
SRR1766447.4917476 chr2 90383109 N chr2 90383206 N DUP 5
SRR1766450.4395789 chr2 90383109 N chr2 90383206 N DUP 5
SRR1766481.10654764 chr2 90383062 N chr2 90383135 N DEL 35
SRR1766442.26962507 chr2 90383114 N chr2 90383241 N DUP 6
SRR1766442.27521889 chr2 90383114 N chr2 90383241 N DUP 6
SRR1766464.8116009 chr2 90383062 N chr2 90383135 N DEL 33
SRR1766461.8465301 chr10 83462788 N chr10 83462853 N DUP 5
SRR1766467.10176985 chr10 83462788 N chr10 83462853 N DUP 5
SRR1766480.2428879 chr10 83462788 N chr10 83462919 N DUP 15
SRR1766481.5204538 chr10 83462829 N chr10 83462919 N DUP 5
SRR1766486.9713072 chr10 83462829 N chr10 83462919 N DUP 5
SRR1766455.8202442 chr10 83462829 N chr10 83462919 N DUP 6
SRR1766462.1054385 chr10 83462829 N chr10 83462919 N DUP 7
SRR1766452.447774 chr10 83462829 N chr10 83462919 N DUP 12
SRR1766447.11314208 chr10 83462899 N chr10 83462964 N DUP 10
SRR1766457.8216012 chr10 83462899 N chr10 83462964 N DUP 10
SRR1766471.2227315 chr10 83462788 N chr10 83462919 N DUP 2
SRR1766485.4060272 chr10 83462788 N chr10 83462853 N DUP 5
SRR1766471.1078669 chr1 3176218 N chr1 3176301 N DUP 2
SRR1766470.1476081 chr1 3176212 N chr1 3176430 N DUP 15
SRR1766477.2715023 chr1 3176257 N chr1 3176308 N DUP 1
SRR1766471.5282663 chr1 3176228 N chr1 3176309 N DEL 8
SRR1766474.10155820 chr1 3176110 N chr1 3176307 N DEL 10
SRR1766455.3959176 chr1 3176302 N chr1 3176428 N DUP 11
SRR1766481.4459235 chr1 3176302 N chr1 3176420 N DUP 2
SRR1766484.8102668 chr1 3176315 N chr1 3176449 N DUP 5
SRR1766446.2714963 chr1 3176302 N chr1 3176436 N DUP 20
SRR1766479.12487080 chr1 3176306 N chr1 3176440 N DUP 15
SRR1766460.7839088 chr1 3176212 N chr1 3176438 N DUP 32
SRR1766455.3605592 chr1 3176329 N chr1 3176413 N DEL 3
SRR1766445.894973 chr16 74110149 N chr16 74110206 N DUP 6
SRR1766473.7451091 chr16 74110149 N chr16 74110206 N DUP 6
SRR1766475.7440242 chr1 1905799 N chr1 1905963 N DUP 5
SRR1766445.2735723 chr1 1905712 N chr1 1905878 N DEL 5
SRR1766486.1914575 chr1 1905717 N chr1 1905883 N DEL 5
SRR1766459.5469991 chr19 46179263 N chr19 46179498 N DEL 1
SRR1766466.9152651 chr19 46179282 N chr19 46179397 N DEL 5
SRR1766470.3357621 chr8 70935280 N chr8 70935363 N DEL 10
SRR1766473.7952460 chr8 70935279 N chr8 70935362 N DEL 11
SRR1766482.9816880 chr8 70935282 N chr8 70935363 N DEL 10
SRR1766476.2528652 chr6 54310806 N chr6 54310872 N DEL 5
SRR1766481.1926376 chr6 54310807 N chr6 54310873 N DEL 6
SRR1766444.2675616 chr6 54310807 N chr6 54310873 N DEL 20
SRR1766484.7499008 chr6 54310807 N chr6 54310873 N DEL 20
SRR1766442.7384271 chr6 54310807 N chr6 54310873 N DEL 25
SRR1766484.1628542 chr6 54310807 N chr6 54310873 N DEL 36
SRR1766442.26017437 chr6 54310807 N chr6 54310873 N DEL 40
SRR1766484.5243983 chr6 54310807 N chr6 54310873 N DEL 43
SRR1766443.5192120 chr6 54310807 N chr6 54310873 N DEL 45
SRR1766442.17971201 chr6 54310807 N chr6 54310873 N DEL 46
SRR1766446.5989979 chr6 54310807 N chr6 54310873 N DEL 49
SRR1766444.2675616 chr6 54310807 N chr6 54310873 N DEL 20
SRR1766442.7384271 chr6 54310807 N chr6 54310873 N DEL 18
SRR1766471.10140423 chr6 54310807 N chr6 54310873 N DEL 16
SRR1766446.2649280 chr6 54310816 N chr6 54310882 N DEL 6
SRR1766442.37386087 chr6 54310820 N chr6 54310886 N DEL 2
SRR1766448.9488474 chr6 54310820 N chr6 54310886 N DEL 2
SRR1766454.3308544 chr6 54310796 N chr6 54311048 N DUP 4
SRR1766464.9081865 chr6 54310796 N chr6 54311048 N DUP 5
SRR1766473.3722528 chr6 54310796 N chr6 54311048 N DUP 6
SRR1766465.1357339 chr6 54310796 N chr6 54311048 N DUP 6
SRR1766462.6687958 chr6 54310796 N chr6 54311048 N DUP 10
SRR1766468.997017 chr6 54310970 N chr6 54311048 N DEL 23
SRR1766449.9094744 chr6 54310813 N chr6 54311061 N DEL 7
SRR1766477.830569 chr6 54310812 N chr6 54311060 N DEL 8
SRR1766483.1013626 chr6 54310812 N chr6 54311060 N DEL 8
SRR1766442.9332335 chr7 155354490 N chr7 155354542 N DEL 1
SRR1766472.2621741 chr7 155354466 N chr7 155354518 N DEL 3
SRR1766482.3714742 chr7 155354466 N chr7 155354518 N DEL 4
SRR1766450.3037937 chr7 155354466 N chr7 155354518 N DEL 8
SRR1766444.5737758 chr7 155354476 N chr7 155354641 N DUP 5
SRR1766470.5693280 chr7 155354477 N chr7 155354642 N DUP 5
SRR1766457.7498004 chr7 155354508 N chr7 155354572 N DUP 24
SRR1766460.5330172 chr7 155354508 N chr7 155354572 N DUP 24
SRR1766464.437873 chr7 155354509 N chr7 155354573 N DUP 23
SRR1766472.164914 chr7 155354509 N chr7 155354573 N DUP 23
SRR1766459.5453688 chr7 155354509 N chr7 155354573 N DUP 22
SRR1766465.1609469 chrX 131137591 N chrX 131137766 N DEL 5
SRR1766471.4680582 chrX 131137445 N chrX 131137548 N DEL 5
SRR1766455.5244457 chrX 131137449 N chrX 131137552 N DEL 5
SRR1766458.8050783 chrX 131137435 N chrX 131137606 N DEL 1
SRR1766481.1037428 chrX 131137841 N chrX 131137936 N DUP 3
SRR1766478.7433986 chrX 131137741 N chrX 131138118 N DEL 5
SRR1766445.8402715 chrX 131138119 N chrX 131138524 N DUP 4
SRR1766482.2157800 chrX 131138107 N chrX 131138174 N DEL 12
SRR1766471.10383777 chrX 131138107 N chrX 131138174 N DEL 9
SRR1766442.44115444 chrX 131138322 N chrX 131138509 N DEL 4
SRR1766442.36906329 chrX 131138290 N chrX 131138509 N DEL 5
SRR1766449.7390739 chr3 98836967 N chr3 98837064 N DUP 5
SRR1766445.5892672 chr3 98837069 N chr3 98837246 N DUP 9
SRR1766478.6655777 chr3 98836939 N chr3 98837163 N DUP 2
SRR1766463.5269002 chr3 98836950 N chr3 98837049 N DEL 5
SRR1766476.8579295 chr3 98837019 N chr3 98837182 N DUP 13
SRR1766442.12693224 chr3 98836980 N chr3 98837206 N DUP 5
SRR1766479.5507843 chr3 98836936 N chr3 98837211 N DUP 5
SRR1766472.8978002 chr3 98836936 N chr3 98837211 N DUP 5
SRR1766462.794707 chr3 98836932 N chr3 98837207 N DUP 10
SRR1766443.9639002 chr3 98836936 N chr3 98837211 N DUP 5
SRR1766480.675749 chr3 98837064 N chr3 98837191 N DUP 11
SRR1766476.8245657 chr3 98836982 N chr3 98837208 N DUP 5
SRR1766453.6517158 chr3 98836976 N chr3 98837202 N DUP 5
SRR1766474.10223131 chr3 98836936 N chr3 98837211 N DUP 15
SRR1766462.1485448 chr3 98836936 N chr3 98837211 N DUP 22
SRR1766474.7634086 chr3 98836936 N chr3 98837211 N DUP 22
SRR1766473.10389319 chr3 98836936 N chr3 98837211 N DUP 22
SRR1766444.1499261 chr3 98836932 N chr3 98837256 N DUP 5
SRR1766458.7059989 chr3 98836967 N chr3 98837242 N DUP 10
SRR1766486.10435513 chr3 98836936 N chr3 98837211 N DUP 28
SRR1766486.3612641 chr3 98836940 N chr3 98837264 N DUP 5
SRR1766477.7862590 chr3 98836932 N chr3 98837256 N DUP 5
SRR1766468.6271492 chr3 98836932 N chr3 98837256 N DUP 5
SRR1766450.4800700 chr11 90155473 N chr11 90155553 N DEL 11
SRR1766442.13480876 chr2 231849126 N chr2 231849256 N DEL 5
SRR1766452.7558339 chr2 231849126 N chr2 231849256 N DEL 5
SRR1766458.2321113 chr2 231849126 N chr2 231849256 N DEL 5
SRR1766464.3696723 chr2 231849126 N chr2 231849256 N DEL 5
SRR1766451.2844129 chr2 231848993 N chr2 231849121 N DUP 10
SRR1766462.10527250 chr2 231849126 N chr2 231849256 N DEL 5
SRR1766453.5278350 chr2 231849128 N chr2 231849258 N DEL 5
SRR1766451.7519367 chr2 231849126 N chr2 231849256 N DEL 5
SRR1766475.1548094 chr2 231849126 N chr2 231849256 N DEL 5
SRR1766467.7577496 chr2 231849126 N chr2 231849256 N DEL 10
SRR1766478.3148213 chr2 231849126 N chr2 231849256 N DEL 10
SRR1766484.39213 chr2 231849159 N chr2 231849289 N DEL 5
SRR1766459.6088788 chr2 231849128 N chr2 231849258 N DEL 5
SRR1766453.3894449 chr2 231849126 N chr2 231849256 N DEL 5
SRR1766473.5973136 chr2 231849060 N chr2 231849188 N DUP 8
SRR1766445.8053166 chr2 231848976 N chr2 231849233 N DUP 10
SRR1766445.10466169 chr2 231849142 N chr2 231849270 N DUP 5
SRR1766462.9641635 chr2 231849142 N chr2 231849270 N DUP 5
SRR1766479.1756897 chr2 231849077 N chr2 231849205 N DUP 6
SRR1766461.1869900 chr2 231849077 N chr2 231849205 N DUP 8
SRR1766484.9262232 chr2 231849172 N chr2 231849300 N DUP 4
SRR1766448.6792094 chr2 231849172 N chr2 231849300 N DUP 5
SRR1766474.4642781 chr2 231849172 N chr2 231849300 N DUP 5
SRR1766469.5750749 chr2 231849172 N chr2 231849300 N DUP 5
SRR1766479.12617993 chr2 231849172 N chr2 231849300 N DUP 5
SRR1766451.2281395 chr2 231849172 N chr2 231849300 N DUP 5
SRR1766463.10364656 chr2 231849174 N chr2 231849302 N DUP 5
SRR1766465.5662069 chr2 231849172 N chr2 231849300 N DUP 5
SRR1766459.10577449 chr5 75271140 N chr5 75271283 N DEL 8
SRR1766467.11522837 chr5 75271287 N chr5 75271411 N DUP 5
SRR1766459.1398121 chr5 75271292 N chr5 75271467 N DEL 2
SRR1766473.1771032 chr5 75271251 N chr5 75271425 N DUP 4
SRR1766451.3582536 chr5 75271095 N chr5 75271459 N DUP 2
SRR1766465.8473923 chr5 75271095 N chr5 75271459 N DUP 3
SRR1766476.9980496 chr5 75271095 N chr5 75271459 N DUP 3
SRR1766453.456379 chr5 75271110 N chr5 75271474 N DUP 5
SRR1766486.4604579 chr5 75271162 N chr5 75271477 N DUP 5
SRR1766481.4689109 chr5 75271162 N chr5 75271477 N DUP 5
SRR1766455.1530288 chr5 75271162 N chr5 75271477 N DUP 5
SRR1766456.3310542 chr5 75271283 N chr5 75271456 N DUP 3
SRR1766457.4151586 chr5 75271152 N chr5 75271420 N DEL 4
SRR1766468.6401342 chr5 75271152 N chr5 75271420 N DEL 4
SRR1766464.2401068 chr5 75271155 N chr5 75271423 N DEL 1
SRR1766457.7277840 chr5 75271153 N chr5 75271421 N DEL 3
SRR1766465.7494245 chr5 75271126 N chr5 75271568 N DUP 5
SRR1766466.3658041 chr5 75271124 N chr5 75271490 N DEL 5
SRR1766480.8464335 chr5 75271124 N chr5 75271490 N DEL 5
SRR1766456.4293555 chr5 75271124 N chr5 75271490 N DEL 5
SRR1766455.2557253 chr5 75271474 N chr5 75271602 N DEL 7
SRR1766478.7428368 chr5 75271409 N chr5 75271683 N DEL 9
SRR1766455.4331604 chr5 75271495 N chr5 75271721 N DEL 5
SRR1766461.5230068 chr5 75271144 N chr5 75271686 N DEL 1
SRR1766450.851328 chr5 75271408 N chr5 75271682 N DEL 5
SRR1766463.4557650 chr5 75271115 N chr5 75271706 N DEL 5
SRR1766477.5630875 chr5 75271190 N chr5 75271732 N DEL 4
SRR1766484.3077561 chr7 74053816 N chr7 74053933 N DEL 10
SRR1766443.7088162 chr13 79373320 N chr13 79373438 N DUP 3
SRR1766472.7457313 chr13 79373361 N chr13 79373571 N DUP 8
SRR1766460.1834256 chr13 79373475 N chr13 79373577 N DUP 9
SRR1766456.586782 chr13 79373475 N chr13 79373577 N DUP 9
SRR1766473.3060644 chr21 41067146 N chr21 41067322 N DEL 5
SRR1766481.5555981 chr21 41067146 N chr21 41067322 N DEL 5
SRR1766453.8992478 chr10 57693297 N chr10 57693358 N DEL 1
SRR1766485.9361892 chr10 57693297 N chr10 57693358 N DEL 1
SRR1766477.8262502 chr10 57693307 N chr10 57693432 N DEL 8
SRR1766454.6137218 chr10 57693307 N chr10 57693432 N DEL 9
SRR1766481.10157706 chr10 57693307 N chr10 57693432 N DEL 9
SRR1766458.584918 chr10 57693307 N chr10 57693432 N DEL 11
SRR1766470.3343466 chr10 57693309 N chr10 57693476 N DEL 12
SRR1766442.38684814 chr10 57693309 N chr10 57693532 N DEL 12
SRR1766474.2405713 chr10 57693309 N chr10 57693532 N DEL 12
SRR1766481.12121069 chr10 57693309 N chr10 57693476 N DEL 19
SRR1766471.10267820 chr10 57693307 N chr10 57693432 N DEL 15
SRR1766466.8655538 chr10 57693307 N chr10 57693432 N DEL 15
SRR1766462.809999 chr10 57693309 N chr10 57693476 N DEL 29
SRR1766486.7915736 chr10 57693144 N chr10 57693431 N DUP 5
SRR1766448.3340831 chr10 57693340 N chr10 57693461 N DUP 5
SRR1766461.5797581 chr10 57693340 N chr10 57693461 N DUP 5
SRR1766481.10157706 chr10 57693340 N chr10 57693461 N DUP 5
SRR1766452.8626167 chr10 57693367 N chr10 57693464 N DUP 6
SRR1766442.24046244 chr10 57693367 N chr10 57693464 N DUP 7
SRR1766442.17174949 chr10 57693367 N chr10 57693464 N DUP 8
SRR1766461.2747020 chr10 57693403 N chr10 57693470 N DUP 32
SRR1766448.1181766 chr10 57693310 N chr10 57693465 N DUP 12
SRR1766476.3000853 chr10 57693403 N chr10 57693470 N DUP 29
SRR1766445.8409272 chr10 57693310 N chr10 57693465 N DUP 13
SRR1766448.10139971 chr10 57693310 N chr10 57693465 N DUP 13
SRR1766459.6753269 chr10 57693403 N chr10 57693470 N DUP 26
SRR1766442.37999359 chr10 57693403 N chr10 57693470 N DUP 24
SRR1766442.38955487 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766464.8804941 chr10 57693406 N chr10 57693481 N DUP 2
SRR1766449.6539435 chr10 57693407 N chr10 57693482 N DUP 3
SRR1766472.8923067 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766477.4716957 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766453.5385784 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766455.1778743 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766448.9008293 chr10 57693434 N chr10 57693573 N DUP 24
SRR1766445.4809961 chr10 57693431 N chr10 57693532 N DEL 8
SRR1766444.2235050 chr10 57693434 N chr10 57693573 N DUP 21
SRR1766456.139808 chr10 57693408 N chr10 57693521 N DUP 11
SRR1766444.4056279 chr10 57693150 N chr10 57693419 N DEL 6
SRR1766444.4934318 chr10 57693403 N chr10 57693470 N DUP 19
SRR1766455.9522319 chr10 57693361 N chr10 57693532 N DEL 8
SRR1766482.3689180 chr10 57693403 N chr10 57693470 N DUP 32
SRR1766451.1700638 chr10 57693403 N chr10 57693470 N DUP 29
SRR1766453.8106407 chr10 57693403 N chr10 57693470 N DUP 29
SRR1766466.8902659 chr10 57693403 N chr10 57693470 N DUP 25
SRR1766483.9385623 chr10 57693434 N chr10 57693559 N DUP 21
SRR1766470.9922797 chr10 57693434 N chr10 57693559 N DUP 20
SRR1766463.2489223 chr10 57693434 N chr10 57693559 N DUP 20
SRR1766483.5544864 chr10 57693434 N chr10 57693559 N DUP 20
SRR1766450.7308757 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766454.6116447 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766442.38955487 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766443.2421400 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766464.10894326 chr10 57693489 N chr10 57693613 N DUP 15
SRR1766468.3716087 chr10 57693472 N chr10 57693624 N DUP 11
SRR1766446.10530166 chr10 57693472 N chr10 57693624 N DUP 17
SRR1766444.4056279 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766463.10909858 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766482.3562229 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766465.1035677 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766457.1363229 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766461.552479 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766448.3340831 chr10 57693472 N chr10 57693624 N DUP 20
SRR1766442.33924965 chr10 57693472 N chr10 57693555 N DUP 19
SRR1766453.8992478 chr10 57693476 N chr10 57693628 N DUP 23
SRR1766443.1159957 chr10 57693472 N chr10 57693555 N DUP 24
SRR1766467.6641138 chr10 57693565 N chr10 57693737 N DEL 41
SRR1766459.204497 chr10 57693565 N chr10 57693737 N DEL 38
SRR1766454.7021792 chr10 57693302 N chr10 57693782 N DUP 2
SRR1766474.3338522 chr10 57693472 N chr10 57693555 N DUP 15
SRR1766470.4773511 chr10 57693537 N chr10 57693737 N DEL 38
SRR1766444.6954974 chr10 57693537 N chr10 57693737 N DEL 38
SRR1766461.2747020 chr10 57693537 N chr10 57693737 N DEL 38
SRR1766484.1893741 chr10 57693537 N chr10 57693737 N DEL 38
SRR1766442.17174949 chr10 57693537 N chr10 57693737 N DEL 37
SRR1766459.4757208 chr10 57693370 N chr10 57693698 N DEL 5
SRR1766475.4260971 chr10 57693370 N chr10 57693698 N DEL 5
SRR1766447.5193368 chr10 57693370 N chr10 57693698 N DEL 5
SRR1766463.2226648 chr10 57693537 N chr10 57693737 N DEL 33
SRR1766483.2455630 chr10 57693370 N chr10 57693698 N DEL 5
SRR1766465.8918817 chr10 57693370 N chr10 57693698 N DEL 5
SRR1766455.9614973 chr10 57693370 N chr10 57693698 N DEL 5
SRR1766448.10391787 chr10 57693370 N chr10 57693698 N DEL 5
SRR1766467.52779 chr10 57693537 N chr10 57693737 N DEL 33
SRR1766447.3931403 chr10 57693509 N chr10 57693737 N DEL 33
SRR1766449.2646646 chr10 57693642 N chr10 57693699 N DEL 5
SRR1766466.11331347 chr10 57693642 N chr10 57693699 N DEL 5
SRR1766483.4020392 chr10 57693509 N chr10 57693737 N DEL 33
SRR1766476.9397200 chr10 57693266 N chr10 57693704 N DEL 5
SRR1766481.9163505 chr10 57693648 N chr10 57693705 N DEL 5
SRR1766448.3603075 chr10 57693363 N chr10 57693737 N DEL 20
SRR1766443.2564668 chr10 57693367 N chr10 57693741 N DEL 11
SRR1766475.2287867 chr10 57693365 N chr10 57693739 N DEL 13
SRR1766459.7905286 chr17 60872551 N chr17 60872658 N DUP 5
SRR1766445.5157270 chr10 1232648 N chr10 1232855 N DEL 2
SRR1766468.986778 chr10 1232682 N chr10 1232741 N DUP 2
SRR1766463.8745275 chr10 1232482 N chr10 1232758 N DUP 10
SRR1766447.7776301 chr10 1232664 N chr10 1232871 N DUP 9
SRR1766446.10585390 chr10 1232664 N chr10 1232871 N DUP 9
SRR1766457.5816053 chr10 1232590 N chr10 1232798 N DUP 5
SRR1766476.3883801 chr10 1232903 N chr10 1233021 N DUP 2
SRR1766480.3029218 chr10 1232904 N chr10 1233022 N DUP 1
SRR1766480.3496822 chr10 1232904 N chr10 1233022 N DUP 1
SRR1766451.6527638 chr10 1232788 N chr10 1232982 N DEL 8
SRR1766451.4993401 chr10 1232879 N chr10 1233017 N DEL 5
SRR1766468.2154801 chr10 1232730 N chr10 1233051 N DEL 5
SRR1766448.10161218 chr12 415452 N chr12 415509 N DEL 11
SRR1766443.3688781 chr12 415452 N chr12 415509 N DEL 11
SRR1766446.4119324 chr12 415452 N chr12 415509 N DEL 11
SRR1766471.4878746 chr12 415435 N chr12 415511 N DEL 3
SRR1766459.6340972 chr12 415564 N chr12 415667 N DEL 5
SRR1766466.5529062 chr12 415565 N chr12 415668 N DEL 5
SRR1766479.2234991 chr10 5052906 N chr10 5053065 N DUP 5
SRR1766448.8377879 chr10 5052906 N chr10 5053065 N DUP 5
SRR1766452.4670150 chr10 133028342 N chr10 133028715 N DEL 13
SRR1766445.6261680 chr10 133028432 N chr10 133028669 N DEL 8
SRR1766462.211532 chr10 133028371 N chr10 133028440 N DEL 5
SRR1766454.6476065 chr10 133028562 N chr10 133028715 N DEL 16
SRR1766466.8830080 chr10 133028636 N chr10 133028721 N DEL 13
SRR1766459.2726208 chr10 133028364 N chr10 133028549 N DEL 3
SRR1766458.166845 chr10 133028583 N chr10 133028834 N DUP 5
SRR1766447.2676565 chr10 133028560 N chr10 133028801 N DEL 5
SRR1766455.1258773 chr10 133028617 N chr10 133028802 N DEL 9
SRR1766442.2026185 chr10 133028374 N chr10 133028811 N DEL 5
SRR1766444.253104 chr17 2226520 N chr17 2226837 N DEL 43
SRR1766482.3528281 chr17 2226162 N chr17 2226755 N DUP 5
SRR1766485.1927755 chr17 2226440 N chr17 2226762 N DEL 3
SRR1766442.44515151 chr17 2226176 N chr17 2226771 N DEL 4
SRR1766486.1825734 chr6 135380069 N chr6 135380179 N DUP 1
SRR1766459.8192040 chr3 152771089 N chr3 152771160 N DEL 7
SRR1766465.4287048 chr3 152771087 N chr3 152771160 N DEL 8
SRR1766467.10338942 chr3 152771088 N chr3 152771161 N DEL 7
SRR1766470.9776822 chr3 152771089 N chr3 152771160 N DEL 6
SRR1766444.1978174 chr3 152771107 N chr3 152771162 N DEL 5
SRR1766453.2150620 chr3 152771111 N chr3 152771166 N DEL 5
SRR1766444.5670414 chr19 19770126 N chr19 19770360 N DEL 11
SRR1766482.3884564 chr19 19770075 N chr19 19770190 N DUP 1
SRR1766447.10080043 chr19 19770112 N chr19 19770229 N DEL 5
SRR1766452.2090012 chr8 93666164 N chr8 93666243 N DEL 21
SRR1766443.10105430 chr8 93666170 N chr8 93666249 N DEL 5
SRR1766455.8616820 chr6 58259507 N chr6 58259961 N DUP 1
SRR1766486.10669182 chr6 58259963 N chr6 58261176 N DEL 5
SRR1766453.10608631 chr6 58259963 N chr6 58261176 N DEL 5
SRR1766463.10312002 chr6 58259983 N chr6 58261194 N DUP 5
SRR1766464.728369 chr6 58259985 N chr6 58261196 N DUP 5
SRR1766475.11450876 chr20 50452230 N chr20 50452296 N DEL 1
SRR1766442.29455733 chr20 50452230 N chr20 50452292 N DEL 5
SRR1766481.12202291 chr20 50452230 N chr20 50452292 N DEL 6
SRR1766462.10877049 chr20 50452230 N chr20 50452292 N DEL 8
SRR1766472.8731080 chr9 129576539 N chr9 129576630 N DUP 1
SRR1766475.4962381 chr18 47982686 N chr18 47982961 N DUP 11
SRR1766480.886026 chr18 47982842 N chr18 47982909 N DEL 29
SRR1766448.2953746 chr18 47982879 N chr18 47982932 N DEL 10
SRR1766445.9014445 chr18 47982842 N chr18 47982923 N DEL 8
SRR1766480.6140780 chr18 47982870 N chr18 47982939 N DEL 5
SRR1766451.6098112 chr18 47982872 N chr18 47982941 N DEL 3
SRR1766453.9095276 chr18 47982847 N chr18 47982942 N DEL 2
SRR1766478.8680833 chrX 153382734 N chrX 153382897 N DUP 15
SRR1766466.6338636 chrX 153382712 N chrX 153382858 N DEL 5
SRR1766457.1764064 chrX 153382865 N chrX 153382968 N DUP 6
SRR1766472.1263479 chrX 153382880 N chrX 153382940 N DUP 5
SRR1766480.3949124 chr13 29492009 N chr13 29492060 N DUP 2
SRR1766476.7371967 chr13 29492025 N chr13 29492138 N DUP 5
SRR1766473.9798208 chr13 29492020 N chr13 29492158 N DUP 5
SRR1766485.10128058 chr13 29491974 N chr13 29492158 N DUP 3
SRR1766442.2631460 chr13 29492157 N chr13 29492280 N DEL 1
SRR1766467.2504130 chr13 29492175 N chr13 29492300 N DEL 8
SRR1766446.10042900 chr13 29492175 N chr13 29492300 N DEL 8
SRR1766459.430459 chr13 29492175 N chr13 29492300 N DEL 13
SRR1766468.2764403 chr13 29492114 N chr13 29492274 N DUP 8
SRR1766461.6057204 chr13 29491989 N chr13 29492171 N DEL 8
SRR1766470.10819057 chr13 29492263 N chr13 29492352 N DEL 6
SRR1766463.5127523 chr13 29492073 N chr13 29492365 N DEL 9
SRR1766442.19180689 chr13 29491961 N chr13 29492368 N DEL 9
SRR1766468.6389248 chr13 29491963 N chr13 29492370 N DEL 8
SRR1766459.1587789 chr13 29492044 N chr13 29492386 N DEL 1
SRR1766448.2514947 chr5 176221689 N chr5 176221850 N DEL 5
SRR1766447.8023820 chr1 17313202 N chr1 17313512 N DUP 9
SRR1766470.10066754 chr1 17313276 N chr1 17313588 N DEL 2
SRR1766481.803067 chr19 46315863 N chr19 46316179 N DUP 4
SRR1766465.11292760 chr11 126214538 N chr11 126214639 N DUP 3
SRR1766451.4029082 chr11 126214538 N chr11 126214645 N DUP 6
SRR1766446.6806400 chr11 126214552 N chr11 126214670 N DEL 5
SRR1766479.849787 chr16 88503535 N chr16 88503612 N DEL 14
SRR1766447.1116039 chr16 88503418 N chr16 88503612 N DEL 11
SRR1766448.7453874 chr16 88503418 N chr16 88503612 N DEL 11
SRR1766446.6629149 chr16 88503352 N chr16 88503624 N DEL 3
SRR1766454.10387899 chr17 513777 N chr17 514376 N DEL 10
SRR1766454.8905852 chr17 513750 N chr17 513841 N DUP 15
SRR1766483.5323667 chr17 513785 N chr17 513876 N DUP 5
SRR1766474.1411407 chr17 513822 N chr17 513913 N DUP 5
SRR1766450.10507364 chr17 513779 N chr17 513872 N DEL 5
SRR1766442.26059876 chr17 513875 N chr17 514058 N DUP 2
SRR1766451.5175205 chr17 513792 N chr17 513885 N DEL 2
SRR1766443.9480016 chr17 513793 N chr17 513886 N DEL 1
SRR1766454.3317024 chr17 513815 N chr17 513908 N DEL 5
SRR1766468.5965867 chr17 513778 N chr17 513917 N DEL 5
SRR1766453.3490162 chr17 513779 N chr17 513918 N DEL 2
SRR1766452.5574745 chr17 513781 N chr17 513920 N DEL 3
SRR1766477.8446947 chr17 513781 N chr17 513920 N DEL 3
SRR1766477.5700713 chr17 513815 N chr17 513908 N DEL 1
SRR1766459.4851646 chr17 513916 N chr17 514375 N DUP 8
SRR1766475.4211247 chr17 513815 N chr17 513908 N DEL 5
SRR1766473.449724 chr17 513822 N chr17 513915 N DEL 5
SRR1766463.9004458 chr17 513815 N chr17 513908 N DEL 5
SRR1766452.5574745 chr17 514000 N chr17 514553 N DEL 15
SRR1766462.6133761 chr17 513815 N chr17 513908 N DEL 5
SRR1766465.7786116 chr17 513815 N chr17 513908 N DEL 5
SRR1766451.6123471 chr17 514008 N chr17 514375 N DUP 5
SRR1766462.293836 chr17 513815 N chr17 514230 N DEL 4
SRR1766460.8809729 chr17 513815 N chr17 514230 N DEL 5
SRR1766455.4603051 chr17 513918 N chr17 514055 N DUP 5
SRR1766449.6367200 chr17 513908 N chr17 514091 N DUP 5
SRR1766474.1411407 chr17 513816 N chr17 514553 N DEL 10
SRR1766442.35057297 chr17 513872 N chr17 514101 N DUP 5
SRR1766464.7266408 chr17 513872 N chr17 514101 N DUP 5
SRR1766482.6382862 chr17 514092 N chr17 514507 N DEL 19
SRR1766444.4244201 chr17 513784 N chr17 514059 N DUP 5
SRR1766459.10019914 chr17 513872 N chr17 514101 N DUP 5
SRR1766442.44866427 chr17 513872 N chr17 514101 N DUP 5
SRR1766442.42990812 chr17 513792 N chr17 514161 N DEL 2
SRR1766462.3947516 chr17 513779 N chr17 513872 N DEL 5
SRR1766484.10769514 chr17 514099 N chr17 514560 N DEL 10
SRR1766449.1996712 chr17 513815 N chr17 514230 N DEL 5
SRR1766484.11434380 chr17 513769 N chr17 514230 N DEL 5
SRR1766485.935551 chr17 513773 N chr17 514234 N DEL 5
SRR1766483.2256060 chr17 513774 N chr17 514235 N DEL 5
SRR1766465.10073698 chr17 514058 N chr17 514243 N DEL 2
SRR1766463.10254058 chr17 513750 N chr17 514347 N DUP 8
SRR1766455.3751661 chr17 513908 N chr17 514091 N DUP 4
SRR1766463.984017 chr17 513872 N chr17 514331 N DUP 10
SRR1766462.1923040 chr17 513815 N chr17 513908 N DEL 5
SRR1766442.3968892 chr17 513815 N chr17 513908 N DEL 5
SRR1766474.628133 chr17 513815 N chr17 513908 N DEL 5
SRR1766459.9807435 chr17 513861 N chr17 514276 N DEL 5
SRR1766459.5800291 chr17 513845 N chr17 514628 N DEL 15
SRR1766485.2648137 chr17 513999 N chr17 514690 N DEL 5
SRR1766459.2743242 chr17 514413 N chr17 514598 N DEL 10
SRR1766458.6279268 chr17 514397 N chr17 514582 N DEL 15
SRR1766460.8809729 chr17 514000 N chr17 514507 N DEL 17
SRR1766465.5874682 chr17 513778 N chr17 514375 N DUP 4
SRR1766454.10387899 chr17 513777 N chr17 514376 N DEL 3
SRR1766450.10471995 chr17 513823 N chr17 514376 N DEL 5
SRR1766444.4244201 chr17 513823 N chr17 514376 N DEL 5
SRR1766483.5323667 chr17 514414 N chr17 514507 N DEL 10
SRR1766456.1210099 chr17 513824 N chr17 514467 N DUP 5
SRR1766454.2335561 chr17 513872 N chr17 514469 N DUP 5
SRR1766469.10663452 chr17 513882 N chr17 514389 N DEL 4
SRR1766465.7786116 chr17 513769 N chr17 514414 N DEL 5
SRR1766471.5622111 chr17 513777 N chr17 514422 N DEL 10
SRR1766484.5300104 chr17 513777 N chr17 514422 N DEL 10
SRR1766443.6384540 chr17 514430 N chr17 514751 N DUP 3
SRR1766478.3338244 chr17 513791 N chr17 514436 N DEL 1
SRR1766451.4955591 chr17 513869 N chr17 514422 N DEL 5
SRR1766475.6312930 chr17 513823 N chr17 514468 N DEL 5
SRR1766483.9072803 chr17 513823 N chr17 514468 N DEL 10
SRR1766481.13060514 chr17 513872 N chr17 514515 N DUP 10
SRR1766464.7266408 chr17 513862 N chr17 514507 N DEL 15
SRR1766459.2533852 chr17 513819 N chr17 514510 N DEL 10
SRR1766482.385766 chr17 513870 N chr17 514469 N DEL 5
SRR1766477.5700713 chr17 513862 N chr17 514507 N DEL 5
SRR1766454.8724154 chr17 513865 N chr17 514510 N DEL 5
SRR1766461.6691777 chr17 513815 N chr17 514506 N DEL 10
SRR1766475.4211247 chr17 513862 N chr17 514553 N DEL 5
SRR1766463.9004458 chr17 513862 N chr17 514553 N DEL 5
SRR1766482.12692664 chr17 513815 N chr17 514552 N DEL 5
SRR1766448.2229688 chr17 513815 N chr17 514552 N DEL 5
SRR1766454.8905852 chr17 513862 N chr17 514553 N DEL 5
SRR1766449.6367200 chr17 513799 N chr17 514582 N DEL 13
SRR1766480.8419087 chr17 513868 N chr17 514559 N DEL 5
SRR1766445.1350308 chr17 513954 N chr17 514599 N DEL 15
SRR1766446.3837643 chr17 513799 N chr17 514582 N DEL 5
SRR1766445.10318933 chr17 514000 N chr17 514645 N DEL 10
SRR1766472.7532989 chr17 513845 N chr17 514628 N DEL 10
SRR1766469.2039799 chr17 513803 N chr17 514586 N DEL 5
SRR1766481.2543704 chr17 513803 N chr17 514586 N DEL 5
SRR1766457.1835406 chr17 513770 N chr17 514599 N DEL 6
SRR1766442.31045508 chr17 513816 N chr17 514645 N DEL 5
SRR1766442.35057297 chr17 513782 N chr17 514611 N DEL 3
SRR1766464.4877394 chr17 513799 N chr17 514628 N DEL 5
SRR1766483.11594712 chr17 513801 N chr17 514630 N DEL 5
SRR1766465.7549356 chr17 513999 N chr17 514690 N DEL 7
SRR1766447.9491750 chr17 513799 N chr17 514674 N DEL 10
SRR1766469.6300760 chr17 513783 N chr17 514658 N DEL 2
SRR1766475.2143380 chr17 513799 N chr17 514674 N DEL 7
SRR1766442.3968892 chr17 513799 N chr17 514674 N DEL 5
SRR1766480.2269130 chr17 513812 N chr17 514687 N DEL 2
SRR1766460.1183346 chr17 513823 N chr17 514698 N DEL 11
SRR1766481.9768781 chr17 513789 N chr17 514710 N DEL 3
SRR1766464.2936417 chr2 238633837 N chr2 238633948 N DUP 5
SRR1766462.3455551 chr2 238633828 N chr2 238633999 N DEL 5
SRR1766458.5901849 chr2 238633800 N chr2 238634029 N DEL 21
SRR1766486.3899436 chr7 44307133 N chr7 44307194 N DEL 13
SRR1766442.34312181 chr7 44307129 N chr7 44307228 N DUP 7
SRR1766442.8726266 chr7 44307047 N chr7 44307145 N DEL 7
SRR1766446.1588920 chr7 44307067 N chr7 44307305 N DEL 5
SRR1766483.6994981 chr7 44307045 N chr7 44307377 N DEL 13
SRR1766470.6803338 chr7 44306887 N chr7 44307377 N DEL 15
SRR1766452.5885207 chr7 44306910 N chr7 44307380 N DEL 7
SRR1766478.1203600 chr7 44307316 N chr7 44307574 N DEL 20
SRR1766457.8515746 chr17 83096612 N chr17 83096684 N DEL 5
SRR1766444.2455469 chr17 83096462 N chr17 83096527 N DEL 2
SRR1766482.12214927 chr5 107848382 N chr5 107848486 N DEL 2
SRR1766479.12574162 chr5 107848382 N chr5 107848486 N DEL 5
SRR1766454.5413134 chr5 107848382 N chr5 107848486 N DEL 5
SRR1766442.10076471 chr5 107848382 N chr5 107848486 N DEL 5
SRR1766469.1286618 chr5 107848382 N chr5 107848486 N DEL 5
SRR1766466.9248054 chr5 107848382 N chr5 107848486 N DEL 5
SRR1766476.5876239 chr5 107848382 N chr5 107848486 N DEL 15
SRR1766469.3822872 chr5 107848382 N chr5 107848486 N DEL 19
SRR1766466.8029342 chr5 107848396 N chr5 107848500 N DEL 1
SRR1766472.3807926 chr5 107848394 N chr5 107848498 N DEL 3
SRR1766442.32605927 chr20 18010549 N chr20 18010675 N DUP 5
SRR1766467.670610 chr20 18010549 N chr20 18010675 N DUP 5
SRR1766472.3180621 chr20 18010598 N chr20 18010894 N DUP 1
SRR1766466.7039552 chr20 18010659 N chr20 18010740 N DUP 5
SRR1766442.17515044 chr20 18010659 N chr20 18010740 N DUP 15
SRR1766475.10891209 chr20 18010522 N chr20 18010779 N DUP 5
SRR1766456.1385979 chr20 18010700 N chr20 18010832 N DEL 6
SRR1766442.17515044 chr20 18010526 N chr20 18010834 N DEL 5
SRR1766442.16712989 chr20 18010616 N chr20 18010952 N DUP 6
SRR1766463.10108778 chr8 19450247 N chr8 19450302 N DEL 12
SRR1766467.10414418 chr5 173285163 N chr5 173285315 N DEL 10
SRR1766474.3753932 chr17 7176592 N chr17 7176655 N DUP 5
SRR1766465.6205749 chr17 7176591 N chr17 7176654 N DUP 10
SRR1766454.8745468 chr3 186601242 N chr3 186601308 N DEL 5
SRR1766478.8704995 chr3 127155508 N chr3 127155625 N DUP 5
SRR1766469.7798101 chr3 127155515 N chr3 127155660 N DUP 2
SRR1766472.1748152 chr3 127155570 N chr3 127155715 N DUP 4
SRR1766467.8649616 chr3 127155601 N chr3 127155752 N DUP 10
SRR1766455.1926442 chr3 127155489 N chr3 127155608 N DEL 8
SRR1766442.29960524 chr3 127155683 N chr3 127155940 N DUP 7
SRR1766448.2660735 chr3 127155683 N chr3 127155940 N DUP 7
SRR1766470.6920485 chr3 127155606 N chr3 127155681 N DEL 5
SRR1766471.6741755 chr3 127155489 N chr3 127155688 N DEL 4
SRR1766468.6727884 chr3 127155498 N chr3 127155823 N DEL 5
SRR1766459.2930480 chr3 127155611 N chr3 127155950 N DUP 7
SRR1766442.33477466 chr3 127155611 N chr3 127155950 N DUP 7
SRR1766453.6138675 chr3 127155611 N chr3 127155950 N DUP 7
SRR1766466.8716389 chr3 127155684 N chr3 127155987 N DUP 1
SRR1766470.5499107 chr3 127155684 N chr3 127155987 N DUP 1
SRR1766461.1455748 chr3 127155623 N chr3 127155916 N DEL 15
SRR1766450.5495346 chr3 127155667 N chr3 127156008 N DUP 10
SRR1766475.7255746 chr1 203781623 N chr1 203781917 N DEL 7
SRR1766483.4033470 chr1 203781624 N chr1 203781927 N DEL 5
SRR1766466.586415 chr1 203781623 N chr1 203781935 N DEL 5
SRR1766471.3912925 chr1 203781660 N chr1 203781969 N DEL 19
SRR1766463.8995767 chr14 86375742 N chr14 86375805 N DUP 5
SRR1766453.10917641 chr7 35682375 N chr7 35682514 N DEL 9
SRR1766443.2384811 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766473.2096586 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766482.10072918 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766469.6508093 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766463.5237044 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766477.1504889 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766469.3245033 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766478.7659731 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766477.10718684 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766442.25599103 chr8 1565024 N chr8 1565103 N DUP 5
SRR1766479.1976983 chr4 3567125 N chr4 3567237 N DUP 1
SRR1766442.1726989 chr4 3567125 N chr4 3567237 N DUP 2
SRR1766467.2978202 chr4 3567125 N chr4 3567237 N DUP 5
SRR1766464.528150 chr4 3567123 N chr4 3567235 N DUP 10
SRR1766478.7053797 chr4 3567123 N chr4 3567235 N DUP 5
SRR1766452.8932261 chr4 3567106 N chr4 3567268 N DUP 5
SRR1766453.8707988 chr4 3567190 N chr4 3567273 N DUP 5
SRR1766451.3815947 chr4 3567106 N chr4 3567268 N DUP 5
SRR1766447.5758201 chr4 3567227 N chr4 3567355 N DUP 5
SRR1766463.4664916 chr4 3567143 N chr4 3567257 N DEL 5
SRR1766463.5329350 chr1 194303974 N chr1 194304045 N DUP 30
SRR1766477.11461267 chr1 194303954 N chr1 194304032 N DUP 18
SRR1766485.7707537 chr1 194303954 N chr1 194304032 N DUP 16
SRR1766474.4138833 chr1 194303974 N chr1 194304045 N DUP 27
SRR1766481.358894 chr1 194303954 N chr1 194304032 N DUP 14
SRR1766461.3794238 chr1 194303974 N chr1 194304045 N DUP 25
SRR1766443.621635 chr1 194303954 N chr1 194304032 N DUP 10
SRR1766446.2074640 chr1 194303974 N chr1 194304045 N DUP 22
SRR1766442.33491480 chr1 194303974 N chr1 194304045 N DUP 22
SRR1766474.5845751 chr1 194303954 N chr1 194304032 N DUP 10
SRR1766480.4817582 chr1 194303954 N chr1 194304032 N DUP 10
SRR1766455.5540420 chr1 194303954 N chr1 194304032 N DUP 10
SRR1766484.11718702 chr1 194303979 N chr1 194304085 N DUP 24
SRR1766477.3912043 chr1 194303974 N chr1 194304045 N DUP 22
SRR1766458.2713721 chr1 194303979 N chr1 194304085 N DUP 21
SRR1766483.2815842 chr1 194303979 N chr1 194304052 N DUP 12
SRR1766482.12070223 chr1 194303978 N chr1 194304088 N DUP 7
SRR1766471.1897321 chr1 194303979 N chr1 194304085 N DUP 21
SRR1766452.9978218 chr1 194303979 N chr1 194304085 N DUP 15
SRR1766457.9333976 chr1 194303978 N chr1 194304088 N DUP 9
SRR1766454.3881683 chr1 194303979 N chr1 194304085 N DUP 17
SRR1766459.9659730 chr1 194303974 N chr1 194304084 N DUP 11
SRR1766462.10934262 chr1 194303979 N chr1 194304085 N DUP 24
SRR1766467.8135243 chr1 194303979 N chr1 194304089 N DUP 10
SRR1766483.6270725 chr1 194303981 N chr1 194304087 N DUP 24
SRR1766463.9385861 chr1 194303954 N chr1 194304069 N DUP 16
SRR1766486.9315120 chr1 194303992 N chr1 194304065 N DUP 8
SRR1766457.753364 chr1 194303975 N chr1 194304048 N DUP 9
SRR1766470.3088814 chr1 194303975 N chr1 194304048 N DUP 9
SRR1766465.3065002 chr1 194303994 N chr1 194304067 N DUP 5
SRR1766466.9430200 chr1 194303974 N chr1 194304045 N DUP 27
SRR1766462.10318776 chr1 194303979 N chr1 194304085 N DUP 26
SRR1766478.8008826 chr1 194303979 N chr1 194304085 N DUP 27
SRR1766445.2556709 chr1 194303979 N chr1 194304052 N DUP 14
SRR1766457.7419715 chr1 194303979 N chr1 194304052 N DUP 15
SRR1766472.5164348 chr1 194303979 N chr1 194304052 N DUP 11
SRR1766479.11822420 chr1 194303937 N chr1 194304098 N DEL 11
SRR1766454.9385242 chr1 194303938 N chr1 194304099 N DEL 10
SRR1766476.2767915 chr13 28633898 N chr13 28634000 N DEL 7
SRR1766481.9867576 chr13 28633898 N chr13 28634000 N DEL 7
SRR1766455.9576174 chr13 28633900 N chr13 28634002 N DEL 7
SRR1766485.5453651 chr13 28633902 N chr13 28634004 N DEL 7
SRR1766481.472272 chr13 28633904 N chr13 28634006 N DEL 7
SRR1766476.6048187 chr13 28633813 N chr13 28634009 N DEL 6
SRR1766447.10467825 chr13 28633815 N chr13 28634011 N DEL 4
SRR1766447.8440982 chr15 99538171 N chr15 99538231 N DUP 4
SRR1766456.3353895 chr15 99538164 N chr15 99538229 N DUP 12
SRR1766453.9802769 chr15 99538164 N chr15 99538234 N DUP 30
SRR1766462.9418870 chr15 99538204 N chr15 99538331 N DUP 9
SRR1766471.7649534 chr15 99538217 N chr15 99538328 N DUP 17
SRR1766448.7118808 chr15 99538185 N chr15 99538242 N DEL 5
SRR1766450.4295297 chr15 99538185 N chr15 99538278 N DEL 5
SRR1766448.3553206 chr15 99538186 N chr15 99538279 N DEL 5
SRR1766466.3420508 chr15 99538189 N chr15 99538282 N DEL 5
SRR1766456.828408 chr18 39802145 N chr18 39802217 N DEL 8
SRR1766471.2721028 chr1 5821474 N chr1 5821571 N DUP 2
SRR1766469.5507709 chr3 53220693 N chr3 53220768 N DUP 3
SRR1766462.7051149 chr3 53220698 N chr3 53220773 N DUP 10
SRR1766471.8810077 chr3 53220693 N chr3 53220768 N DUP 6
SRR1766473.11161244 chr3 53220693 N chr3 53220768 N DUP 6
SRR1766482.6765648 chr3 53220693 N chr3 53220768 N DUP 7
SRR1766463.7825909 chr3 53220693 N chr3 53220768 N DUP 9
SRR1766450.2468939 chr3 53220693 N chr3 53220768 N DUP 11
SRR1766445.3229622 chr3 53220693 N chr3 53220768 N DUP 11
SRR1766473.10806054 chr3 53220693 N chr3 53220768 N DUP 17
SRR1766455.9494665 chr4 151732108 N chr4 151732201 N DUP 11
SRR1766443.3675115 chr4 151732089 N chr4 151732182 N DUP 5
SRR1766458.356231 chr4 151732092 N chr4 151732185 N DUP 5
SRR1766472.5292795 chr4 151732108 N chr4 151732201 N DUP 6
SRR1766458.356231 chr4 151732084 N chr4 151732177 N DUP 5
SRR1766483.8017323 chr4 151732125 N chr4 151732219 N DUP 14
SRR1766449.5351571 chr4 151732125 N chr4 151732219 N DUP 15
SRR1766473.7014302 chr14 41808350 N chr14 41808476 N DUP 10
SRR1766465.9403511 chr14 41808350 N chr14 41808492 N DUP 5
SRR1766442.37667490 chr14 41808350 N chr14 41808476 N DUP 5
SRR1766447.10229442 chr13 108013563 N chr13 108013653 N DUP 5
SRR1766452.6164498 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766471.697922 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766479.11559321 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766476.222021 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766484.7408776 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766478.338504 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766463.2790873 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766480.7357442 chr3 60860445 N chr3 60860532 N DUP 10
SRR1766485.12066027 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766485.10768909 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766457.6262873 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766458.9287330 chr3 60860467 N chr3 60860532 N DUP 10
SRR1766480.3000600 chr3 60860467 N chr3 60860532 N DUP 7
SRR1766483.11240195 chr3 60860439 N chr3 60860550 N DEL 5
SRR1766442.40836406 chr3 60860439 N chr3 60860550 N DEL 5
SRR1766447.8688072 chr3 60860708 N chr3 60861327 N DEL 6
SRR1766442.15157501 chr3 60860708 N chr3 60861352 N DEL 9
SRR1766445.7457421 chr3 60860708 N chr3 60861352 N DEL 9
SRR1766485.1816155 chr3 60860671 N chr3 60860889 N DEL 9
SRR1766481.3283283 chr3 60860671 N chr3 60860889 N DEL 10
SRR1766483.5993109 chr3 60860671 N chr3 60860889 N DEL 13
SRR1766448.1799644 chr3 60860671 N chr3 60860889 N DEL 14
SRR1766462.4903994 chr3 60860671 N chr3 60860889 N DEL 14
SRR1766471.11733694 chr3 60860671 N chr3 60860889 N DEL 15
SRR1766462.2354933 chr3 60860671 N chr3 60860889 N DEL 15
SRR1766442.15233988 chr3 60860671 N chr3 60860889 N DEL 15
SRR1766442.38204776 chr3 60860671 N chr3 60860889 N DEL 15
SRR1766442.9842272 chr3 60860671 N chr3 60860889 N DEL 9
SRR1766452.75794 chr3 60860671 N chr3 60860889 N DEL 9
SRR1766463.3610676 chr3 60860671 N chr3 60860889 N DEL 9
SRR1766449.1101688 chr3 60860671 N chr3 60860889 N DEL 9
SRR1766485.12066027 chr3 60860671 N chr3 60860889 N DEL 9
SRR1766462.666280 chr3 60860643 N chr3 60860708 N DEL 9
SRR1766466.5425960 chr3 60860645 N chr3 60860710 N DEL 9
SRR1766476.4922483 chr3 60860645 N chr3 60860710 N DEL 9
SRR1766461.9564372 chr3 60860653 N chr3 60860718 N DEL 4
SRR1766471.7923542 chr3 60860888 N chr3 60861013 N DEL 16
SRR1766465.1580462 chr3 60860800 N chr3 60860861 N DUP 12
SRR1766448.1799644 chr3 60860819 N chr3 60860911 N DUP 21
SRR1766477.3672114 chr3 60860955 N chr3 60861327 N DEL 3
SRR1766447.10529974 chr3 60860800 N chr3 60860861 N DUP 2
SRR1766463.4530372 chr3 60860819 N chr3 60860911 N DUP 18
SRR1766451.5226196 chr3 60860911 N chr3 60860976 N DEL 24
SRR1766474.837542 chr3 60860911 N chr3 60860976 N DEL 27
SRR1766462.2354933 chr3 60860911 N chr3 60860976 N DEL 20
SRR1766456.4561025 chr3 60860911 N chr3 60860976 N DEL 13
SRR1766445.3556066 chr3 60860911 N chr3 60860976 N DEL 12
SRR1766451.9911731 chr3 60860911 N chr3 60860976 N DEL 12
SRR1766473.817752 chr3 60860911 N chr3 60860976 N DEL 11
SRR1766442.29031690 chr3 60860976 N chr3 60861370 N DUP 11
SRR1766442.21664132 chr3 60860976 N chr3 60861370 N DUP 10
SRR1766457.1737569 chr3 60860849 N chr3 60861005 N DEL 20
SRR1766463.10281596 chr3 60860787 N chr3 60861004 N DEL 9
SRR1766453.8305262 chr3 60860787 N chr3 60861004 N DEL 9
SRR1766483.12388682 chr3 60861325 N chr3 60861374 N DUP 19
SRR1766443.5382570 chr3 60861325 N chr3 60861374 N DUP 23
SRR1766484.5797667 chr3 60861331 N chr3 60861397 N DUP 13
SRR1766460.997619 chr3 60861331 N chr3 60861397 N DUP 14
SRR1766466.5425960 chr3 60861331 N chr3 60861397 N DUP 15
SRR1766469.4226798 chr3 60861325 N chr3 60861374 N DUP 15
SRR1766449.1972374 chr3 60861363 N chr3 60861418 N DUP 45
SRR1766454.867446 chr3 60861363 N chr3 60861418 N DUP 49
SRR1766442.31422660 chr3 60861363 N chr3 60861418 N DUP 50
SRR1766464.1820646 chr3 60861363 N chr3 60861418 N DUP 50
SRR1766476.518582 chr3 60861363 N chr3 60861418 N DUP 43
SRR1766472.4426684 chr3 60861363 N chr3 60861418 N DUP 32
SRR1766475.7945408 chr3 60861363 N chr3 60861418 N DUP 30
SRR1766462.5828437 chr3 60861363 N chr3 60861418 N DUP 30
SRR1766442.179443 chr3 60861339 N chr3 60861402 N DEL 9
SRR1766449.6707718 chr3 60861338 N chr3 60861410 N DEL 5
SRR1766459.9083631 chr3 60861340 N chr3 60861412 N DEL 5
SRR1766448.2603475 chr8 92949820 N chr8 92949935 N DEL 1
SRR1766461.7446069 chr8 92949737 N chr8 92949832 N DUP 5
SRR1766454.8399615 chr8 92949696 N chr8 92949789 N DEL 1
SRR1766442.44601420 chr8 92949822 N chr8 92949931 N DUP 1
SRR1766479.12526102 chr8 92949831 N chr8 92949944 N DEL 17
SRR1766442.12497524 chr8 92949831 N chr8 92949940 N DEL 13
SRR1766456.15467 chr8 92949831 N chr8 92949940 N DEL 13
SRR1766471.7744362 chr8 92949831 N chr8 92949944 N DEL 17
SRR1766459.281501 chr8 92949831 N chr8 92949944 N DEL 17
SRR1766483.8249271 chr8 92949831 N chr8 92949940 N DEL 13
SRR1766442.1491400 chr8 92949831 N chr8 92949944 N DEL 17
SRR1766482.12930706 chr8 92949831 N chr8 92949940 N DEL 13
SRR1766442.26922800 chr8 92949950 N chr8 92950062 N DUP 12
SRR1766449.4978335 chr8 92949679 N chr8 92949950 N DEL 5
SRR1766460.6231183 chr8 92949679 N chr8 92949954 N DEL 5
SRR1766461.5403136 chr3 60553589 N chr3 60553645 N DUP 9
SRR1766471.4246382 chr3 60553589 N chr3 60553645 N DUP 9
SRR1766454.8041048 chr9 137346675 N chr9 137346755 N DUP 3
SRR1766449.6914977 chr9 137346675 N chr9 137346755 N DUP 5
SRR1766467.5683003 chr9 137346675 N chr9 137346755 N DUP 5
SRR1766465.3998335 chr9 137346675 N chr9 137346755 N DUP 6
SRR1766477.5342213 chr9 137346675 N chr9 137346755 N DUP 7
SRR1766442.5990419 chr9 137346675 N chr9 137346755 N DUP 7
SRR1766463.9811517 chr9 137346675 N chr9 137346755 N DUP 7
SRR1766467.553454 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766454.3934622 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766452.5436474 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766470.2893510 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766462.3998730 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766464.709182 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766448.630881 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766442.44025291 chr9 137346675 N chr9 137346755 N DUP 12
SRR1766466.5871898 chr9 137346675 N chr9 137346755 N DUP 15
SRR1766442.9207384 chr9 137346675 N chr9 137346755 N DUP 15
SRR1766452.5061677 chr9 137346675 N chr9 137346755 N DUP 17
SRR1766459.11523964 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766465.485204 chr9 137346675 N chr9 137346755 N DUP 14
SRR1766465.8611863 chr9 137346675 N chr9 137346755 N DUP 16
SRR1766473.438832 chr9 137346675 N chr9 137346755 N DUP 18
SRR1766453.649293 chr9 137346677 N chr9 137346757 N DUP 5
SRR1766458.8534101 chr9 137346679 N chr9 137346759 N DUP 5
SRR1766451.3158204 chr9 137346675 N chr9 137346755 N DUP 10
SRR1766450.9886743 chr9 137346675 N chr9 137346755 N DUP 11
SRR1766482.6846727 chr9 137346686 N chr9 137346766 N DUP 4
SRR1766486.1270104 chr9 137346675 N chr9 137346755 N DUP 17
SRR1766477.4644375 chr9 137346675 N chr9 137346755 N DUP 18
SRR1766478.6821376 chr9 137346675 N chr9 137346755 N DUP 25
SRR1766482.9248942 chr9 137346675 N chr9 137346755 N DUP 29
SRR1766456.5732290 chr9 137346675 N chr9 137346755 N DUP 31
SRR1766449.1322370 chr9 137346675 N chr9 137346755 N DUP 32
SRR1766442.17412559 chr9 137346675 N chr9 137346755 N DUP 34
SRR1766454.3361702 chr17 17486990 N chr17 17487108 N DUP 4
SRR1766471.9901825 chr16 34941880 N chr16 34942237 N DUP 5
SRR1766446.338854 chr16 34941880 N chr16 34942237 N DUP 5
SRR1766484.4039994 chr16 89118061 N chr16 89118387 N DEL 5
SRR1766455.134915 chr16 89118072 N chr16 89118127 N DEL 3
SRR1766467.7578342 chr16 89118184 N chr16 89118237 N DUP 5
SRR1766455.4979907 chr16 89118096 N chr16 89118368 N DEL 10
SRR1766442.29107285 chr1 246783094 N chr1 246783149 N DEL 6
SRR1766444.4345832 chr1 246783143 N chr1 246783198 N DEL 5
SRR1766442.17801777 chr1 246783177 N chr1 246783720 N DEL 5
SRR1766478.855463 chr1 246783161 N chr1 246783272 N DEL 6
SRR1766475.7758344 chr1 246783161 N chr1 246783272 N DEL 7
SRR1766465.11264477 chr1 246783161 N chr1 246783272 N DEL 12
SRR1766461.4373721 chr1 246783161 N chr1 246783272 N DEL 12
SRR1766475.9939127 chr1 246783162 N chr1 246783273 N DEL 5
SRR1766474.6356817 chr1 246783144 N chr1 246783255 N DEL 10
SRR1766486.11441733 chr1 246783143 N chr1 246783254 N DEL 6
SRR1766460.8066768 chr1 246783178 N chr1 246783611 N DUP 5
SRR1766469.2045721 chr1 246783161 N chr1 246783272 N DEL 12
SRR1766447.10432918 chr1 246783109 N chr1 246783274 N DEL 5
SRR1766453.471251 chr1 246783110 N chr1 246783275 N DEL 5
SRR1766478.1149973 chr1 246783124 N chr1 246783611 N DUP 5
SRR1766447.11089647 chr1 246783161 N chr1 246783272 N DEL 12
SRR1766478.1433909 chr1 246783341 N chr1 246783666 N DEL 5
SRR1766472.7305625 chr1 246783161 N chr1 246783542 N DEL 5
SRR1766471.6438661 chr1 246783121 N chr1 246783556 N DEL 1
SRR1766445.3828254 chr1 246783143 N chr1 246783578 N DEL 5
SRR1766450.9647453 chr1 246783185 N chr1 246783672 N DUP 5
SRR1766462.3878972 chr1 246783185 N chr1 246783672 N DUP 5
SRR1766448.4417635 chr1 246783241 N chr1 246783672 N DUP 5
SRR1766451.8627045 chr1 246783211 N chr1 246783646 N DEL 5
SRR1766442.29107285 chr1 246783211 N chr1 246783646 N DEL 5
SRR1766479.11196940 chr1 246783658 N chr1 246783711 N DUP 10
SRR1766462.9745035 chr1 246783284 N chr1 246783663 N DEL 1
SRR1766442.26007885 chr1 246783137 N chr1 246783680 N DEL 6
SRR1766482.12139146 chr1 246783271 N chr1 246783704 N DEL 9
SRR1766442.36133833 chr1 246783215 N chr1 246783704 N DEL 5
SRR1766467.4678479 chr1 246783216 N chr1 246783705 N DEL 5
SRR1766482.10113521 chr1 246783215 N chr1 246783704 N DEL 5
SRR1766442.38142669 chr1 246783216 N chr1 246783705 N DEL 5
SRR1766486.11441733 chr1 246783162 N chr1 246783705 N DEL 5
SRR1766463.9581663 chr1 246783138 N chr1 246783735 N DEL 5
SRR1766468.3913814 chr22 35343026 N chr22 35343145 N DEL 10
SRR1766476.11029581 chr22 35342916 N chr22 35343158 N DUP 4
SRR1766480.607020 chr22 35343029 N chr22 35343148 N DEL 10
SRR1766483.4128890 chr22 35342943 N chr22 35343108 N DUP 10
SRR1766453.4484805 chr22 35342929 N chr22 35343055 N DEL 1
SRR1766465.9205454 chr22 35343132 N chr22 35343609 N DUP 8
SRR1766445.7386224 chr22 35342967 N chr22 35343139 N DEL 1
SRR1766442.37064475 chr22 35342967 N chr22 35343139 N DEL 1
SRR1766449.1467942 chr22 35343255 N chr22 35343475 N DEL 5
SRR1766465.6230714 chr22 35343280 N chr22 35343496 N DEL 1
SRR1766480.3699349 chr22 35343420 N chr22 35343845 N DEL 2
SRR1766477.3325424 chr22 35343423 N chr22 35343886 N DEL 5
SRR1766452.9795082 chr22 35343229 N chr22 35343444 N DUP 3
SRR1766443.5069973 chr22 35343444 N chr22 35343562 N DUP 15
SRR1766475.1516000 chr22 35343444 N chr22 35343562 N DUP 18
SRR1766468.2071797 chr22 35343450 N chr22 35343568 N DUP 8
SRR1766442.9296832 chr22 35342948 N chr22 35343411 N DEL 9
SRR1766464.1006011 chr22 35343353 N chr22 35343471 N DUP 6
SRR1766477.768154 chr22 35343353 N chr22 35343471 N DUP 19
SRR1766450.8110981 chr22 35343484 N chr22 35343668 N DEL 9
SRR1766469.858437 chr22 35343444 N chr22 35343562 N DUP 13
SRR1766442.21849910 chr22 35342940 N chr22 35343520 N DUP 9
SRR1766447.3643589 chr22 35343425 N chr22 35343541 N DUP 2
SRR1766461.9619339 chr22 35343425 N chr22 35343541 N DUP 2
SRR1766443.5069973 chr22 35343425 N chr22 35343541 N DUP 2
SRR1766474.827521 chr22 35343127 N chr22 35343462 N DEL 1
SRR1766448.2499982 chr22 35343125 N chr22 35343460 N DEL 4
SRR1766454.3890269 chr22 35343001 N chr22 35343460 N DEL 2
SRR1766465.6443837 chr22 35343252 N chr22 35343588 N DUP 5
SRR1766479.12844044 chr22 35343222 N chr22 35343632 N DUP 6
SRR1766472.5279979 chr22 35342901 N chr22 35343666 N DUP 5
SRR1766442.14051561 chr22 35343222 N chr22 35343663 N DUP 7
SRR1766451.3378260 chr22 35343242 N chr22 35343721 N DUP 8
SRR1766486.701308 chr22 35343084 N chr22 35343798 N DUP 5
SRR1766478.11889826 chr22 35343099 N chr22 35343813 N DUP 5
SRR1766453.757372 chr22 35343894 N chr22 35344118 N DUP 3
SRR1766472.4162160 chr22 35343485 N chr22 35344059 N DUP 2
SRR1766479.12844044 chr22 35343477 N chr22 35344043 N DEL 1
SRR1766472.787716 chr22 35343508 N chr22 35344084 N DEL 5
SRR1766451.8109115 chr22 35343508 N chr22 35344084 N DEL 5
SRR1766464.9814916 chr22 35342927 N chr22 35344084 N DEL 5
SRR1766454.1108230 chr22 35342930 N chr22 35344087 N DEL 5
SRR1766442.22647289 chr22 35342932 N chr22 35344089 N DEL 5
SRR1766458.704410 chr22 35343528 N chr22 35344100 N DEL 1
SRR1766445.4255998 chr22 35342971 N chr22 35344190 N DEL 5
SRR1766451.6128293 chr2 117643574 N chr2 117643742 N DEL 1
SRR1766461.9241348 chr2 117643574 N chr2 117643742 N DEL 2
SRR1766469.5288738 chr2 117643589 N chr2 117643669 N DEL 13
SRR1766467.4962233 chr2 117643589 N chr2 117643669 N DEL 14
SRR1766484.7938859 chr2 117643589 N chr2 117643669 N DEL 14
SRR1766450.4983810 chr2 117643600 N chr2 117643742 N DEL 15
SRR1766442.41170099 chr2 117643612 N chr2 117643669 N DEL 13
SRR1766479.3488358 chr2 117643563 N chr2 117643630 N DUP 26
SRR1766459.3930887 chr2 117643612 N chr2 117643716 N DEL 22
SRR1766450.4935025 chr2 117643642 N chr2 117643744 N DEL 9
SRR1766478.2952910 chr2 117643563 N chr2 117643630 N DUP 26
SRR1766447.7657057 chr2 117643581 N chr2 117643651 N DUP 14
SRR1766475.321428 chr2 117643581 N chr2 117643651 N DUP 14
SRR1766473.6403983 chr2 117643588 N chr2 117643663 N DUP 18
SRR1766443.6199221 chr2 117643583 N chr2 117643643 N DEL 10
SRR1766481.830855 chr2 117643579 N chr2 117643674 N DEL 6
SRR1766475.11318762 chr2 117643579 N chr2 117643747 N DEL 9
SRR1766442.37490237 chr2 117643666 N chr2 117643743 N DEL 13
SRR1766464.8795132 chr4 186129119 N chr4 186129316 N DEL 5
SRR1766461.5189018 chr7 144859583 N chr7 144859676 N DEL 7
SRR1766446.554344 chr7 144859583 N chr7 144859676 N DEL 7
SRR1766467.1298611 chr11 69398338 N chr11 69398470 N DUP 5
SRR1766481.7647243 chr11 69398353 N chr11 69398487 N DEL 1
SRR1766450.7320547 chr11 69398445 N chr11 69398526 N DEL 5
SRR1766460.6171667 chr11 69398350 N chr11 69398587 N DEL 2
SRR1766442.44296059 chr11 69398455 N chr11 69398599 N DEL 5
SRR1766482.5913511 chr11 69398359 N chr11 69398690 N DEL 5
SRR1766464.4190977 chr14 106309111 N chr14 106309189 N DUP 1
SRR1766474.3331344 chr16 15518017 N chr16 15518086 N DUP 1
SRR1766480.982051 chr16 15518011 N chr16 15518086 N DEL 6
SRR1766442.16062081 chr16 15518124 N chr16 15518173 N DUP 5
SRR1766449.1724361 chr16 15518068 N chr16 15518141 N DEL 5
SRR1766476.6192138 chr16 33385929 N chr16 33386038 N DEL 4
SRR1766463.961025 chr16 33385861 N chr16 33386050 N DUP 4
SRR1766448.11039860 chr7 98242604 N chr7 98242983 N DEL 5
SRR1766474.3247988 chr7 98242707 N chr7 98243192 N DEL 3
SRR1766484.4424215 chr7 98242710 N chr7 98242916 N DEL 5
SRR1766444.1873712 chr7 98242708 N chr7 98242898 N DEL 5
SRR1766442.30077399 chr7 98242722 N chr7 98242936 N DEL 2
SRR1766459.7648564 chr7 98242710 N chr7 98242916 N DEL 10
SRR1766449.1934320 chr7 98242677 N chr7 98243204 N DUP 10
SRR1766450.10299331 chr7 98242740 N chr7 98242950 N DEL 16
SRR1766466.6080538 chr7 98242740 N chr7 98242950 N DEL 10
SRR1766471.2511842 chr7 98242854 N chr7 98243190 N DEL 2
SRR1766459.11334197 chr7 98242582 N chr7 98242752 N DEL 4
SRR1766463.9569264 chr7 98242635 N chr7 98242805 N DEL 3
SRR1766451.8430121 chr7 98242722 N chr7 98242888 N DEL 10
SRR1766475.72241 chr7 98242729 N chr7 98243136 N DUP 23
SRR1766446.3423439 chr7 98242729 N chr7 98243136 N DUP 26
SRR1766451.8963773 chr7 98242720 N chr7 98242882 N DEL 14
SRR1766483.7689659 chr7 98242697 N chr7 98242907 N DEL 4
SRR1766482.10862535 chr7 98242738 N chr7 98242932 N DEL 5
SRR1766483.2533620 chr7 98242585 N chr7 98242932 N DEL 10
SRR1766442.36839067 chr7 98242580 N chr7 98242939 N DEL 5
SRR1766458.7674319 chr7 98242705 N chr7 98243062 N DUP 2
SRR1766469.9836517 chr7 98242705 N chr7 98243062 N DUP 4
SRR1766482.9868772 chr7 98242580 N chr7 98242955 N DEL 4
SRR1766475.3910586 chr7 98242680 N chr7 98243069 N DUP 9
SRR1766452.5261696 chr7 98242901 N chr7 98243073 N DUP 23
SRR1766486.5729006 chr7 98242680 N chr7 98243069 N DUP 17
SRR1766445.3465306 chr7 98242680 N chr7 98243069 N DUP 17
SRR1766459.5195443 chr7 98242680 N chr7 98243069 N DUP 17
SRR1766445.3465306 chr7 98242710 N chr7 98243099 N DUP 16
SRR1766481.2920189 chr7 98242680 N chr7 98243069 N DUP 17
SRR1766472.319119 chr7 98242631 N chr7 98243010 N DEL 10
SRR1766477.3241455 chr7 98242912 N chr7 98243104 N DUP 5
SRR1766465.6082402 chr7 98242623 N chr7 98243002 N DEL 6
SRR1766483.4972764 chr7 98243151 N chr7 98243236 N DEL 13
SRR1766445.2933269 chr7 98242933 N chr7 98243125 N DUP 10
SRR1766473.7601517 chr7 98242912 N chr7 98243134 N DUP 1
SRR1766442.30077399 chr7 98242920 N chr7 98243138 N DUP 7
SRR1766445.10598649 chr7 98243175 N chr7 98243286 N DUP 9
SRR1766460.7656836 chr7 98243143 N chr7 98243197 N DUP 13
SRR1766475.8964712 chr7 98242588 N chr7 98243186 N DEL 11
SRR1766461.4851364 chr7 98242859 N chr7 98243215 N DEL 10
SRR1766479.7612018 chr7 98243185 N chr7 98243242 N DEL 5
SRR1766478.7636865 chr7 98242583 N chr7 98243245 N DEL 15
SRR1766454.1422690 chr7 98243196 N chr7 98243253 N DEL 4
SRR1766472.11992491 chr7 98242762 N chr7 98243255 N DEL 5
SRR1766477.11377730 chr7 98243199 N chr7 98243256 N DEL 1
SRR1766454.6385194 chr7 98242687 N chr7 98243264 N DEL 7
SRR1766476.10898224 chr7 98242578 N chr7 98243264 N DEL 3
SRR1766452.73185 chr7 98242580 N chr7 98243274 N DEL 4
SRR1766448.6005268 chr2 90385464 N chr2 90385649 N DUP 1
SRR1766482.3425912 chr2 90385464 N chr2 90385649 N DUP 1
SRR1766442.36322747 chr2 90385338 N chr2 90385540 N DUP 1
SRR1766451.4623070 chr2 90385338 N chr2 90385540 N DUP 1
SRR1766478.10126501 chr2 90385338 N chr2 90385540 N DUP 1
SRR1766478.884379 chr2 90385411 N chr2 90385505 N DUP 5
SRR1766456.5712240 chr2 90385556 N chr2 90385607 N DUP 2
SRR1766468.6957284 chr2 90385324 N chr2 90385656 N DUP 5
SRR1766470.2970001 chr2 90385341 N chr2 90385569 N DUP 5
SRR1766452.3711307 chr2 90385520 N chr2 90385649 N DUP 5
SRR1766465.6947226 chr2 90385316 N chr2 90385485 N DUP 1
SRR1766451.7449198 chr2 90385324 N chr2 90385656 N DUP 5
SRR1766481.5925425 chr2 90385324 N chr2 90385656 N DUP 5
SRR1766451.6562554 chr7 56374456 N chr7 56374635 N DUP 5
SRR1766477.2086417 chr7 56374482 N chr7 56374579 N DUP 5
SRR1766483.7744340 chr7 56374508 N chr7 56374638 N DUP 5
SRR1766442.47066220 chr7 56374501 N chr7 56374631 N DUP 5
SRR1766442.333445 chr7 56374501 N chr7 56374631 N DUP 5
SRR1766472.8106085 chr7 56374505 N chr7 56374635 N DUP 5
SRR1766484.11544905 chr7 56374505 N chr7 56374635 N DUP 5
SRR1766485.8900953 chr7 56374505 N chr7 56374635 N DUP 5
SRR1766482.12349739 chr7 56374508 N chr7 56374638 N DUP 5
SRR1766465.10512950 chr7 56374508 N chr7 56374638 N DUP 5
SRR1766448.10254267 chr7 56374510 N chr7 56374640 N DUP 5
SRR1766482.10472016 chr7 56374510 N chr7 56374640 N DUP 5
SRR1766459.1327909 chr7 56374511 N chr7 56374641 N DUP 5
SRR1766463.8453321 chr7 56374434 N chr7 56374532 N DEL 1
SRR1766442.5856380 chr7 56374462 N chr7 56374561 N DEL 5
SRR1766463.10821881 chr7 56374462 N chr7 56374561 N DEL 5
SRR1766449.10083364 chr7 56374466 N chr7 56374565 N DEL 5
SRR1766485.10489570 chr7 56374464 N chr7 56374563 N DEL 5
SRR1766484.4849709 chr7 56374466 N chr7 56374565 N DEL 5
SRR1766482.7184330 chr7 56374471 N chr7 56374570 N DEL 5
SRR1766480.6377997 chr7 56374474 N chr7 56374573 N DEL 3
SRR1766453.7105339 chr7 56374476 N chr7 56374575 N DEL 1
SRR1766469.4359348 chr7 56374476 N chr7 56374575 N DEL 1
SRR1766486.2282401 chr7 56374476 N chr7 56374575 N DEL 1
SRR1766480.5170612 chr7 56374442 N chr7 56374589 N DEL 5
SRR1766444.5917304 chr7 56374478 N chr7 56374610 N DEL 1
SRR1766450.2912706 chr7 56374444 N chr7 56374624 N DEL 5
SRR1766478.4704905 chr7 56374502 N chr7 56374634 N DEL 5
SRR1766442.34405836 chr14 105693685 N chr14 105693776 N DUP 13
SRR1766456.1765955 chr14 105693591 N chr14 105693682 N DEL 13
SRR1766483.3675680 chr14 105693504 N chr14 105693690 N DEL 9
SRR1766477.7985835 chr14 105693773 N chr14 105693850 N DUP 30
SRR1766465.4756042 chr14 105693514 N chr14 105693782 N DEL 1
SRR1766469.1574397 chr14 105693724 N chr14 105693849 N DUP 13
SRR1766483.10386505 chr14 105693724 N chr14 105693849 N DUP 13
SRR1766444.6154220 chr14 105693632 N chr14 105693799 N DUP 8
SRR1766455.8863995 chr14 105693695 N chr14 105694434 N DUP 2
SRR1766449.35250 chr14 105693695 N chr14 105694434 N DUP 2
SRR1766442.41494110 chr14 105693815 N chr14 105694234 N DEL 2
SRR1766451.9882016 chr14 105693807 N chr14 105694226 N DEL 5
SRR1766482.6452191 chr14 105693685 N chr14 105693776 N DUP 18
SRR1766467.6138329 chr14 105693767 N chr14 105693898 N DEL 13
SRR1766485.5430354 chr14 105693685 N chr14 105693776 N DUP 23
SRR1766456.1765955 chr14 105693767 N chr14 105693898 N DEL 13
SRR1766480.7451536 chr14 105693767 N chr14 105693898 N DEL 13
SRR1766447.11079155 chr14 105693625 N chr14 105693844 N DUP 1
SRR1766450.5905352 chr14 105693849 N chr14 105694641 N DEL 9
SRR1766470.5418221 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766453.1635179 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766461.3897103 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766482.7587429 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766447.6165974 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766460.2399364 chr14 105693624 N chr14 105693991 N DUP 15
SRR1766466.2330993 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766483.2379837 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766475.4980514 chr14 105693734 N chr14 105693911 N DEL 3
SRR1766479.4308506 chr14 105693991 N chr14 105694226 N DEL 7
SRR1766463.1477430 chr14 105693721 N chr14 105693898 N DEL 13
SRR1766462.3769719 chr14 105694008 N chr14 105694175 N DEL 12
SRR1766474.1253906 chr14 105693764 N chr14 105693993 N DUP 14
SRR1766479.848576 chr14 105693636 N chr14 105693899 N DEL 13
SRR1766485.10482168 chr14 105693586 N chr14 105693913 N DEL 1
SRR1766442.15504051 chr14 105693640 N chr14 105693903 N DEL 10
SRR1766453.2862649 chr14 105694027 N chr14 105694725 N DEL 5
SRR1766474.3952943 chr14 105693488 N chr14 105693904 N DUP 11
SRR1766442.40174251 chr14 105694033 N chr14 105695209 N DEL 8
SRR1766446.2436237 chr14 105694035 N chr14 105694226 N DEL 4
SRR1766480.5161219 chr14 105694035 N chr14 105694226 N DEL 4
SRR1766480.5435223 chr14 105693632 N chr14 105694075 N DUP 5
SRR1766486.2134703 chr14 105694080 N chr14 105694640 N DEL 9
SRR1766467.11257614 chr14 105693971 N chr14 105694254 N DUP 5
SRR1766470.230018 chr14 105693756 N chr14 105694063 N DUP 1
SRR1766479.5959405 chr14 105693680 N chr14 105694075 N DUP 1
SRR1766454.4159986 chr14 105693775 N chr14 105693998 N DEL 5
SRR1766442.2051280 chr14 105694118 N chr14 105694245 N DEL 10
SRR1766460.754203 chr14 105693713 N chr14 105694032 N DEL 5
SRR1766451.416995 chr14 105693713 N chr14 105694032 N DEL 5
SRR1766482.7318132 chr14 105693643 N chr14 105694040 N DEL 5
SRR1766458.8115922 chr14 105693647 N chr14 105694086 N DEL 1
SRR1766463.2498035 chr14 105693660 N chr14 105694229 N DUP 3
SRR1766481.2270202 chr14 105694231 N chr14 105695093 N DEL 5
SRR1766462.9636172 chr14 105694345 N chr14 105694462 N DEL 1
SRR1766456.5459490 chr14 105694201 N chr14 105694410 N DEL 15
SRR1766442.40990022 chr14 105693788 N chr14 105694750 N DUP 15
SRR1766484.4321590 chr14 105694649 N chr14 105694784 N DUP 5
SRR1766446.2603995 chr14 105694158 N chr14 105694860 N DUP 10
SRR1766481.11539659 chr14 105694783 N chr14 105695064 N DUP 4
SRR1766471.7234007 chr14 105694764 N chr14 105695037 N DEL 5
SRR1766443.2468488 chr2 29393136 N chr2 29393186 N DUP 8
SRR1766467.7750244 chr1 153575119 N chr1 153575393 N DEL 5
SRR1766452.9594788 chr1 153575049 N chr1 153575564 N DUP 1
SRR1766453.5631924 chr1 153575044 N chr1 153575601 N DEL 3
SRR1766442.30736685 chr11 38147208 N chr11 38147263 N DUP 10
SRR1766448.4024225 chrX 766364 N chrX 766637 N DUP 5
SRR1766457.9349281 chrX 766444 N chrX 766582 N DEL 5
SRR1766469.6909650 chr11 3359329 N chr11 3359498 N DEL 5
SRR1766442.46591202 chr11 3359330 N chr11 3359497 N DUP 1
SRR1766471.7602032 chr11 3359330 N chr11 3359497 N DUP 5
SRR1766482.10034420 chr1 2976660 N chr1 2976884 N DEL 7
SRR1766454.10962373 chr1 2976705 N chr1 2977962 N DUP 5
SRR1766469.6243408 chr1 2976990 N chr1 2977255 N DEL 5
SRR1766476.11179653 chr1 2976843 N chr1 2977372 N DUP 2
SRR1766452.9897100 chr1 2977693 N chr1 2977772 N DUP 34
SRR1766478.4781638 chr1 2977476 N chr1 2978018 N DUP 7
SRR1766475.11251595 chr1 2977608 N chr1 2977913 N DEL 3
SRR1766442.37323400 chr1 2976954 N chr1 2978074 N DEL 1
SRR1766458.8687225 chr1 2977522 N chr1 2978110 N DEL 11
SRR1766464.7820864 chr14 100546482 N chr14 100546602 N DEL 3
SRR1766457.3759168 chr14 100546569 N chr14 100546620 N DEL 7
SRR1766475.1560710 chr14 100546488 N chr14 100546608 N DEL 15
SRR1766449.8325027 chr9 134636930 N chr9 134636989 N DUP 2
SRR1766476.7426164 chr9 134636930 N chr9 134637009 N DUP 5
SRR1766485.2021711 chr9 134636945 N chr9 134637044 N DUP 6
SRR1766445.1904144 chr7 62441954 N chr7 62442120 N DEL 3
SRR1766451.2227258 chr7 62441866 N chr7 62441960 N DEL 5
SRR1766452.8384836 chr7 62441866 N chr7 62441960 N DEL 5
SRR1766482.1701519 chr7 62441868 N chr7 62441962 N DEL 5
SRR1766449.1033935 chr7 62442006 N chr7 62442124 N DUP 1
SRR1766443.10178981 chr7 62442169 N chr7 62442624 N DEL 5
SRR1766446.2238516 chr7 62442169 N chr7 62442624 N DEL 5
SRR1766475.5293393 chr7 62442169 N chr7 62442624 N DEL 5
SRR1766469.2136012 chr7 62442193 N chr7 62442646 N DUP 4
SRR1766456.1017640 chr7 62442193 N chr7 62442646 N DUP 4
SRR1766447.1810928 chr7 62442193 N chr7 62442261 N DUP 2
SRR1766455.4722542 chr7 62442193 N chr7 62442261 N DUP 1
SRR1766453.128358 chr7 62441836 N chr7 62442285 N DEL 15
SRR1766472.8443588 chr7 62441885 N chr7 62442413 N DUP 5
SRR1766464.5343314 chr7 62441903 N chr7 62442454 N DUP 3
SRR1766452.8384836 chr7 62441903 N chr7 62442454 N DUP 3
SRR1766476.8389588 chr7 62441903 N chr7 62442454 N DUP 4
SRR1766486.1120897 chr7 62441903 N chr7 62442454 N DUP 7
SRR1766447.3670339 chr7 62442456 N chr7 62442751 N DEL 15
SRR1766450.1049268 chr7 62442454 N chr7 62442698 N DUP 21
SRR1766442.39480516 chr7 62442460 N chr7 62442580 N DUP 7
SRR1766451.1203630 chr7 62441910 N chr7 62442463 N DEL 1
SRR1766470.1050489 chr7 62441909 N chr7 62442462 N DEL 2
SRR1766455.4473224 chr7 62442468 N chr7 62442637 N DUP 5
SRR1766465.11230860 chr7 62441916 N chr7 62442590 N DEL 10
SRR1766469.5913933 chr7 62441870 N chr7 62442583 N DEL 8
SRR1766478.191833 chr7 62441916 N chr7 62442590 N DEL 10
SRR1766478.362698 chr7 62441874 N chr7 62442587 N DEL 3
SRR1766484.206190 chr7 62441874 N chr7 62442587 N DEL 3
SRR1766460.5835705 chr7 62441856 N chr7 62442714 N DUP 5
SRR1766442.28974248 chr7 62441834 N chr7 62442596 N DEL 1
SRR1766442.46964375 chr7 62442623 N chr7 62442720 N DUP 4
SRR1766485.4736569 chr7 62441961 N chr7 62442630 N DEL 8
SRR1766471.2210920 chr7 62442660 N chr7 62442734 N DUP 25
SRR1766466.3515121 chr2 206372205 N chr2 206372276 N DEL 2
SRR1766481.7166101 chr2 206372205 N chr2 206372276 N DEL 3
SRR1766485.4397259 chr2 206372215 N chr2 206372414 N DEL 5
SRR1766442.4616750 chr2 206372285 N chr2 206372350 N DEL 2
SRR1766463.3542640 chr2 206372285 N chr2 206372350 N DEL 2
SRR1766442.41340391 chr2 206372285 N chr2 206372350 N DEL 5
SRR1766481.5444875 chr2 206372285 N chr2 206372350 N DEL 5
SRR1766442.698419 chr2 206372218 N chr2 206372321 N DEL 12
SRR1766451.6006236 chr2 206372162 N chr2 206372327 N DEL 6
SRR1766453.5812362 chr2 206372218 N chr2 206372321 N DEL 12
SRR1766454.9060274 chr2 206372220 N chr2 206372323 N DEL 10
SRR1766453.5600855 chr2 206372218 N chr2 206372321 N DEL 12
SRR1766454.10025593 chr2 206372344 N chr2 206372407 N DUP 5
SRR1766442.23888005 chr2 206372344 N chr2 206372407 N DUP 5
SRR1766460.1216866 chr2 206372344 N chr2 206372407 N DUP 5
SRR1766445.727337 chr2 206372347 N chr2 206372410 N DUP 5
SRR1766469.5953152 chr2 206372348 N chr2 206372411 N DUP 5
SRR1766466.9554349 chr2 206372352 N chr2 206372415 N DUP 5
SRR1766473.11191124 chr2 206372354 N chr2 206372417 N DUP 5
SRR1766478.5996974 chr2 206372354 N chr2 206372417 N DUP 5
SRR1766486.5142640 chr2 206372358 N chr2 206372421 N DUP 1
SRR1766449.479769 chr4 70516455 N chr4 70516554 N DEL 4
SRR1766453.10872049 chr4 70516452 N chr4 70516561 N DEL 8
SRR1766479.2594768 chr4 70516460 N chr4 70516561 N DEL 10
SRR1766462.776988 chr4 70516460 N chr4 70516561 N DEL 12
SRR1766473.10455670 chr4 70516460 N chr4 70516561 N DEL 13
SRR1766466.5291348 chr4 70516459 N chr4 70516538 N DEL 18
SRR1766456.2374242 chr4 70516461 N chr4 70516562 N DEL 7
SRR1766462.2101035 chr4 70516462 N chr4 70516563 N DEL 6
SRR1766464.1177064 chr4 70516455 N chr4 70516556 N DEL 13
SRR1766473.8503848 chr4 70516459 N chr4 70516560 N DEL 9
SRR1766485.7186165 chr4 70516455 N chr4 70516556 N DEL 13
SRR1766460.8528614 chr4 70516458 N chr4 70516563 N DEL 7
SRR1766473.808173 chr4 70516455 N chr4 70516564 N DEL 10
SRR1766486.4249754 chr4 70516465 N chr4 70516585 N DEL 6
SRR1766447.3559350 chr4 70516475 N chr4 70516587 N DEL 6
SRR1766470.6985422 chr22 38807029 N chr22 38807303 N DEL 1
SRR1766453.3771907 chr22 38806854 N chr22 38807322 N DUP 5
SRR1766443.8920110 chr2 64375734 N chr2 64375823 N DEL 2
SRR1766467.9128986 chr2 64375753 N chr2 64376213 N DEL 24
SRR1766443.179353 chr2 64375753 N chr2 64376213 N DEL 29
SRR1766442.8935067 chr2 64375803 N chr2 64375868 N DEL 13
SRR1766442.45717887 chr2 64375788 N chr2 64375868 N DEL 5
SRR1766464.4429184 chr2 64375746 N chr2 64376215 N DEL 8
SRR1766470.4626732 chr2 64375858 N chr2 64376377 N DEL 13
SRR1766456.6162646 chr2 64375868 N chr2 64375952 N DUP 19
SRR1766461.8014131 chr2 64375795 N chr2 64376208 N DEL 24
SRR1766479.1785907 chr2 64375822 N chr2 64375950 N DUP 11
SRR1766468.7482571 chr2 64375735 N chr2 64375872 N DUP 9
SRR1766445.7757027 chr2 64375878 N chr2 64376298 N DUP 8
SRR1766456.2984199 chr2 64375822 N chr2 64375883 N DUP 9
SRR1766478.3040180 chr2 64375800 N chr2 64376035 N DEL 19
SRR1766482.4175847 chr2 64375740 N chr2 64375815 N DUP 10
SRR1766448.2893483 chr2 64375739 N chr2 64375917 N DUP 7
SRR1766452.5794147 chr2 64375786 N chr2 64375917 N DUP 4
SRR1766443.8429926 chr2 64375748 N chr2 64375917 N DUP 17
SRR1766479.12516280 chr2 64375838 N chr2 64376193 N DEL 13
SRR1766476.2181495 chr2 64375766 N chr2 64376092 N DEL 18
SRR1766456.1368625 chr2 64375800 N chr2 64375880 N DEL 13
SRR1766484.11814463 chr2 64375788 N chr2 64375868 N DEL 5
SRR1766447.7497881 chr2 64375897 N chr2 64376202 N DEL 11
SRR1766482.7255812 chr2 64375803 N chr2 64375960 N DUP 5
SRR1766482.10989921 chr2 64375749 N chr2 64375876 N DEL 10
SRR1766469.1311668 chr2 64376173 N chr2 64376289 N DUP 13
SRR1766455.658195 chr2 64375751 N chr2 64375881 N DEL 7
SRR1766471.10368059 chr2 64375770 N chr2 64375905 N DEL 2
SRR1766466.2982883 chr2 64375915 N chr2 64376221 N DUP 10
SRR1766450.6851033 chr2 64375735 N chr2 64375974 N DUP 5
SRR1766442.29805931 chr2 64375901 N chr2 64376283 N DUP 6
SRR1766476.2181495 chr2 64375859 N chr2 64375980 N DEL 5
SRR1766457.5161250 chr2 64375782 N chr2 64375906 N DEL 1
SRR1766446.5868090 chr2 64375763 N chr2 64375999 N DUP 9
SRR1766459.3574931 chr2 64375794 N chr2 64375921 N DEL 8
SRR1766467.11058203 chr2 64375918 N chr2 64376069 N DUP 11
SRR1766463.318073 chr2 64375874 N chr2 64376338 N DUP 13
SRR1766446.8520773 chr2 64375900 N chr2 64375975 N DUP 10
SRR1766454.435312 chr2 64375807 N chr2 64376005 N DUP 9
SRR1766447.4097105 chr2 64375735 N chr2 64375977 N DUP 18
SRR1766473.8323290 chr2 64375797 N chr2 64376187 N DEL 11
SRR1766483.6953215 chr2 64375747 N chr2 64375989 N DUP 11
SRR1766445.8500216 chr2 64375828 N chr2 64376345 N DUP 13
SRR1766476.9592672 chr2 64375874 N chr2 64375952 N DUP 13
SRR1766465.992677 chr2 64375874 N chr2 64375990 N DUP 16
SRR1766472.10661683 chr2 64375750 N chr2 64375912 N DEL 3
SRR1766454.770780 chr2 64375874 N chr2 64376338 N DUP 9
SRR1766469.8584880 chr2 64375874 N chr2 64376338 N DUP 13
SRR1766478.10710367 chr2 64375944 N chr2 64376173 N DEL 13
SRR1766456.5515521 chr2 64375958 N chr2 64376187 N DEL 3
SRR1766456.5515521 chr2 64375874 N chr2 64376069 N DUP 10
SRR1766473.8323290 chr2 64375838 N chr2 64375956 N DEL 8
SRR1766455.2164592 chr2 64375735 N chr2 64376059 N DUP 4
SRR1766480.2497720 chr2 64375813 N chr2 64376039 N DEL 24
SRR1766479.5991748 chr2 64375958 N chr2 64376187 N DEL 9
SRR1766453.3260526 chr2 64375824 N chr2 64376016 N DUP 11
SRR1766477.3223782 chr2 64375736 N chr2 64376086 N DUP 16
SRR1766480.3121727 chr2 64375825 N chr2 64376017 N DUP 10
SRR1766452.4615466 chr2 64375874 N chr2 64375990 N DUP 10
SRR1766476.6838937 chr2 64375874 N chr2 64376256 N DUP 14
SRR1766442.7354464 chr2 64375874 N chr2 64375987 N DUP 13
SRR1766478.9075524 chr2 64375886 N chr2 64376347 N DUP 10
SRR1766456.3795525 chr2 64375874 N chr2 64375990 N DUP 10
SRR1766443.2878377 chr2 64376020 N chr2 64376208 N DEL 7
SRR1766453.3864471 chr2 64375874 N chr2 64375990 N DUP 10
SRR1766480.4931241 chr2 64375874 N chr2 64375987 N DUP 13
SRR1766478.2533618 chr2 64375824 N chr2 64376098 N DUP 3
SRR1766443.853062 chr2 64375944 N chr2 64376173 N DEL 6
SRR1766446.5563350 chr2 64375868 N chr2 64375952 N DUP 11
SRR1766455.1791120 chr2 64375794 N chr2 64375921 N DEL 8
SRR1766452.8880707 chr2 64375780 N chr2 64376208 N DEL 16
SRR1766478.9243993 chr2 64375794 N chr2 64375880 N DEL 5
SRR1766460.1816860 chr2 64375739 N chr2 64376139 N DUP 8
SRR1766476.11115489 chr2 64375735 N chr2 64376147 N DUP 9
SRR1766450.8013720 chr2 64376058 N chr2 64376139 N DUP 7
SRR1766481.3941539 chr2 64375737 N chr2 64376093 N DUP 13
SRR1766453.3880162 chr2 64375795 N chr2 64376145 N DUP 12
SRR1766447.10281777 chr2 64375874 N chr2 64375987 N DUP 8
SRR1766455.3219840 chr2 64375944 N chr2 64376135 N DEL 11
SRR1766442.31007132 chr2 64375736 N chr2 64376212 N DUP 4
SRR1766455.3924306 chr2 64375967 N chr2 64376219 N DEL 29
SRR1766446.5082191 chr2 64375874 N chr2 64376215 N DUP 8
SRR1766472.3668981 chr2 64375782 N chr2 64375874 N DEL 11
SRR1766469.11046682 chr2 64375747 N chr2 64375989 N DUP 18
SRR1766484.10342390 chr2 64375936 N chr2 64376203 N DEL 7
SRR1766458.1451090 chr2 64375737 N chr2 64375856 N DUP 13
SRR1766481.9487105 chr2 64375791 N chr2 64375874 N DEL 13
SRR1766456.5934369 chr2 64375737 N chr2 64375979 N DUP 18
SRR1766479.3600612 chr2 64375884 N chr2 64376218 N DEL 15
SRR1766456.3609411 chr2 64375750 N chr2 64376187 N DEL 6
SRR1766473.3927163 chr2 64375747 N chr2 64376071 N DUP 6
SRR1766443.4327616 chr2 64375880 N chr2 64376221 N DUP 8
SRR1766474.7707327 chr2 64375918 N chr2 64376259 N DUP 8
SRR1766455.8841869 chr2 64376174 N chr2 64376290 N DUP 10
SRR1766464.4429184 chr2 64375900 N chr2 64375972 N DUP 8
SRR1766478.9075524 chr2 64375947 N chr2 64376018 N DEL 22
SRR1766457.4284435 chr2 64375737 N chr2 64375979 N DUP 15
SRR1766448.10928298 chr2 64375812 N chr2 64375975 N DUP 13
SRR1766469.6997753 chr2 64375737 N chr2 64375979 N DUP 17
SRR1766452.8798532 chr2 64375801 N chr2 64376344 N DUP 13
SRR1766457.8770427 chr2 64375982 N chr2 64376173 N DEL 8
SRR1766472.5977698 chr2 64375807 N chr2 64376116 N DUP 11
SRR1766483.11075530 chr2 64375795 N chr2 64376069 N DUP 13
SRR1766485.7896807 chr2 64375944 N chr2 64376018 N DEL 16
SRR1766442.31898883 chr2 64375838 N chr2 64376231 N DEL 16
SRR1766445.9821722 chr2 64376005 N chr2 64376193 N DEL 10
SRR1766447.8266882 chr2 64375758 N chr2 64376310 N DUP 12
SRR1766468.5671200 chr2 64375786 N chr2 64376214 N DEL 9
SRR1766445.9506881 chr2 64375751 N chr2 64376214 N DEL 8
SRR1766446.6181696 chr2 64375882 N chr2 64376216 N DEL 7
SRR1766482.2343075 chr2 64375791 N chr2 64376219 N DEL 4
SRR1766484.31648 chr2 64375944 N chr2 64376018 N DEL 12
SRR1766447.8266882 chr2 64375759 N chr2 64376308 N DUP 14
SRR1766484.10428003 chr2 64375746 N chr2 64376295 N DUP 11
SRR1766454.3658398 chr2 64375822 N chr2 64376333 N DUP 9
SRR1766481.2994782 chr2 64375739 N chr2 64376323 N DUP 8
SRR1766450.8013720 chr2 64375862 N chr2 64376173 N DEL 10
SRR1766448.3886690 chr2 64375874 N chr2 64376297 N DUP 17
SRR1766478.4083906 chr2 64375735 N chr2 64376346 N DUP 7
SRR1766442.43832294 chr2 64375761 N chr2 64376247 N DEL 8
SRR1766479.4471343 chr2 64375874 N chr2 64376145 N DUP 18
SRR1766463.1685291 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766478.6116256 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766481.409521 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766463.2518470 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766445.4818764 chr2 64375798 N chr2 64376308 N DEL 10
SRR1766460.8782180 chr2 64375757 N chr2 64376308 N DEL 7
SRR1766442.20259212 chr2 64375758 N chr2 64376309 N DEL 5
SRR1766461.1758616 chr2 64375754 N chr2 64376311 N DEL 5
SRR1766474.6821041 chr2 64375754 N chr2 64376352 N DEL 5
SRR1766449.5423178 chr2 94283690 N chr2 94283788 N DEL 10
SRR1766479.4667760 chrX 1735658 N chrX 1735815 N DEL 2
SRR1766471.8460006 chrX 35692462 N chrX 35692559 N DUP 31
SRR1766483.6209409 chrX 35692537 N chrX 35692610 N DUP 31
SRR1766477.7315024 chrX 35692492 N chrX 35692559 N DUP 28
SRR1766447.3730770 chrX 35692492 N chrX 35692559 N DUP 41
SRR1766461.9713008 chrX 35692492 N chrX 35692559 N DUP 41
SRR1766475.7968703 chrX 35692492 N chrX 35692559 N DUP 34
SRR1766455.386080 chrX 35692492 N chrX 35692559 N DUP 31
SRR1766460.3099710 chrX 35692492 N chrX 35692559 N DUP 40
SRR1766477.943855 chrX 35692503 N chrX 35692560 N DUP 20
SRR1766462.10448532 chrX 35692503 N chrX 35692560 N DUP 19
SRR1766479.9065739 chrX 35692503 N chrX 35692560 N DUP 16
SRR1766482.12448661 chrX 35692503 N chrX 35692610 N DUP 19
SRR1766442.25600171 chrX 35692503 N chrX 35692610 N DUP 19
SRR1766472.6339022 chr4 123498553 N chr4 123498747 N DEL 9
SRR1766471.11969579 chr4 123498716 N chr4 123498874 N DUP 6
SRR1766469.481458 chr8 2448044 N chr8 2448116 N DEL 5
SRR1766454.6312347 chr8 2447983 N chr8 2448055 N DUP 5
SRR1766480.809303 chr8 2447983 N chr8 2448055 N DUP 5
SRR1766484.1451048 chr8 2447999 N chr8 2448073 N DEL 4
SRR1766442.1184542 chrX 1472802 N chrX 1472960 N DUP 12
SRR1766481.4523254 chrX 1472956 N chrX 1473199 N DEL 2
SRR1766451.9472057 chrX 1473000 N chrX 1473199 N DEL 13
SRR1766482.6957216 chrX 1472867 N chrX 1473034 N DUP 11
SRR1766448.9250568 chrX 1472917 N chrX 1473202 N DUP 4
SRR1766484.1660444 chrX 1472959 N chrX 1473161 N DUP 8
SRR1766445.4822830 chrX 1473013 N chrX 1473139 N DUP 15
SRR1766477.5946920 chr20 18539123 N chr20 18539424 N DEL 6
SRR1766462.6271552 chr20 18539123 N chr20 18539424 N DEL 7
SRR1766474.8742642 chr20 18539213 N chr20 18539673 N DUP 1
SRR1766442.42441363 chr20 18539319 N chr20 18539618 N DEL 5
SRR1766454.5293583 chr20 18539212 N chr20 18539674 N DEL 1
SRR1766476.5571681 chr5 138143756 N chr5 138143823 N DEL 58
SRR1766484.9328623 chr1 8301322 N chr1 8301463 N DEL 5
SRR1766468.1854140 chr1 8301316 N chr1 8301597 N DEL 34
SRR1766467.10459469 chr1 8301352 N chr1 8301437 N DEL 5
SRR1766466.7843751 chr1 8301356 N chr1 8301441 N DEL 1
SRR1766469.1386354 chr1 8301400 N chr1 8301485 N DEL 5
SRR1766454.8447095 chr1 8301356 N chr1 8301441 N DEL 10
SRR1766455.96219 chr1 8301390 N chr1 8301811 N DEL 5
SRR1766442.40547766 chr1 8301411 N chr1 8301468 N DEL 5
SRR1766446.3687314 chr1 8301356 N chr1 8301441 N DEL 1
SRR1766452.5510176 chr1 8301356 N chr1 8301441 N DEL 12
SRR1766486.8460964 chr1 8301356 N chr1 8301441 N DEL 5
SRR1766461.8633633 chr1 8301484 N chr1 8302044 N DEL 5
SRR1766450.6225578 chr1 8301482 N chr1 8301931 N DEL 11
SRR1766474.4394840 chr1 8301462 N chr1 8301659 N DEL 10
SRR1766446.1088376 chr1 8301456 N chr1 8301653 N DEL 8
SRR1766447.1099627 chr1 8301430 N chr1 8301851 N DEL 10
SRR1766457.5066481 chr1 8301505 N chr1 8301926 N DEL 11
SRR1766467.3794240 chr1 8301437 N chr1 8301548 N DUP 13
SRR1766480.2029925 chr1 8301505 N chr1 8301588 N DUP 10
SRR1766461.2630096 chr1 8301501 N chr1 8301584 N DUP 5
SRR1766471.2724162 chr1 8301428 N chr1 8301567 N DUP 10
SRR1766457.5628980 chr1 8301501 N chr1 8301584 N DUP 5
SRR1766454.847125 chr1 8301542 N chr1 8301961 N DUP 10
SRR1766454.8816610 chr1 8301393 N chr1 8301534 N DEL 4
SRR1766466.9790793 chr1 8301634 N chr1 8301915 N DEL 10
SRR1766478.7043699 chr1 8301658 N chr1 8301939 N DEL 5
SRR1766447.6477887 chr1 8301394 N chr1 8301563 N DEL 1
SRR1766478.2071916 chr1 8301680 N chr1 8302072 N DEL 1
SRR1766468.1854140 chr1 8301301 N chr1 8301582 N DEL 21
SRR1766477.9827703 chr1 8301653 N chr1 8301960 N DUP 10
SRR1766480.6327103 chr1 8301521 N chr1 8301634 N DEL 20
SRR1766473.11015767 chr1 8301497 N chr1 8301666 N DEL 2
SRR1766473.8438433 chr1 8301389 N chr1 8301670 N DEL 5
SRR1766479.13807250 chr1 8301596 N chr1 8301709 N DEL 5
SRR1766482.8668446 chr1 8301457 N chr1 8301710 N DEL 5
SRR1766453.9216938 chr1 8301460 N chr1 8301713 N DEL 5
SRR1766463.7328244 chr1 8301821 N chr1 8302073 N DEL 1
SRR1766450.6225578 chr1 8301379 N chr1 8301716 N DEL 5
SRR1766475.4855356 chr1 8301565 N chr1 8301734 N DEL 5
SRR1766468.2872500 chr1 8301341 N chr1 8301734 N DEL 5
SRR1766485.4436147 chr1 8301393 N chr1 8301758 N DEL 10
SRR1766445.7914758 chr1 8301785 N chr1 8301952 N DUP 30
SRR1766469.631126 chr1 8301380 N chr1 8301745 N DEL 4
SRR1766485.4460136 chr1 8301589 N chr1 8301758 N DEL 12
SRR1766442.4413872 chr1 8301781 N chr1 8301948 N DUP 15
SRR1766463.6086776 chr1 8301586 N chr1 8301783 N DEL 12
SRR1766486.8460964 chr1 8301502 N chr1 8301783 N DEL 10
SRR1766474.2525743 chr1 8301794 N chr1 8301905 N DUP 1
SRR1766444.5759840 chr1 8301690 N chr1 8301831 N DEL 5
SRR1766455.7760761 chr1 8301487 N chr1 8301852 N DEL 5
SRR1766477.4719669 chr1 8301483 N chr1 8301848 N DEL 25
SRR1766442.40547766 chr1 8301486 N chr1 8301851 N DEL 16
SRR1766454.5673377 chr1 8301486 N chr1 8301851 N DEL 16
SRR1766472.6181988 chr1 8301851 N chr1 8301934 N DUP 30
SRR1766461.8633633 chr1 8301486 N chr1 8301851 N DEL 20
SRR1766475.8036736 chr1 8301709 N chr1 8301878 N DEL 11
SRR1766474.8666197 chr1 8301541 N chr1 8301878 N DEL 10
SRR1766442.6311373 chr1 8301709 N chr1 8301878 N DEL 9
SRR1766481.13004859 chr1 8301880 N chr1 8301963 N DUP 5
SRR1766442.1420060 chr1 8301887 N chr1 8301970 N DUP 5
SRR1766472.4891251 chr1 8301906 N chr1 8301961 N DUP 5
SRR1766459.1078409 chr1 8301494 N chr1 8301915 N DEL 5
SRR1766467.5122452 chr1 8301389 N chr1 8302033 N DEL 10
SRR1766450.9037220 chr2 121777114 N chr2 121777207 N DEL 5
SRR1766460.424437 chr2 121777117 N chr2 121777168 N DUP 5
SRR1766459.1363886 chr2 121777156 N chr2 121777221 N DUP 8
SRR1766484.1797632 chr2 121777159 N chr2 121777244 N DUP 1
SRR1766473.4348518 chr11 71124166 N chr11 71124339 N DUP 1
SRR1766458.2207851 chr8 132187850 N chr8 132187959 N DEL 2
SRR1766456.4528995 chr8 132187841 N chr8 132187944 N DEL 5
SRR1766452.8361062 chr8 132187854 N chr8 132187957 N DEL 5
SRR1766475.4503166 chr8 132187863 N chr8 132188005 N DEL 7
SRR1766460.2163640 chr8 132187901 N chr8 132187983 N DEL 25
SRR1766458.3312228 chr8 132187932 N chr8 132188029 N DEL 10
SRR1766451.5424159 chr8 132187947 N chr8 132188000 N DUP 10
SRR1766442.15546467 chr8 132188012 N chr8 132188083 N DUP 5
SRR1766485.4977296 chr8 132187791 N chr8 132188011 N DEL 14
SRR1766464.9104850 chr8 132187788 N chr8 132188017 N DEL 3
SRR1766459.1325541 chr8 132187782 N chr8 132188065 N DEL 5
SRR1766484.7598318 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766476.5880276 chr5 180615360 N chr5 180615464 N DEL 15
SRR1766456.6470003 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766452.7138667 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766484.7138450 chr5 180615503 N chr5 180615562 N DEL 22
SRR1766472.2125366 chr5 180615386 N chr5 180615548 N DEL 10
SRR1766447.2809373 chr5 180615335 N chr5 180615437 N DUP 13
SRR1766442.9426009 chr5 180615317 N chr5 180615522 N DUP 15
SRR1766448.1807269 chr5 180615318 N chr5 180615420 N DUP 10
SRR1766442.3611502 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766454.4593470 chr5 180615347 N chr5 180615451 N DEL 15
SRR1766474.3271898 chr5 180615347 N chr5 180615451 N DEL 5
SRR1766442.24573789 chr5 180615448 N chr5 180615653 N DUP 4
SRR1766465.9482057 chr5 180615347 N chr5 180615451 N DEL 5
SRR1766486.11910309 chr5 180615347 N chr5 180615451 N DEL 5
SRR1766472.7458730 chr5 180615347 N chr5 180615451 N DEL 5
SRR1766462.7972114 chr5 180615347 N chr5 180615451 N DEL 5
SRR1766453.480081 chr5 180615352 N chr5 180615456 N DEL 5
SRR1766486.9579523 chr5 180615309 N chr5 180615458 N DEL 5
SRR1766455.198855 chr5 180615465 N chr5 180615624 N DUP 30
SRR1766465.5023132 chr5 180615372 N chr5 180615521 N DEL 10
SRR1766451.6290074 chr5 180615445 N chr5 180615591 N DUP 6
SRR1766444.6610758 chr5 180615317 N chr5 180615522 N DUP 20
SRR1766480.2452568 chr5 180615445 N chr5 180615591 N DUP 9
SRR1766481.6316063 chr5 180615420 N chr5 180615611 N DUP 24
SRR1766449.4575616 chr8 22371578 N chr8 22371906 N DEL 6
SRR1766486.3306821 chr8 22371772 N chr8 22372085 N DEL 5
SRR1766463.900643 chr8 22371772 N chr8 22372085 N DEL 5
SRR1766483.4288774 chr8 22371772 N chr8 22372085 N DEL 5
SRR1766467.8090688 chr8 22371773 N chr8 22372086 N DEL 5
SRR1766474.2229789 chr8 22371776 N chr8 22372089 N DEL 5
SRR1766481.10151039 chr8 22371796 N chr8 22372109 N DEL 1
SRR1766442.37695204 chr3 137956899 N chr3 137956974 N DEL 4
SRR1766454.7761521 chr3 137956901 N chr3 137956989 N DUP 2
SRR1766486.5231049 chr3 137956915 N chr3 137957004 N DEL 2
SRR1766473.4435826 chr22 18370593 N chr22 18370646 N DUP 2
SRR1766465.6219816 chr22 18370651 N chr22 18370706 N DEL 25
SRR1766485.11657075 chr22 18370651 N chr22 18370706 N DEL 15
SRR1766480.6806500 chr22 18370628 N chr22 18370710 N DEL 10
SRR1766468.1820484 chr22 18370633 N chr22 18370715 N DEL 6
SRR1766456.5493097 chr22 18370638 N chr22 18370720 N DEL 1
SRR1766453.1413062 chr10 27783269 N chr10 27783634 N DEL 4
SRR1766465.2967605 chr10 27783324 N chr10 27783596 N DEL 2
SRR1766471.11446939 chr10 27783331 N chr10 27783791 N DEL 5
SRR1766483.2500958 chr10 27783459 N chr10 27783640 N DUP 5
SRR1766451.203247 chr10 27783207 N chr10 27783483 N DEL 5
SRR1766455.4469518 chr10 27783414 N chr10 27783593 N DEL 5
SRR1766442.3815949 chr10 27783617 N chr10 27783710 N DUP 3
SRR1766442.46039148 chr10 27783277 N chr10 27783611 N DEL 5
SRR1766459.10523175 chr10 27783627 N chr10 27783844 N DUP 1
SRR1766451.233145 chr10 27783604 N chr10 27783667 N DEL 5
SRR1766453.1544534 chr10 27783635 N chr10 27783762 N DEL 5
SRR1766460.6462817 chr10 27783434 N chr10 27783774 N DEL 3
SRR1766443.636141 chr10 27783513 N chr10 27783791 N DEL 6
SRR1766476.6313398 chr11 3174069 N chr11 3174191 N DEL 5
SRR1766469.9155466 chr2 225783072 N chr2 225783687 N DUP 12
SRR1766442.34340362 chr2 225783082 N chr2 225783681 N DUP 2
SRR1766460.7446245 chr2 225782846 N chr2 225783338 N DEL 5
SRR1766477.7574171 chr2 225783280 N chr2 225783342 N DEL 5
SRR1766442.43672654 chr2 225783087 N chr2 225783376 N DEL 5
SRR1766447.7976738 chr2 225783087 N chr2 225783376 N DEL 5
SRR1766485.11927016 chr2 225783191 N chr2 225783521 N DEL 9
SRR1766475.4779788 chr12 48664595 N chr12 48664900 N DEL 16
SRR1766469.7178186 chr12 48664442 N chr12 48664609 N DEL 2
SRR1766447.9952138 chr12 48664915 N chr12 48665054 N DUP 8
SRR1766458.6594155 chr12 48664740 N chr12 48665041 N DEL 3
SRR1766483.1458972 chr12 48664443 N chr12 48665032 N DEL 12
SRR1766454.9797345 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766458.4243773 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766474.3321557 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766486.11116663 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766484.6698605 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766477.2534543 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766482.7155531 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766468.6151140 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766453.7676675 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766458.1319368 chr21 40821220 N chr21 40821287 N DEL 9
SRR1766445.6153449 chr21 40821194 N chr21 40821287 N DEL 9
SRR1766467.7651482 chr21 40821194 N chr21 40821287 N DEL 9
SRR1766464.9185942 chr21 40821195 N chr21 40821288 N DEL 9
SRR1766480.2981406 chr21 40821196 N chr21 40821289 N DEL 9
SRR1766448.9726418 chr21 40821200 N chr21 40821293 N DEL 9
SRR1766446.7561168 chr21 40821201 N chr21 40821294 N DEL 8
SRR1766447.10229442 chr13 108013563 N chr13 108013653 N DUP 5
SRR1766467.1798646 chr10 68946105 N chr10 68946264 N DUP 5
SRR1766459.4694282 chr10 68946105 N chr10 68946264 N DUP 5
SRR1766442.33222737 chr10 2871852 N chr10 2871910 N DEL 2
SRR1766459.2254822 chr10 2871852 N chr10 2871910 N DEL 3
SRR1766477.3247718 chr10 2871852 N chr10 2871910 N DEL 3
SRR1766478.11701309 chr10 2871852 N chr10 2871910 N DEL 37
SRR1766442.17362191 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766450.2437205 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766451.10089738 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766461.4433608 chr10 2871852 N chr10 2871910 N DEL 49
SRR1766485.9023809 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766456.4442558 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766461.388165 chr10 2871852 N chr10 2871910 N DEL 39
SRR1766453.9816872 chr10 2871859 N chr10 2871942 N DUP 5
SRR1766463.5413813 chr10 2871859 N chr10 2871942 N DUP 7
SRR1766464.2928886 chr10 2871859 N chr10 2871942 N DUP 6
SRR1766474.8808373 chr10 2871859 N chr10 2871942 N DUP 6
SRR1766482.3788811 chr10 2871865 N chr10 2871948 N DUP 3
SRR1766443.6051216 chr10 2871932 N chr10 2872047 N DEL 5
SRR1766460.7725590 chr10 2871986 N chr10 2872099 N DUP 8
SRR1766477.7256797 chr10 2872086 N chr10 2872144 N DEL 5
SRR1766463.5413813 chr10 2871944 N chr10 2872200 N DEL 5
SRR1766462.7897352 chr2 10291518 N chr2 10291583 N DUP 4
SRR1766449.9144307 chr2 10291518 N chr2 10291583 N DUP 8
SRR1766467.7479950 chr2 10291518 N chr2 10291583 N DUP 9
SRR1766456.639110 chr14 74245027 N chr14 74245164 N DEL 8
SRR1766475.3441543 chr6 22792114 N chr6 22792186 N DEL 4
SRR1766477.6967252 chr6 22792114 N chr6 22792186 N DEL 4
SRR1766456.4051609 chr6 22792205 N chr6 22792291 N DEL 8
SRR1766481.3188801 chr10 49105042 N chr10 49105155 N DUP 9
SRR1766453.6126579 chr10 49105155 N chr10 49105275 N DEL 8
SRR1766447.3884509 chr10 49104954 N chr10 49105159 N DUP 4
SRR1766481.6056795 chr10 49104954 N chr10 49105159 N DUP 5
SRR1766467.622409 chr10 49104954 N chr10 49105159 N DUP 7
SRR1766476.1026075 chr10 49105183 N chr10 49105333 N DEL 12
SRR1766471.10114334 chr10 49105226 N chr10 49105361 N DEL 7
SRR1766465.792244 chr10 49104928 N chr10 49105224 N DUP 5
SRR1766473.10797123 chr10 49105274 N chr10 49105359 N DEL 5
SRR1766442.30169593 chr10 49104982 N chr10 49105188 N DEL 2
SRR1766453.10336138 chr10 49104978 N chr10 49105184 N DEL 7
SRR1766477.10830749 chr10 49104978 N chr10 49105184 N DEL 7
SRR1766461.10068879 chr10 49104979 N chr10 49105185 N DEL 7
SRR1766468.1748711 chr10 49104984 N chr10 49105190 N DEL 7
SRR1766458.3279031 chr10 49105335 N chr10 49105422 N DUP 9
SRR1766485.1266714 chr10 49105117 N chr10 49105341 N DEL 3
SRR1766478.6787392 chr10 49105380 N chr10 49105486 N DUP 3
SRR1766486.1036844 chr15 101763544 N chr15 101763731 N DUP 5
SRR1766447.2750525 chr15 101763550 N chr15 101763737 N DUP 8
SRR1766483.7404021 chr15 101763553 N chr15 101763740 N DUP 5
SRR1766473.5023340 chr15 101763542 N chr15 101763634 N DEL 10
SRR1766471.4159492 chr15 101763538 N chr15 101763816 N DUP 10
SRR1766478.2321437 chr15 101763529 N chr15 101763898 N DUP 5
SRR1766451.1635891 chr15 101763789 N chr15 101763881 N DEL 5
SRR1766463.5347317 chr15 101763733 N chr15 101763979 N DUP 5
SRR1766442.13863827 chr15 101763726 N chr15 101763972 N DUP 5
SRR1766478.11492364 chr15 101763733 N chr15 101763979 N DUP 5
SRR1766445.9509672 chr15 101763733 N chr15 101763979 N DUP 5
SRR1766478.6369112 chr15 101763733 N chr15 101763979 N DUP 5
SRR1766480.168118 chr15 101763771 N chr15 101764017 N DUP 4
SRR1766444.3613729 chr15 101763835 N chr15 101763990 N DUP 15
SRR1766461.7482410 chr15 101763700 N chr15 101764037 N DUP 7
SRR1766467.839787 chr15 101763552 N chr15 101763923 N DEL 5
SRR1766456.2068414 chr15 101763557 N chr15 101763928 N DEL 5
SRR1766457.8535198 chr15 101763708 N chr15 101764045 N DUP 15
SRR1766442.5056389 chr11 50210445 N chr11 50210506 N DEL 7
SRR1766445.4550658 chr11 50210445 N chr11 50210506 N DEL 7
SRR1766476.8083468 chr2 91411569 N chr2 91411720 N DEL 12
SRR1766457.6475972 chr2 91411569 N chr2 91411720 N DEL 14
SRR1766482.7385798 chr2 91411561 N chr2 91411637 N DEL 15
SRR1766442.9203551 chr2 91411561 N chr2 91411637 N DEL 16
SRR1766442.5604741 chr2 91411561 N chr2 91411637 N DEL 16
SRR1766455.9284697 chr2 91411477 N chr2 91411623 N DUP 9
SRR1766473.5844795 chr2 91411478 N chr2 91411725 N DUP 5
SRR1766446.9040484 chr2 91411600 N chr2 91411653 N DEL 4
SRR1766465.9461494 chr2 91411600 N chr2 91411653 N DEL 4
SRR1766472.1173620 chr2 91411600 N chr2 91411653 N DEL 3
SRR1766442.8615401 chr2 91411589 N chr2 91411642 N DEL 14
SRR1766442.28051979 chr2 91411589 N chr2 91411642 N DEL 14
SRR1766442.45350726 chr2 91411600 N chr2 91411653 N DEL 10
SRR1766471.6464001 chr2 91411600 N chr2 91411653 N DEL 8
SRR1766450.9897887 chr2 91411600 N chr2 91411653 N DEL 11
SRR1766456.5372149 chr2 91411600 N chr2 91411653 N DEL 12
SRR1766462.84490 chr2 91411600 N chr2 91411653 N DEL 12
SRR1766442.474109 chr13 99620946 N chr13 99620995 N DUP 10
SRR1766464.5004418 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766464.1312386 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766462.11166545 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766470.8699690 chr10 58708156 N chr10 58708299 N DEL 16
SRR1766454.8558581 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766472.11610492 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766443.4177231 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766449.3936321 chr10 58708156 N chr10 58708299 N DEL 17
SRR1766453.10001715 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766445.2605719 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766449.1496577 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766449.2454599 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766484.5634435 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766449.4918813 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766460.10997639 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766463.6155653 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766456.836855 chr10 58708270 N chr10 58708419 N DEL 5
SRR1766460.5763000 chr10 58708123 N chr10 58708419 N DEL 5
SRR1766466.3143481 chr10 58708123 N chr10 58708419 N DEL 5
SRR1766457.7199640 chr10 58708124 N chr10 58708420 N DEL 5
SRR1766486.7492795 chr10 58708132 N chr10 58708428 N DEL 5
SRR1766470.4263651 chr10 58708135 N chr10 58708431 N DEL 3
SRR1766473.2168284 chr6 36363978 N chr6 36364139 N DEL 5
SRR1766483.2040401 chr6 36364101 N chr6 36364262 N DEL 10
SRR1766442.20972254 chr13 18468131 N chr13 18469131 N DEL 3
SRR1766442.32226422 chr13 18468158 N chr13 18469156 N DUP 5
SRR1766449.942050 chr13 18468158 N chr13 18469156 N DUP 5
SRR1766476.476450 chr13 18468158 N chr13 18469156 N DUP 5
SRR1766465.1168276 chr13 18468160 N chr13 18469158 N DUP 5
SRR1766485.10527728 chr13 18468275 N chr13 18469696 N DEL 5
SRR1766447.4917925 chr13 18468275 N chr13 18469696 N DEL 5
SRR1766472.8655288 chr13 18468293 N chr13 18469712 N DUP 1
SRR1766469.4749135 chr13 18468405 N chr13 18468985 N DEL 9
SRR1766451.10072901 chr13 18468465 N chr13 18469633 N DEL 5
SRR1766464.613337 chr13 18468465 N chr13 18469633 N DEL 5
SRR1766451.10040829 chr13 18468465 N chr13 18469633 N DEL 5
SRR1766463.7256560 chr13 18468465 N chr13 18469633 N DEL 5
SRR1766449.942050 chr13 18468425 N chr13 18469003 N DUP 5
SRR1766471.12209535 chr13 18468425 N chr13 18469003 N DUP 5
SRR1766476.7742735 chr13 18468425 N chr13 18469003 N DUP 5
SRR1766462.9939431 chr13 18468425 N chr13 18469003 N DUP 5
SRR1766472.8549226 chr13 18468425 N chr13 18469003 N DUP 5
SRR1766476.225344 chr13 18468425 N chr13 18469003 N DUP 5
SRR1766456.4556662 chr13 18468425 N chr13 18469003 N DUP 8
SRR1766444.5727483 chr13 18468425 N chr13 18469003 N DUP 7
SRR1766447.348021 chr13 18468439 N chr13 18469437 N DUP 1
SRR1766477.10703311 chr13 18468484 N chr13 18469650 N DUP 4
SRR1766480.6019018 chr13 18469113 N chr13 18469450 N DEL 5
SRR1766464.1184363 chr13 18468490 N chr13 18469070 N DEL 5
SRR1766449.5793786 chr13 18468420 N chr13 18469084 N DEL 14
SRR1766451.4962205 chr13 18468491 N chr13 18469575 N DEL 5
SRR1766452.7664534 chr13 18468491 N chr13 18469575 N DEL 5
SRR1766447.5459916 chr13 18468574 N chr13 18469576 N DEL 5
SRR1766464.496106 chr13 18468325 N chr13 18469827 N DUP 3
SRR1766449.9118484 chr10 83585241 N chr10 83585319 N DEL 31
SRR1766484.2236619 chr10 83585233 N chr10 83585348 N DUP 21
SRR1766446.2853833 chr10 83585201 N chr10 83585311 N DUP 2
SRR1766445.3062325 chr10 83585215 N chr10 83585292 N DEL 9
SRR1766461.10657587 chr10 83585215 N chr10 83585292 N DEL 9
SRR1766479.7061399 chr10 83585215 N chr10 83585312 N DEL 13
SRR1766443.4056017 chr10 83585260 N chr10 83585312 N DEL 19
SRR1766465.9769986 chr10 83585215 N chr10 83585312 N DEL 12
SRR1766447.9802070 chr10 83585216 N chr10 83585313 N DEL 12
SRR1766472.9956458 chr10 83585264 N chr10 83585316 N DEL 11
SRR1766478.3536599 chr10 83585266 N chr10 83585318 N DEL 9
SRR1766443.3331832 chr10 114737114 N chr10 114737248 N DUP 2
SRR1766446.6989397 chr4 45024481 N chr4 45024572 N DUP 5
SRR1766449.3355157 chr4 45024483 N chr4 45024574 N DUP 5
SRR1766460.10986091 chr4 45024485 N chr4 45024576 N DUP 5
SRR1766467.10819439 chr4 45024485 N chr4 45024576 N DUP 5
SRR1766473.3499570 chr4 45024485 N chr4 45024576 N DUP 5
SRR1766442.35752459 chr4 45024486 N chr4 45024605 N DUP 5
SRR1766463.6022293 chr4 45024702 N chr4 45024763 N DEL 3
SRR1766446.2834015 chr17 41123840 N chr17 41123916 N DEL 4
SRR1766453.6951404 chr17 41124011 N chr17 41124132 N DEL 2
SRR1766445.5609964 chr17 41124012 N chr17 41124133 N DEL 3
SRR1766476.5739410 chr17 41124011 N chr17 41124132 N DEL 4
SRR1766453.3959204 chr17 41124011 N chr17 41124132 N DEL 5
SRR1766469.1381832 chr17 41124059 N chr17 41124180 N DEL 5
SRR1766475.10768449 chr17 41124060 N chr17 41124179 N DUP 5
SRR1766482.4584152 chr17 41123984 N chr17 41124105 N DEL 7
SRR1766464.7738294 chr17 41123984 N chr17 41124105 N DEL 6
SRR1766480.4128761 chr17 41123864 N chr17 41124105 N DEL 5
SRR1766467.11122595 chr17 41123891 N chr17 41124132 N DEL 10
SRR1766469.5487914 chr17 41123891 N chr17 41124132 N DEL 10
SRR1766453.8800494 chr17 41123891 N chr17 41124132 N DEL 10
SRR1766454.218979 chr17 41123891 N chr17 41124132 N DEL 10
SRR1766478.669465 chr17 41123891 N chr17 41124132 N DEL 9
SRR1766453.1220644 chr17 41123891 N chr17 41124132 N DEL 5
SRR1766483.5898113 chr17 41123891 N chr17 41124132 N DEL 5
SRR1766477.10070576 chr2 233035819 N chr2 233035886 N DUP 7
SRR1766449.6559513 chr7 61803568 N chr7 61803908 N DUP 5
SRR1766442.10733765 chr7 61803716 N chr7 61803886 N DUP 5
SRR1766475.10595440 chr7 61803545 N chr7 61804393 N DEL 5
SRR1766456.5814328 chr13 27748106 N chr13 27748267 N DEL 5
SRR1766445.7527746 chr13 27748144 N chr13 27748305 N DEL 1
SRR1766481.5581138 chr13 27747910 N chr13 27748188 N DUP 5
SRR1766474.9424075 chr17 10475742 N chr17 10475797 N DUP 19
SRR1766455.5567930 chr7 111539297 N chr7 111539354 N DEL 15
SRR1766473.4109352 chr21 40364843 N chr21 40364910 N DUP 6
SRR1766466.39818 chr14 47139953 N chr14 47140010 N DEL 5
SRR1766463.1755430 chr19 53559050 N chr19 53559157 N DUP 17
SRR1766475.5827848 chr19 53559050 N chr19 53559157 N DUP 16
SRR1766482.11081530 chr19 53559050 N chr19 53559157 N DUP 16
SRR1766465.10807234 chr19 53559064 N chr19 53559241 N DUP 1
SRR1766464.7735615 chr19 53559021 N chr19 53559104 N DEL 8
SRR1766445.6110651 chr19 53559022 N chr19 53559105 N DEL 8
SRR1766443.8981208 chr19 53559024 N chr19 53559107 N DEL 6
SRR1766480.7428873 chr19 53559229 N chr19 53559348 N DEL 7
SRR1766442.41474231 chr19 53559226 N chr19 53559343 N DUP 5
SRR1766481.1530174 chr19 53559272 N chr19 53559387 N DUP 5
SRR1766477.6875400 chr19 53559281 N chr19 53559398 N DUP 5
SRR1766483.7102010 chr19 53559022 N chr19 53559300 N DEL 3
SRR1766443.4797883 chr1 191828617 N chr1 191828736 N DEL 14
SRR1766452.8612104 chr1 191828611 N chr1 191828736 N DEL 14
SRR1766466.5250270 chr1 191828611 N chr1 191828738 N DEL 13
SRR1766450.1975808 chr8 14847784 N chr8 14847891 N DUP 5
SRR1766450.10077471 chr12 131247281 N chr12 131247393 N DEL 2
SRR1766480.6065734 chr22 32329737 N chr22 32330066 N DEL 2
SRR1766446.8077423 chr22 32329947 N chr22 32331286 N DEL 1
SRR1766456.5063869 chr22 32329881 N chr22 32330167 N DUP 21
SRR1766456.311475 chr22 32330193 N chr22 32330414 N DUP 6
SRR1766443.1483676 chr22 32329781 N chr22 32330227 N DEL 1
SRR1766442.12898336 chr22 32330421 N chr22 32330861 N DEL 1
SRR1766461.3313195 chr22 32330694 N chr22 32330952 N DEL 10
SRR1766445.7399666 chr22 32329857 N chr22 32330695 N DEL 6
SRR1766481.1735460 chr22 32329729 N chr22 32330695 N DEL 8
SRR1766453.10923412 chr22 32329787 N chr22 32330928 N DUP 5
SRR1766455.2442462 chr22 32330065 N chr22 32330918 N DUP 1
SRR1766453.9584636 chr22 32330717 N chr22 32330985 N DUP 5
SRR1766477.169762 chr22 32329804 N chr22 32331093 N DUP 5
SRR1766469.7646005 chr22 32330227 N chr22 32331116 N DUP 10
SRR1766451.4648276 chr22 32330057 N chr22 32331102 N DUP 5
SRR1766484.3511511 chr22 32330744 N chr22 32331014 N DEL 11
SRR1766456.2004508 chr22 32331018 N chr22 32331093 N DUP 5
SRR1766447.7705951 chr22 32330050 N chr22 32331116 N DUP 5
SRR1766451.6534568 chr22 32330100 N chr22 32331304 N DEL 29
SRR1766452.4833591 chr22 32329821 N chr22 32331337 N DEL 11
SRR1766473.6322467 chr19 33536496 N chr19 33536553 N DUP 5
SRR1766466.28321 chr20 57453562 N chr20 57453872 N DEL 3
SRR1766483.1473463 chr20 61444892 N chr20 61445029 N DEL 5
SRR1766471.10757781 chr13 84125790 N chr13 84125882 N DUP 10
SRR1766467.11087533 chr13 84125842 N chr13 84126007 N DUP 5
SRR1766460.1761163 chr13 111197272 N chr13 111197409 N DUP 1
SRR1766442.2890192 chr13 111197272 N chr13 111197409 N DUP 1
SRR1766476.3006525 chr13 111197294 N chr13 111197433 N DEL 5
SRR1766451.9845037 chr13 111197294 N chr13 111197433 N DEL 5
SRR1766480.7970230 chr13 111197294 N chr13 111197433 N DEL 5
SRR1766456.5689171 chr13 111197299 N chr13 111197438 N DEL 5
SRR1766464.10636960 chr10 110411892 N chr10 110411965 N DUP 7
SRR1766478.4536335 chr10 110411897 N chr10 110412044 N DUP 9
SRR1766442.18914588 chr10 110411888 N chr10 110411961 N DUP 6
SRR1766450.5530687 chr10 110411888 N chr10 110411961 N DUP 13
SRR1766459.7854122 chr10 110411971 N chr10 110412044 N DUP 5
SRR1766451.9033452 chr9 89671689 N chr9 89671819 N DEL 18
SRR1766461.6554851 chr9 89671689 N chr9 89671819 N DEL 32
SRR1766483.11646071 chr9 89671698 N chr9 89671748 N DUP 15
SRR1766442.15415282 chr9 89671740 N chr9 89671895 N DUP 15
SRR1766450.81952 chr9 89671770 N chr9 89671826 N DUP 19
SRR1766472.9302579 chr9 89671769 N chr9 89671819 N DUP 1
SRR1766483.186203 chr9 89671770 N chr9 89671877 N DUP 17
SRR1766442.27168270 chr9 89671692 N chr9 89671871 N DUP 20
SRR1766453.6777803 chr9 89671710 N chr9 89671868 N DUP 27
SRR1766465.3894362 chr9 89671698 N chr9 89671808 N DUP 18
SRR1766442.43397043 chr9 89671656 N chr9 89671793 N DUP 13
SRR1766460.5257654 chr9 89671713 N chr9 89671871 N DUP 6
SRR1766442.31375677 chr9 89671738 N chr9 89671923 N DUP 10
SRR1766442.34575855 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766483.2545094 chr9 89671664 N chr9 89671825 N DUP 6
SRR1766453.6777803 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766471.11994022 chr9 89671710 N chr9 89671781 N DUP 9
SRR1766442.3282057 chr9 89671713 N chr9 89671769 N DUP 17
SRR1766474.9109956 chr9 89671692 N chr9 89671802 N DUP 14
SRR1766455.4344450 chr9 89671692 N chr9 89671937 N DUP 23
SRR1766468.7418887 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766462.6278994 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766467.648867 chr9 89671742 N chr9 89671945 N DUP 10
SRR1766460.2499286 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766482.10510174 chr9 89671701 N chr9 89671850 N DUP 15
SRR1766479.889896 chr9 89671755 N chr9 89671859 N DUP 12
SRR1766445.3147857 chr9 89671755 N chr9 89671859 N DUP 12
SRR1766472.10619239 chr9 89671713 N chr9 89671769 N DUP 17
SRR1766464.1845413 chr9 89671770 N chr9 89671877 N DUP 20
SRR1766473.5048874 chr9 89671713 N chr9 89671871 N DUP 27
SRR1766458.2726627 chr9 89671692 N chr9 89671802 N DUP 14
SRR1766481.97153 chr9 89671770 N chr9 89671826 N DUP 23
SRR1766459.10678798 chr9 89671692 N chr9 89671837 N DUP 24
SRR1766455.1511834 chr9 89671818 N chr9 89671874 N DUP 22
SRR1766475.9514433 chr9 89671772 N chr9 89671849 N DUP 20
SRR1766473.5048874 chr9 89671770 N chr9 89671877 N DUP 24
SRR1766468.6203617 chr9 89671729 N chr9 89671782 N DUP 16
SRR1766453.4804902 chr9 89671692 N chr9 89671802 N DUP 19
SRR1766442.36499330 chr9 89671729 N chr9 89671833 N DUP 10
SRR1766460.6361669 chr9 89671729 N chr9 89671833 N DUP 15
SRR1766472.1245181 chr9 89671771 N chr9 89671878 N DUP 17
SRR1766450.7868999 chr9 89671729 N chr9 89671833 N DUP 23
SRR1766470.5022487 chr9 89671692 N chr9 89671802 N DUP 19
SRR1766442.21049350 chr9 89671676 N chr9 89671749 N DEL 6
SRR1766466.8258181 chr9 89671676 N chr9 89671749 N DEL 6
SRR1766484.3901896 chr9 89671729 N chr9 89671782 N DUP 15
SRR1766471.11994022 chr9 89671701 N chr9 89671859 N DUP 17
SRR1766473.6578963 chr9 89671698 N chr9 89671775 N DUP 17
SRR1766481.10663315 chr9 89671770 N chr9 89671877 N DUP 22
SRR1766473.8097852 chr9 89671680 N chr9 89671753 N DEL 2
SRR1766450.5021997 chr9 89671692 N chr9 89671802 N DUP 23
SRR1766463.633447 chr9 89671781 N chr9 89671936 N DUP 8
SRR1766475.9199244 chr9 89671753 N chr9 89671884 N DUP 2
SRR1766486.7288799 chr9 89671753 N chr9 89671884 N DUP 3
SRR1766466.9088531 chr9 89671701 N chr9 89671859 N DUP 19
SRR1766471.2137093 chr9 89671705 N chr9 89671812 N DUP 10
SRR1766447.2003579 chr9 89671692 N chr9 89671853 N DUP 11
SRR1766478.9056447 chr9 89671770 N chr9 89671877 N DUP 26
SRR1766450.1914612 chr9 89671792 N chr9 89671878 N DUP 12
SRR1766483.8401693 chr9 89671818 N chr9 89671874 N DUP 19
SRR1766449.1978826 chr9 89671818 N chr9 89671874 N DUP 27
SRR1766457.3867954 chr9 89671720 N chr9 89671793 N DEL 12
SRR1766471.4303433 chr9 89671738 N chr9 89671893 N DUP 24
SRR1766447.10681820 chr9 89671690 N chr9 89671935 N DUP 17
SRR1766442.17130031 chr9 89671743 N chr9 89671841 N DUP 12
SRR1766462.9338154 chr9 89671675 N chr9 89671778 N DEL 7
SRR1766447.443044 chr9 89671770 N chr9 89671877 N DUP 28
SRR1766482.5794508 chr9 89671692 N chr9 89671853 N DUP 31
SRR1766476.10484931 chr9 89671724 N chr9 89671818 N DEL 5
SRR1766462.9665532 chr9 89671864 N chr9 89671932 N DUP 5
SRR1766461.10271180 chr9 89671734 N chr9 89671843 N DEL 5
SRR1766456.5141629 chr9 89671829 N chr9 89671881 N DEL 10
SRR1766485.3052228 chr9 89671724 N chr9 89671884 N DEL 12
SRR1766462.9256981 chr9 89671766 N chr9 89671890 N DEL 5
SRR1766442.10108642 chr9 89671767 N chr9 89671891 N DEL 4
SRR1766460.2093877 chr9 89671678 N chr9 89671904 N DEL 1
SRR1766472.3515691 chr9 89671871 N chr9 89671923 N DEL 8
SRR1766477.1372195 chr9 89671673 N chr9 89671935 N DEL 3
SRR1766455.3042337 chr6 89125587 N chr6 89126778 N DEL 4
SRR1766478.748849 chr6 89125628 N chr6 89125934 N DEL 5
SRR1766474.6189546 chr6 89125640 N chr6 89125944 N DUP 9
SRR1766452.2872880 chr6 89126071 N chr6 89126670 N DEL 3
SRR1766444.4934578 chr6 89125933 N chr6 89126832 N DUP 11
SRR1766442.31832656 chr6 89125947 N chr6 89126831 N DEL 2
SRR1766479.6714728 chr1 207315826 N chr1 207315923 N DEL 5
SRR1766471.10456104 chr1 207315729 N chr1 207315818 N DEL 7
SRR1766442.30039505 chr1 207315772 N chr1 207315827 N DEL 5
SRR1766449.5469315 chr1 207315767 N chr1 207315892 N DEL 2
SRR1766462.8922206 chr1 207315827 N chr1 207315944 N DEL 3
SRR1766472.4939874 chr13 52818024 N chr13 52818451 N DEL 7
SRR1766469.8335865 chr13 52818046 N chr13 52818471 N DUP 9
SRR1766456.6423839 chr13 52818047 N chr13 52818472 N DUP 8
SRR1766453.7115105 chr13 52818165 N chr13 52818474 N DUP 5
SRR1766469.7369787 chr22 48858033 N chr22 48858232 N DUP 5
SRR1766483.10634864 chr22 48857991 N chr22 48858042 N DEL 9
SRR1766443.9191301 chr22 48858144 N chr22 48858243 N DUP 10
SRR1766465.1487523 chr22 48858144 N chr22 48858193 N DUP 5
SRR1766442.33948611 chr22 48858144 N chr22 48858193 N DUP 5
SRR1766460.1206443 chr22 48858137 N chr22 48858236 N DUP 5
SRR1766479.11356186 chr22 48858137 N chr22 48858236 N DUP 5
SRR1766467.4395583 chr22 48858141 N chr22 48858240 N DUP 5
SRR1766459.3947627 chr22 48858144 N chr22 48858193 N DUP 5
SRR1766455.4443474 chr22 48858009 N chr22 48858160 N DEL 5
SRR1766442.17217561 chr13 92297394 N chr13 92297555 N DEL 5
SRR1766463.7196809 chr22 36434243 N chr22 36434385 N DUP 12
SRR1766474.7663017 chr22 36434342 N chr22 36434399 N DUP 22
SRR1766458.1222399 chr22 36434323 N chr22 36434386 N DUP 10
SRR1766442.4509105 chr22 36434260 N chr22 36434359 N DEL 10
SRR1766478.6579743 chr22 36434260 N chr22 36434359 N DEL 10
SRR1766450.7669133 chr22 36434248 N chr22 36434375 N DEL 8
SRR1766483.10563390 chr1 5804559 N chr1 5804714 N DUP 2
SRR1766454.1096888 chr1 96153244 N chr1 96153309 N DUP 3
SRR1766476.6618191 chr1 96153244 N chr1 96153309 N DUP 5
SRR1766477.198242 chr1 96153244 N chr1 96153309 N DUP 5
SRR1766448.9788747 chr1 96153244 N chr1 96153309 N DUP 25
SRR1766450.8675057 chr1 96153244 N chr1 96153309 N DUP 32
SRR1766444.6197180 chr1 96153244 N chr1 96153309 N DUP 30
SRR1766445.10309417 chr1 96153244 N chr1 96153309 N DUP 29
SRR1766481.11244748 chr1 96153244 N chr1 96153309 N DUP 25
SRR1766455.93041 chr1 96153244 N chr1 96153309 N DUP 8
SRR1766443.9470226 chr1 96153244 N chr1 96153309 N DUP 25
SRR1766442.9972324 chr1 96153244 N chr1 96153309 N DUP 25
SRR1766475.5016149 chr1 96153244 N chr1 96153309 N DUP 23
SRR1766477.7379421 chr1 96153244 N chr1 96153309 N DUP 12
SRR1766481.6612261 chr1 96153244 N chr1 96153309 N DUP 13
SRR1766442.24511617 chr1 96153244 N chr1 96153309 N DUP 19
SRR1766448.3634630 chr1 96153244 N chr1 96153309 N DUP 18
SRR1766463.3962757 chr1 96153244 N chr1 96153309 N DUP 18
SRR1766476.10068121 chr1 96153244 N chr1 96153309 N DUP 20
SRR1766456.1000680 chr1 96153244 N chr1 96153309 N DUP 7
SRR1766453.867901 chr1 96153252 N chr1 96153317 N DUP 5
SRR1766482.12656170 chr1 96153244 N chr1 96153309 N DUP 26
SRR1766471.11558901 chr1 96153244 N chr1 96153309 N DUP 30
SRR1766479.8424729 chr1 96153244 N chr1 96153309 N DUP 30
SRR1766483.10966137 chr1 96153237 N chr1 96153329 N DEL 9
SRR1766456.5549548 chrX 143492665 N chrX 143492759 N DEL 10
SRR1766484.10336819 chr11 82625107 N chr11 82625168 N DUP 4
SRR1766443.10808698 chr11 82625189 N chr11 82625252 N DEL 5
SRR1766445.9449135 chr11 82625189 N chr11 82625252 N DEL 5
SRR1766486.164433 chr11 82625189 N chr11 82625252 N DEL 5
SRR1766478.2733615 chr11 82625189 N chr11 82625252 N DEL 5
SRR1766457.7135441 chr11 82625158 N chr11 82625252 N DEL 5
SRR1766479.11249282 chr11 82625158 N chr11 82625252 N DEL 5
SRR1766452.4779377 chr11 82625158 N chr11 82625252 N DEL 5
SRR1766442.2915091 chr11 82625174 N chr11 82625609 N DEL 6
SRR1766485.1103097 chr11 82625158 N chr11 82625252 N DEL 5
SRR1766485.6845551 chr11 82625143 N chr11 82625578 N DEL 7
SRR1766470.1526638 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766442.26159733 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766457.4828538 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766466.5100626 chr11 82625639 N chr11 82625700 N DUP 5
SRR1766446.5275326 chr11 82625144 N chr11 82625298 N DEL 5
SRR1766461.7208748 chr11 82625144 N chr11 82625298 N DEL 5
SRR1766443.1243459 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766454.9923865 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766467.1150909 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766467.10006278 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766471.3995506 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766481.5327801 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766466.2465400 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766464.3919215 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766454.1319920 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766469.1075203 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766475.7121725 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766479.1857319 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766485.9433274 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766471.9509743 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766479.919869 chr11 82625144 N chr11 82625298 N DEL 5
SRR1766447.615898 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766476.1429636 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766456.5622208 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766461.8878019 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766472.1657650 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766479.8296166 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766473.10714094 chr11 82625268 N chr11 82625701 N DUP 5
SRR1766452.10027210 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766446.2667981 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766474.6858171 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766449.1384187 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766460.4451839 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766448.6009477 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766449.5443472 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766453.3937140 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766442.27603532 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766475.10552943 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766470.4046916 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766458.2836886 chr11 82625268 N chr11 82625577 N DEL 5
SRR1766442.32875246 chr11 82625268 N chr11 82625577 N DEL 5
SRR1766470.2401346 chr11 82625268 N chr11 82625577 N DEL 5
SRR1766445.3944385 chr11 82625239 N chr11 82625701 N DUP 11
SRR1766484.10336819 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766442.23272736 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766451.8943180 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766448.4917194 chr11 82625239 N chr11 82625701 N DUP 12
SRR1766471.660448 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766479.1857319 chr11 82625144 N chr11 82625298 N DEL 5
SRR1766450.2529431 chr11 82625268 N chr11 82625639 N DEL 15
SRR1766479.7871069 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766450.8302904 chr11 82625298 N chr11 82625700 N DUP 5
SRR1766481.5327801 chr11 82625144 N chr11 82625298 N DEL 5
SRR1766471.3810130 chr11 82625144 N chr11 82625298 N DEL 5
SRR1766447.615898 chr11 82625268 N chr11 82625701 N DUP 5
SRR1766461.10958631 chr11 82625086 N chr11 82625776 N DEL 8
SRR1766449.9895207 chr5 58889084 N chr5 58889192 N DUP 7
SRR1766466.9561632 chr7 26620013 N chr7 26620157 N DEL 4
SRR1766470.10170800 chr1 67930134 N chr1 67930185 N DEL 16
SRR1766442.28711279 chr1 67930132 N chr1 67930188 N DEL 12
SRR1766459.4334118 chr1 67930132 N chr1 67930188 N DEL 12
SRR1766442.36425228 chr1 67930133 N chr1 67930189 N DEL 11
SRR1766448.2886559 chr1 67930133 N chr1 67930194 N DEL 6
SRR1766468.7320823 chr1 67930133 N chr1 67930194 N DEL 6
SRR1766473.7086936 chr1 67930134 N chr1 67930195 N DEL 5
SRR1766480.5814775 chr1 67930133 N chr1 67930199 N DEL 1
SRR1766452.10494590 chr9 129075407 N chr9 129075538 N DUP 3
SRR1766457.1770646 chr9 129075426 N chr9 129075559 N DEL 5
SRR1766442.46399505 chr9 129075433 N chr9 129075566 N DEL 5
SRR1766453.453629 chr6 64296679 N chr6 64296774 N DEL 13
SRR1766474.10119312 chr6 64296679 N chr6 64296774 N DEL 13
SRR1766442.30041039 chr18 79631201 N chr18 79631557 N DEL 1
SRR1766485.9274433 chr18 79631238 N chr18 79631421 N DEL 5
SRR1766442.31667097 chr18 79631143 N chr18 79631305 N DUP 10
SRR1766455.9012160 chr18 79631217 N chr18 79631408 N DUP 2
SRR1766442.299375 chr18 79631096 N chr18 79631349 N DEL 3
SRR1766468.4850778 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766463.3065180 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766472.12030894 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766482.6565003 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766459.2999629 chr20 22378545 N chr20 22378668 N DEL 10
SRR1766474.1018088 chr20 22378591 N chr20 22378658 N DEL 14
SRR1766442.4714973 chr20 22378591 N chr20 22378658 N DEL 15
SRR1766448.10370720 chr20 22378581 N chr20 22378638 N DEL 15
SRR1766463.7254966 chr20 22378615 N chr20 22378744 N DEL 12
SRR1766479.11251285 chr20 22378581 N chr20 22378638 N DEL 20
SRR1766469.8627368 chr20 22378581 N chr20 22378638 N DEL 25
SRR1766443.6222788 chr20 22378605 N chr20 22378730 N DUP 5
SRR1766447.6572847 chr20 21537794 N chr20 21537865 N DEL 6
SRR1766444.6096505 chr20 21537813 N chr20 21537864 N DEL 7
SRR1766461.1932418 chr11 132162754 N chr11 132162869 N DUP 18
SRR1766465.10263446 chr11 132162725 N chr11 132162930 N DUP 4
SRR1766459.2603290 chr2 5172401 N chr2 5172504 N DUP 10
SRR1766446.8099319 chr2 5172521 N chr2 5172749 N DEL 1
SRR1766479.7833899 chr2 5172452 N chr2 5172521 N DUP 5
SRR1766477.2438837 chr2 5172521 N chr2 5172749 N DEL 8
SRR1766464.6095762 chr2 5172452 N chr2 5172521 N DUP 10
SRR1766474.10122045 chr2 5172452 N chr2 5172521 N DUP 5
SRR1766451.2656153 chr2 5172441 N chr2 5172667 N DUP 14
SRR1766464.6888983 chr2 5172375 N chr2 5172548 N DUP 5
SRR1766458.5366035 chr2 5172479 N chr2 5172548 N DUP 11
SRR1766481.8272481 chr2 5172511 N chr2 5172667 N DUP 5
SRR1766474.3278831 chr2 5172391 N chr2 5172566 N DEL 1
SRR1766456.5567803 chr2 5172391 N chr2 5172566 N DEL 1
SRR1766481.3273931 chr2 5172536 N chr2 5172624 N DEL 6
SRR1766478.2884598 chr2 5172404 N chr2 5172734 N DUP 5
SRR1766457.9502353 chr2 5172404 N chr2 5172734 N DUP 5
SRR1766466.3030116 chr2 5172375 N chr2 5172637 N DEL 5
SRR1766454.930909 chr2 5172406 N chr2 5172668 N DEL 5
SRR1766472.11983339 chr2 5172576 N chr2 5172681 N DEL 3
SRR1766464.5250533 chr2 5172442 N chr2 5172738 N DUP 13
SRR1766485.7867618 chr2 5172442 N chr2 5172738 N DUP 14
SRR1766458.5405039 chr2 5172712 N chr2 5172781 N DUP 5
SRR1766482.7999140 chr2 5172442 N chr2 5172738 N DUP 15
SRR1766468.4452065 chr2 5172439 N chr2 5172701 N DEL 5
SRR1766456.5749530 chr2 5172749 N chr2 5172818 N DUP 5
SRR1766465.611496 chr2 5172457 N chr2 5172823 N DUP 5
SRR1766465.4066721 chr2 5172453 N chr2 5172819 N DUP 10
SRR1766466.10070456 chr2 5172457 N chr2 5172823 N DUP 5
SRR1766455.6003896 chr2 5172457 N chr2 5172823 N DUP 5
SRR1766465.3727250 chr2 5172457 N chr2 5172823 N DUP 5
SRR1766456.1598082 chr7 66231173 N chr7 66231334 N DEL 5
SRR1766467.10739014 chr7 66231134 N chr7 66231295 N DEL 5
SRR1766463.5796289 chr4 149047120 N chr4 149047347 N DEL 3
SRR1766446.4855979 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766442.26025961 chr4 149047120 N chr4 149047347 N DEL 6
SRR1766481.220266 chr4 149047120 N chr4 149047347 N DEL 7
SRR1766442.13367979 chr4 149047120 N chr4 149047347 N DEL 7
SRR1766455.2447653 chr4 149047120 N chr4 149047347 N DEL 7
SRR1766479.3624000 chr4 149047120 N chr4 149047347 N DEL 7
SRR1766442.36615782 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766471.7468403 chr4 149047120 N chr4 149047347 N DEL 7
SRR1766442.38688191 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766442.17467967 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766442.35403156 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766470.8640406 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766461.6322797 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766449.4493670 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766442.21808024 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766482.1410844 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766482.2039014 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766442.18317366 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766459.6210399 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766467.9952947 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766459.8065812 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766475.4821277 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766484.4940572 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766486.9936453 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766459.1247659 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766483.10996278 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766442.22343347 chr4 149047088 N chr4 149047347 N DEL 7
SRR1766474.2603167 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766453.10069926 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766485.10570042 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766481.4877153 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766446.1145365 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766459.10052551 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766471.6713084 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766442.30046645 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766467.8022230 chr4 149047056 N chr4 149047347 N DEL 7
SRR1766447.3939850 chr4 149047030 N chr4 149047353 N DEL 7
SRR1766448.9531825 chr7 72255251 N chr7 72255555 N DUP 4
SRR1766467.375395 chr7 72255269 N chr7 72255599 N DEL 20
SRR1766470.10878154 chr4 1652179 N chr4 1652707 N DEL 5
SRR1766471.5715339 chr4 1652203 N chr4 1652384 N DEL 7
SRR1766478.6416402 chr4 1652212 N chr4 1652711 N DEL 15
SRR1766483.10468105 chr4 1652233 N chr4 1652733 N DEL 12
SRR1766460.10149699 chr4 1652251 N chr4 1653072 N DEL 8
SRR1766444.3148256 chr4 1652332 N chr4 1652384 N DEL 10
SRR1766452.8202823 chr4 1652204 N chr4 1652350 N DUP 9
SRR1766455.2767194 chr4 1652164 N chr4 1652350 N DUP 9
SRR1766445.862033 chr4 1652305 N chr4 1652427 N DUP 3
SRR1766472.5122422 chr4 1652379 N chr4 1652875 N DUP 9
SRR1766447.183552 chr4 1652525 N chr4 1652579 N DEL 7
SRR1766464.4990011 chr4 1652362 N chr4 1652543 N DUP 9
SRR1766450.10170017 chr4 1652285 N chr4 1652595 N DUP 12
SRR1766475.8899743 chr4 1652615 N chr4 1653151 N DEL 1
SRR1766479.1077914 chr4 1652198 N chr4 1652585 N DEL 5
SRR1766468.5748843 chr4 1652573 N chr4 1652740 N DUP 3
SRR1766442.43087218 chr4 1652299 N chr4 1652627 N DEL 9
SRR1766479.4628079 chr4 1652631 N chr4 1653165 N DUP 6
SRR1766442.32025554 chr4 1652385 N chr4 1652752 N DUP 11
SRR1766475.8193333 chr4 1652624 N chr4 1652788 N DUP 12
SRR1766442.20982458 chr4 1652791 N chr4 1652929 N DEL 11
SRR1766470.2492378 chr4 1652144 N chr4 1652934 N DUP 5
SRR1766444.168556 chr4 1652837 N chr4 1653019 N DUP 5
SRR1766448.8707697 chr4 1652301 N chr4 1652908 N DEL 1
SRR1766482.8155477 chr4 1652928 N chr4 1653363 N DUP 8
SRR1766482.8965201 chr4 1652601 N chr4 1652972 N DEL 22
SRR1766447.183552 chr4 1652197 N chr4 1652969 N DEL 6
SRR1766464.4990011 chr4 1653007 N chr4 1653276 N DUP 1
SRR1766486.5304800 chr4 1652852 N chr4 1653022 N DEL 1
SRR1766450.10170017 chr4 1652252 N chr4 1653126 N DEL 4
SRR1766471.11924537 chr4 1652321 N chr4 1653153 N DEL 5
SRR1766469.4785279 chr5 29743712 N chr5 29743790 N DUP 6
SRR1766477.5301882 chr5 29743712 N chr5 29743790 N DUP 12
SRR1766465.9281932 chr10 17629553 N chr10 17629750 N DEL 10
SRR1766465.4026573 chr10 17629449 N chr10 17629530 N DEL 1
SRR1766475.6868300 chr10 17629696 N chr10 17629853 N DEL 5
SRR1766481.1744450 chr7 116768118 N chr7 116768191 N DUP 8
SRR1766482.6212979 chr6 104424259 N chr6 104424392 N DEL 4
SRR1766459.6384534 chr6 104424259 N chr6 104424392 N DEL 7
SRR1766462.7797835 chr6 104424368 N chr6 104424501 N DEL 11
SRR1766463.5418275 chr6 104424259 N chr6 104424400 N DEL 25
SRR1766442.967555 chr6 104424329 N chr6 104424462 N DEL 18
SRR1766473.4522759 chr6 104424329 N chr6 104424462 N DEL 18
SRR1766445.8931811 chr6 104424329 N chr6 104424462 N DEL 18
SRR1766442.24393412 chr6 104424190 N chr6 104424475 N DEL 2
SRR1766445.1846767 chr6 104424332 N chr6 104424501 N DEL 5
SRR1766444.532132 chr6 104424448 N chr6 104424549 N DEL 16
SRR1766464.8385957 chr6 104424385 N chr6 104424566 N DEL 13
SRR1766485.9612350 chr6 104424385 N chr6 104424566 N DEL 13
SRR1766483.517225 chr6 104424385 N chr6 104424566 N DEL 13
SRR1766461.7506131 chr3 122780251 N chr3 122780350 N DEL 5
SRR1766457.1495452 chr3 122780252 N chr3 122780351 N DEL 10
SRR1766472.10202845 chr3 122780329 N chr3 122780427 N DUP 7
SRR1766460.2390377 chr3 122780285 N chr3 122780431 N DUP 5
SRR1766442.19190595 chr3 122780339 N chr3 122780388 N DUP 2
SRR1766477.673845 chr3 122780338 N chr3 122780389 N DEL 6
SRR1766478.1461263 chr3 122780291 N chr3 122780390 N DEL 5
SRR1766442.36034386 chr3 122780195 N chr3 122780565 N DUP 1
SRR1766474.5536027 chr3 122780195 N chr3 122780419 N DUP 3
SRR1766463.10429696 chr3 122780204 N chr3 122780574 N DUP 2
SRR1766486.6006713 chr3 122780273 N chr3 122780519 N DEL 5
SRR1766460.7475219 chr3 122780329 N chr3 122780649 N DUP 5
SRR1766473.2291270 chr3 122780276 N chr3 122780648 N DEL 5
SRR1766442.24341092 chr3 122780279 N chr3 122780651 N DEL 4
SRR1766486.4183173 chr3 122780546 N chr3 122780721 N DEL 10
SRR1766449.5453261 chr3 122780339 N chr3 122780806 N DUP 7
SRR1766481.332204 chr3 122780339 N chr3 122780806 N DUP 7
SRR1766483.6427839 chr3 122780546 N chr3 122780721 N DEL 15
SRR1766450.5770543 chr3 122780365 N chr3 122780833 N DEL 5
SRR1766477.6589296 chr3 181743074 N chr3 181743217 N DEL 16
SRR1766482.795057 chr3 181743062 N chr3 181743157 N DEL 15
SRR1766457.7759522 chr3 181743053 N chr3 181743112 N DUP 25
SRR1766481.2321111 chr15 84672847 N chr15 84672964 N DEL 3
SRR1766466.1381218 chr15 84672895 N chr15 84673012 N DEL 13
SRR1766486.6995240 chr15 84672963 N chr15 84673080 N DEL 5
SRR1766481.1943707 chr15 84672901 N chr15 84673210 N DUP 5
SRR1766447.4043922 chr15 84673061 N chr15 84673259 N DEL 6
SRR1766461.475316 chrY 10750602 N chrY 10750701 N DUP 10
SRR1766485.11627066 chrY 10750588 N chrY 10750724 N DEL 3
SRR1766447.5041538 chr19 108019 N chr19 108076 N DUP 12
SRR1766477.4433814 chr19 108019 N chr19 108076 N DUP 14
SRR1766447.1495805 chr19 108019 N chr19 108076 N DUP 20
SRR1766461.3872695 chr19 107980 N chr19 108037 N DUP 25
SRR1766462.8314030 chr19 108019 N chr19 108076 N DUP 23
SRR1766475.1018103 chr19 107980 N chr19 108037 N DUP 28
SRR1766458.3804696 chr19 108015 N chr19 108082 N DUP 3
SRR1766486.11960780 chr19 108015 N chr19 108082 N DUP 3
SRR1766464.1816599 chr19 108015 N chr19 108082 N DUP 8
SRR1766442.16085073 chr19 108015 N chr19 108082 N DUP 5
SRR1766464.4285568 chr19 108015 N chr19 108082 N DUP 6
SRR1766467.5463105 chr19 108015 N chr19 108082 N DUP 6
SRR1766458.3282239 chr19 108015 N chr19 108082 N DUP 10
SRR1766472.10946882 chr19 107980 N chr19 108081 N DUP 20
SRR1766461.7452503 chr19 107980 N chr19 108081 N DUP 22
SRR1766445.5725495 chr19 107980 N chr19 108081 N DUP 28
SRR1766448.6909808 chr19 108001 N chr19 108106 N DUP 27
SRR1766445.641220 chr19 108001 N chr19 108106 N DUP 28
SRR1766455.7004062 chr19 108020 N chr19 108277 N DUP 5
SRR1766478.10914553 chr19 108120 N chr19 108206 N DEL 12
SRR1766465.7444298 chr19 108043 N chr19 108100 N DEL 18
SRR1766442.26622570 chr19 108120 N chr19 108206 N DEL 12
SRR1766459.736160 chr19 108152 N chr19 108319 N DEL 5
SRR1766460.5868200 chr19 108152 N chr19 108340 N DEL 7
SRR1766442.24412388 chr19 108120 N chr19 108206 N DEL 12
SRR1766477.11480372 chr19 108093 N chr19 108365 N DUP 6
SRR1766442.18570184 chr19 108076 N chr19 108245 N DUP 17
SRR1766482.10962747 chr19 108014 N chr19 108167 N DUP 19
SRR1766451.2923848 chr19 108014 N chr19 108167 N DUP 19
SRR1766453.3918307 chr19 108014 N chr19 108167 N DUP 19
SRR1766472.9551699 chr19 108100 N chr19 108187 N DUP 5
SRR1766477.9531331 chr19 108014 N chr19 108167 N DUP 24
SRR1766472.8870166 chr19 108014 N chr19 108167 N DUP 29
SRR1766467.1248967 chr19 108093 N chr19 108348 N DUP 7
SRR1766460.1425148 chr19 108093 N chr19 108348 N DUP 8
SRR1766453.3911643 chr19 107913 N chr19 108087 N DEL 11
SRR1766471.6541267 chr19 107972 N chr19 108093 N DEL 4
SRR1766443.9102227 chr19 108091 N chr19 108363 N DUP 5
SRR1766455.7824443 chr19 108091 N chr19 108363 N DUP 6
SRR1766446.7019254 chr19 107972 N chr19 108098 N DEL 1
SRR1766453.10539642 chr19 108118 N chr19 108200 N DUP 10
SRR1766442.34695860 chr19 108025 N chr19 108239 N DUP 5
SRR1766442.25468777 chr19 108153 N chr19 108273 N DUP 5
SRR1766466.8700754 chr19 108153 N chr19 108273 N DUP 5
SRR1766482.9261177 chr19 107966 N chr19 108156 N DEL 5
SRR1766471.5895040 chr19 108036 N chr19 108271 N DEL 2
SRR1766460.6211909 chrX 129154199 N chrX 129154250 N DUP 5
SRR1766451.6734027 chrX 129154206 N chrX 129154347 N DUP 2
SRR1766468.5320785 chrX 129154206 N chrX 129154347 N DUP 5
SRR1766471.12078432 chrX 129154206 N chrX 129154347 N DUP 5
SRR1766442.38665176 chrX 129154206 N chrX 129154347 N DUP 7
SRR1766458.4708992 chrX 129154206 N chrX 129154347 N DUP 7
SRR1766448.260965 chr1 47122119 N chr1 47122175 N DUP 5
SRR1766444.948662 chr8 93734279 N chr8 93734350 N DUP 5
SRR1766447.9573370 chr12 98846114 N chr12 98846173 N DUP 2
SRR1766482.8767373 chr6 38103525 N chr6 38103618 N DUP 2
SRR1766442.40732873 chr6 38103525 N chr6 38103618 N DUP 3
SRR1766469.9347513 chr6 38103525 N chr6 38103618 N DUP 5
SRR1766449.10487788 chr6 38103619 N chr6 38103674 N DEL 13
SRR1766474.6505441 chr6 38103619 N chr6 38103674 N DEL 13
SRR1766476.3675767 chr6 38103619 N chr6 38103674 N DEL 57
SRR1766484.7238743 chr6 38103619 N chr6 38103674 N DEL 43
SRR1766449.2476763 chr6 38103619 N chr6 38103674 N DEL 43
SRR1766460.1082899 chr6 38103619 N chr6 38103674 N DEL 37
SRR1766443.5964584 chr6 38103553 N chr6 38103614 N DEL 6
SRR1766483.1665888 chr6 38103619 N chr6 38103674 N DEL 33
SRR1766448.7012654 chr6 38103619 N chr6 38103674 N DEL 32
SRR1766474.7268480 chr6 38103619 N chr6 38103674 N DEL 30
SRR1766442.11322981 chr6 38103619 N chr6 38103674 N DEL 30
SRR1766459.2346732 chr6 38103619 N chr6 38103674 N DEL 46
SRR1766473.1415475 chr6 38103619 N chr6 38103674 N DEL 14
SRR1766443.5246386 chr6 38103602 N chr6 38103685 N DEL 4
SRR1766450.3860702 chr6 38103597 N chr6 38103680 N DEL 9
SRR1766456.1045756 chr6 38103604 N chr6 38103687 N DEL 2
SRR1766486.1205355 chr7 47736300 N chr7 47736411 N DEL 4
SRR1766444.4120140 chr7 47736367 N chr7 47736539 N DUP 15
SRR1766483.8237834 chr7 47736313 N chr7 47736368 N DEL 4
SRR1766442.27609945 chrX 30602966 N chrX 30603145 N DEL 1
SRR1766456.5270421 chrX 30602965 N chrX 30603015 N DUP 5
SRR1766469.1576879 chrX 30602965 N chrX 30603015 N DUP 5
SRR1766451.10133926 chrX 30603027 N chrX 30603510 N DEL 5
SRR1766448.4797181 chrX 30602902 N chrX 30603030 N DUP 5
SRR1766442.10596542 chrX 30603032 N chrX 30603261 N DEL 5
SRR1766465.3833772 chrX 30602948 N chrX 30603076 N DUP 1
SRR1766442.27358825 chrX 30602948 N chrX 30603076 N DUP 2
SRR1766472.11698995 chrX 30602906 N chrX 30603036 N DEL 5
SRR1766473.8540541 chrX 30602965 N chrX 30603420 N DUP 10
SRR1766485.6897542 chrX 30602996 N chrX 30603126 N DEL 5
SRR1766477.9796129 chrX 30602859 N chrX 30603115 N DEL 5
SRR1766476.1349411 chrX 30602860 N chrX 30603116 N DEL 5
SRR1766448.8688647 chrX 30603179 N chrX 30603404 N DUP 12
SRR1766446.7503658 chrX 30602837 N chrX 30603192 N DEL 1
SRR1766454.2787157 chrX 30602887 N chrX 30603243 N DUP 5
SRR1766456.1890393 chrX 30602889 N chrX 30603245 N DUP 10
SRR1766474.1160062 chrX 30603176 N chrX 30603228 N DEL 6
SRR1766486.2945426 chrX 30603022 N chrX 30603251 N DEL 5
SRR1766456.5270421 chrX 30603022 N chrX 30603251 N DEL 5
SRR1766464.5717867 chrX 30603145 N chrX 30603323 N DUP 7
SRR1766456.660630 chrX 30603145 N chrX 30603323 N DUP 7
SRR1766452.6303539 chrX 30603145 N chrX 30603323 N DUP 7
SRR1766474.7201539 chrX 30603003 N chrX 30603360 N DEL 7
SRR1766453.559428 chrX 30602824 N chrX 30603405 N DUP 5
SRR1766462.7762510 chrX 30602984 N chrX 30603391 N DEL 11
SRR1766464.4629912 chrX 30602906 N chrX 30603391 N DEL 7
SRR1766455.1373640 chr18 62384542 N chr18 62384643 N DUP 1
SRR1766478.7693658 chr1 247091704 N chr1 247091881 N DUP 6
SRR1766461.3889564 chr9 90997439 N chr9 90997496 N DUP 6
SRR1766463.6667281 chr9 90997437 N chr9 90997496 N DUP 8
SRR1766474.6239594 chr9 90997449 N chr9 90997516 N DEL 7
SRR1766473.7923431 chr9 90997450 N chr9 90997521 N DEL 2
SRR1766478.2781509 chr9 90997450 N chr9 90997519 N DEL 4
SRR1766443.6484668 chr6 25206628 N chr6 25206711 N DEL 4
SRR1766476.3014034 chr6 25206628 N chr6 25206711 N DEL 7
SRR1766455.3486668 chr6 25206656 N chr6 25206733 N DUP 24
SRR1766451.858048 chr6 25206655 N chr6 25206732 N DUP 13
SRR1766466.4973155 chr6 25206655 N chr6 25206732 N DUP 15
SRR1766451.4105653 chr6 25206681 N chr6 25206731 N DUP 27
SRR1766469.1862069 chr6 25206656 N chr6 25206733 N DUP 24
SRR1766476.4947481 chr6 25206644 N chr6 25206699 N DUP 13
SRR1766470.8296467 chr6 25206583 N chr6 25206773 N DUP 5
SRR1766465.9915501 chr6 25206713 N chr6 25206784 N DUP 27
SRR1766457.2866596 chr6 25206713 N chr6 25206784 N DUP 25
SRR1766442.47090403 chr6 25206702 N chr6 25206775 N DUP 17
SRR1766485.823053 chr6 25206728 N chr6 25206799 N DUP 8
SRR1766466.9439057 chr6 25206727 N chr6 25206798 N DUP 9
SRR1766447.8831279 chr6 25206659 N chr6 25206737 N DEL 11
SRR1766465.4195719 chr6 25206657 N chr6 25206767 N DEL 16
SRR1766483.11930667 chr6 25206657 N chr6 25206767 N DEL 16
SRR1766470.241301 chr14 76609856 N chr14 76609920 N DEL 5
SRR1766449.6003900 chrX 114387073 N chrX 114387670 N DEL 5
SRR1766442.46609057 chrX 114387100 N chrX 114387232 N DEL 11
SRR1766462.3490905 chrX 114387100 N chrX 114387232 N DEL 11
SRR1766473.11346133 chrX 114387100 N chrX 114387232 N DEL 13
SRR1766442.31322311 chrX 114387100 N chrX 114387232 N DEL 18
SRR1766467.11197680 chrX 114387100 N chrX 114387232 N DEL 19
SRR1766481.10066704 chrX 114387100 N chrX 114387232 N DEL 12
SRR1766471.10706270 chrX 114387100 N chrX 114387232 N DEL 19
SRR1766461.6166102 chrX 114387045 N chrX 114387676 N DUP 23
SRR1766482.10018456 chrX 114387045 N chrX 114387176 N DUP 10
SRR1766449.5694974 chrX 114387043 N chrX 114387387 N DUP 9
SRR1766462.10247388 chrX 114387129 N chrX 114387595 N DEL 11
SRR1766442.45939718 chrX 114387042 N chrX 114387195 N DUP 11
SRR1766450.6626251 chrX 114387120 N chrX 114387406 N DEL 20
SRR1766455.3927219 chrX 114387148 N chrX 114387240 N DEL 20
SRR1766442.43858060 chrX 114387075 N chrX 114387475 N DEL 10
SRR1766479.2283950 chrX 114387120 N chrX 114387406 N DEL 19
SRR1766467.4995991 chrX 114387054 N chrX 114387158 N DUP 6
SRR1766485.943342 chrX 114387063 N chrX 114387387 N DUP 18
SRR1766470.1011863 chrX 114387178 N chrX 114387241 N DEL 11
SRR1766482.8774494 chrX 114387178 N chrX 114387241 N DEL 11
SRR1766462.1869508 chrX 114387159 N chrX 114387401 N DUP 9
SRR1766445.2706233 chrX 114387199 N chrX 114387641 N DUP 28
SRR1766453.9217813 chrX 114387182 N chrX 114387266 N DUP 17
SRR1766454.9028196 chrX 114387199 N chrX 114387641 N DUP 26
SRR1766446.1980675 chrX 114387240 N chrX 114387339 N DEL 1
SRR1766472.8561265 chrX 114387190 N chrX 114387394 N DUP 2
SRR1766445.9650319 chrX 114387221 N chrX 114387385 N DUP 20
SRR1766462.3490905 chrX 114387198 N chrX 114387299 N DEL 14
SRR1766460.6309865 chrX 114387244 N chrX 114387566 N DUP 18
SRR1766472.10854182 chrX 114387221 N chrX 114387385 N DUP 19
SRR1766454.2139521 chrX 114387265 N chrX 114387320 N DUP 12
SRR1766442.5682528 chrX 114387261 N chrX 114387336 N DUP 19
SRR1766467.864445 chrX 114387281 N chrX 114387336 N DUP 8
SRR1766482.8353578 chrX 114387085 N chrX 114387237 N DEL 6
SRR1766481.6934418 chrX 114387221 N chrX 114387385 N DUP 8
SRR1766481.9076653 chrX 114387221 N chrX 114387385 N DUP 13
SRR1766446.5267646 chrX 114387114 N chrX 114387293 N DEL 8
SRR1766442.44913756 chrX 114387315 N chrX 114387541 N DEL 17
SRR1766479.6862988 chrX 114387308 N chrX 114387474 N DUP 21
SRR1766447.1511369 chrX 114387258 N chrX 114387323 N DEL 13
SRR1766472.8561265 chrX 114387175 N chrX 114387342 N DEL 14
SRR1766446.7168921 chrX 114387045 N chrX 114387356 N DUP 1
SRR1766462.10247388 chrX 114387053 N chrX 114387357 N DUP 14
SRR1766443.7709385 chrX 114387321 N chrX 114387505 N DEL 17
SRR1766484.8442413 chrX 114387043 N chrX 114387365 N DUP 6
SRR1766485.2651990 chrX 114387199 N chrX 114387385 N DUP 9
SRR1766465.4836281 chrX 114387199 N chrX 114387385 N DUP 9
SRR1766443.992595 chrX 114387199 N chrX 114387385 N DUP 12
SRR1766442.12813109 chrX 114387199 N chrX 114387385 N DUP 13
SRR1766461.10309545 chrX 114387324 N chrX 114387503 N DEL 12
SRR1766486.1008721 chrX 114387199 N chrX 114387385 N DUP 13
SRR1766442.22025397 chrX 114387063 N chrX 114387366 N DUP 10
SRR1766460.4809186 chrX 114387199 N chrX 114387385 N DUP 13
SRR1766454.5525715 chrX 114387199 N chrX 114387385 N DUP 16
SRR1766465.10827398 chrX 114387199 N chrX 114387385 N DUP 17
SRR1766453.5861128 chrX 114387059 N chrX 114387183 N DUP 20
SRR1766467.864445 chrX 114387178 N chrX 114387299 N DEL 11
SRR1766476.5818927 chrX 114387219 N chrX 114387271 N DEL 5
SRR1766447.986226 chrX 114387221 N chrX 114387385 N DUP 20
SRR1766481.5985479 chrX 114387221 N chrX 114387385 N DUP 21
SRR1766477.10961291 chrX 114387199 N chrX 114387641 N DUP 23
SRR1766477.8918353 chrX 114387080 N chrX 114387323 N DEL 16
SRR1766454.6029977 chrX 114387324 N chrX 114387376 N DEL 8
SRR1766459.6544722 chrX 114387281 N chrX 114387376 N DUP 16
SRR1766484.2316801 chrX 114387190 N chrX 114387280 N DUP 7
SRR1766455.4469180 chrX 114387089 N chrX 114387297 N DEL 11
SRR1766474.5712184 chrX 114387252 N chrX 114387405 N DUP 6
SRR1766473.7390007 chrX 114387258 N chrX 114387341 N DEL 15
SRR1766486.1274959 chrX 114387247 N chrX 114387403 N DUP 17
SRR1766473.9805277 chrX 114387339 N chrX 114387392 N DUP 10
SRR1766443.10125434 chrX 114387120 N chrX 114387406 N DEL 19
SRR1766450.6363542 chrX 114387221 N chrX 114387385 N DUP 11
SRR1766475.948443 chrX 114387342 N chrX 114387395 N DUP 6
SRR1766479.10999255 chrX 114387065 N chrX 114387503 N DUP 7
SRR1766467.9461684 chrX 114387115 N chrX 114387497 N DUP 11
SRR1766469.1993856 chrX 114387221 N chrX 114387385 N DUP 19
SRR1766480.3075486 chrX 114387378 N chrX 114387533 N DEL 16
SRR1766454.10503428 chrX 114387061 N chrX 114387209 N DEL 7
SRR1766445.8908361 chrX 114387352 N chrX 114387576 N DEL 17
SRR1766467.1549694 chrX 114387386 N chrX 114387585 N DUP 22
SRR1766450.6626251 chrX 114387198 N chrX 114387633 N DEL 9
SRR1766456.3887543 chrX 114387198 N chrX 114387633 N DEL 9
SRR1766474.5059490 chrX 114387198 N chrX 114387633 N DEL 9
SRR1766485.2651990 chrX 114387178 N chrX 114387633 N DEL 9
SRR1766445.4499448 chrX 114387082 N chrX 114387633 N DEL 9
SRR1766444.5557979 chrX 114387084 N chrX 114387635 N DEL 9
SRR1766442.12813109 chrX 114387085 N chrX 114387636 N DEL 9
SRR1766479.11426768 chrX 114387085 N chrX 114387636 N DEL 9
SRR1766450.757285 chrX 114387091 N chrX 114387642 N DEL 6
SRR1766451.5714116 chrX 114387057 N chrX 114387646 N DEL 2
SRR1766467.1848268 chr7 577119 N chr7 577230 N DEL 5
SRR1766475.1670285 chr1 104712550 N chr1 104712611 N DEL 7
SRR1766468.7762353 chr1 104712552 N chr1 104712613 N DEL 7
SRR1766459.2333772 chr1 104712553 N chr1 104712614 N DEL 7
SRR1766445.8250367 chr1 104712556 N chr1 104712617 N DEL 5
SRR1766468.6325797 chr8 140120705 N chr8 140120870 N DEL 41
SRR1766477.11085877 chr8 140120731 N chr8 140120784 N DEL 6
SRR1766482.4114782 chr8 140120705 N chr8 140120870 N DEL 12
SRR1766473.4727613 chr8 140120804 N chr8 140120968 N DUP 5
SRR1766466.3542217 chr8 140120661 N chr8 140120970 N DUP 5
SRR1766479.11341268 chr8 140120878 N chr8 140121004 N DUP 4
SRR1766471.1081450 chr8 140120758 N chr8 140120892 N DEL 9
SRR1766465.4070334 chr8 140120706 N chr8 140121019 N DUP 5
SRR1766465.1469828 chr8 140120718 N chr8 140120964 N DEL 5
SRR1766479.5058398 chr8 140120712 N chr8 140121023 N DEL 5
SRR1766473.7101736 chr8 140120912 N chr8 140121059 N DEL 5
SRR1766461.10779610 chr22 11330017 N chr22 11330201 N DUP 9
SRR1766463.3131326 chr22 11330112 N chr22 11330207 N DUP 9
SRR1766482.11513602 chr22 11330017 N chr22 11330201 N DUP 9
SRR1766477.6411351 chr22 11330112 N chr22 11330207 N DUP 10
SRR1766461.1126524 chr22 11330112 N chr22 11330207 N DUP 10
SRR1766478.978308 chr22 11330112 N chr22 11330207 N DUP 5
SRR1766473.8286729 chr22 11330112 N chr22 11330207 N DUP 5
SRR1766442.44900526 chr22 11330112 N chr22 11330207 N DUP 5
SRR1766474.468699 chr22 11330112 N chr22 11330207 N DUP 5
SRR1766479.9239418 chr22 11330112 N chr22 11330207 N DUP 5
SRR1766469.621422 chr22 11330112 N chr22 11330207 N DUP 5
SRR1766458.1610780 chr22 11330117 N chr22 11330212 N DUP 7
SRR1766446.5957593 chr22 11330115 N chr22 11330210 N DUP 5
SRR1766458.6544205 chr22 11330117 N chr22 11330212 N DUP 5
SRR1766462.5862358 chr22 11330117 N chr22 11330212 N DUP 5
SRR1766469.7285934 chr22 11330117 N chr22 11330212 N DUP 5
SRR1766479.2718368 chr22 11330117 N chr22 11330212 N DUP 5
SRR1766443.221821 chr22 11330126 N chr22 11330221 N DUP 6
SRR1766449.529047 chr22 11330126 N chr22 11330221 N DUP 6
SRR1766477.6270182 chr22 11330126 N chr22 11330221 N DUP 6
SRR1766442.5720809 chr22 11330123 N chr22 11330218 N DUP 9
SRR1766442.10339754 chr22 11330119 N chr22 11330214 N DUP 14
SRR1766442.46585745 chr22 11330120 N chr22 11330215 N DUP 12
SRR1766453.3022385 chr22 11330119 N chr22 11330214 N DUP 14
SRR1766455.2889090 chr22 11330122 N chr22 11330217 N DUP 10
SRR1766465.9343204 chr22 11330119 N chr22 11330214 N DUP 13
SRR1766469.7777432 chr22 11330124 N chr22 11330219 N DUP 8
SRR1766482.8128168 chr22 11330119 N chr22 11330214 N DUP 14
SRR1766451.3757380 chr22 11330118 N chr22 11330213 N DUP 4
SRR1766454.6074728 chr22 11330119 N chr22 11330214 N DUP 14
SRR1766476.2525848 chr22 11330064 N chr22 11330248 N DUP 3
SRR1766458.3000531 chr22 11330158 N chr22 11330253 N DUP 4
SRR1766457.3807398 chr22 11330112 N chr22 11330255 N DUP 3
SRR1766473.3213478 chr22 11330158 N chr22 11330253 N DUP 5
SRR1766485.2375891 chr22 11330158 N chr22 11330253 N DUP 5
SRR1766453.2258056 chr22 11330158 N chr22 11330253 N DUP 6
SRR1766449.9862107 chr22 11330158 N chr22 11330253 N DUP 7
SRR1766484.4122207 chr22 11330158 N chr22 11330253 N DUP 7
SRR1766471.9921091 chr22 11330074 N chr22 11330258 N DUP 14
SRR1766466.9241412 chr22 11329930 N chr22 11330265 N DUP 1
SRR1766442.37699834 chr22 11329930 N chr22 11330265 N DUP 5
SRR1766443.8824166 chr22 11329930 N chr22 11330265 N DUP 5
SRR1766462.6168466 chr22 11329930 N chr22 11330265 N DUP 5
SRR1766445.724582 chr22 11329930 N chr22 11330265 N DUP 1
SRR1766442.28315841 chr22 11329930 N chr22 11330265 N DUP 5
SRR1766480.3338276 chr22 11330085 N chr22 11330223 N DEL 5
SRR1766446.1583450 chr22 11330127 N chr22 11330224 N DEL 10
SRR1766448.6459079 chr22 11330045 N chr22 11330231 N DEL 5
SRR1766464.3060280 chr22 11330046 N chr22 11330232 N DEL 5
SRR1766442.4227131 chr12 6884811 N chr12 6884861 N DUP 5
SRR1766442.20095216 chr12 6884811 N chr12 6884861 N DUP 5
SRR1766447.9504807 chr12 6884811 N chr12 6884861 N DUP 5
SRR1766442.36429439 chr12 6884831 N chr12 6884883 N DEL 5
SRR1766442.28306341 chr16 36201564 N chr16 36201929 N DEL 5
SRR1766448.9999981 chr16 36201610 N chr16 36201875 N DUP 5
SRR1766469.7515687 chr2 2536967 N chr2 2537150 N DUP 5
SRR1766459.1808856 chr2 2536967 N chr2 2537150 N DUP 5
SRR1766484.9834079 chr2 2536967 N chr2 2537150 N DUP 5
SRR1766460.523256 chr6 139308114 N chr6 139308165 N DEL 3
SRR1766471.9230917 chr6 139308121 N chr6 139308172 N DEL 5
SRR1766477.9859847 chr6 139308115 N chr6 139308166 N DEL 11
SRR1766478.979686 chr6 139308121 N chr6 139308173 N DEL 14
SRR1766462.3627008 chr6 139308114 N chr6 139308165 N DEL 19
SRR1766444.7308254 chr6 139308124 N chr6 139308175 N DEL 5
SRR1766472.10395538 chr10 132124664 N chr10 132124803 N DUP 5
SRR1766473.10807103 chr4 127417316 N chr4 127417375 N DEL 12
SRR1766476.9377565 chr4 127417316 N chr4 127417375 N DEL 10
SRR1766463.4556652 chr4 127417349 N chr4 127417400 N DUP 9
SRR1766464.4648920 chr4 127417350 N chr4 127417451 N DUP 17
SRR1766471.11284481 chr4 127417364 N chr4 127417415 N DEL 1
SRR1766447.6353005 chr10 33028397 N chr10 33028456 N DEL 12
SRR1766452.1366004 chr10 33028397 N chr10 33028456 N DEL 12
SRR1766465.6949820 chr10 33028393 N chr10 33028456 N DEL 12
SRR1766484.47055 chr10 33028389 N chr10 33028456 N DEL 9
SRR1766448.2835657 chr10 33028347 N chr10 33028455 N DEL 12
SRR1766449.7536950 chr10 33028345 N chr10 33028465 N DEL 6
SRR1766473.2061138 chr10 33028345 N chr10 33028465 N DEL 6
SRR1766484.2727896 chr10 33028346 N chr10 33028466 N DEL 5
SRR1766461.8582858 chr2 871439 N chr2 871549 N DUP 10
SRR1766465.8217467 chr2 871273 N chr2 871439 N DEL 5
SRR1766466.10359749 chr11 98763181 N chr11 98763341 N DUP 5
SRR1766476.10193702 chr11 98763181 N chr11 98763341 N DUP 5
SRR1766482.2649817 chr11 98763181 N chr11 98763341 N DUP 5
SRR1766471.10125929 chr11 98763181 N chr11 98763341 N DUP 5
SRR1766470.6382796 chr11 98763181 N chr11 98763341 N DUP 5
SRR1766450.4025174 chr11 98763181 N chr11 98763341 N DUP 5
SRR1766454.6832720 chr11 98763181 N chr11 98763341 N DUP 5
SRR1766469.6377863 chr7 104824854 N chr7 104824921 N DEL 6
SRR1766474.3588684 chr7 104824856 N chr7 104824923 N DEL 4
SRR1766454.1405065 chr7 31239682 N chr7 31239792 N DEL 8
SRR1766482.4358026 chr7 31239683 N chr7 31239793 N DEL 7
SRR1766455.1058291 chr6 14301674 N chr6 14301845 N DEL 5
SRR1766461.8757488 chr6 14301674 N chr6 14301845 N DEL 5
SRR1766455.9603798 chr6 14301690 N chr6 14301859 N DUP 5
SRR1766452.1494075 chr6 14301698 N chr6 14301867 N DUP 1
SRR1766470.8710263 chr6 14301732 N chr6 14301815 N DUP 5
SRR1766467.1203306 chr6 14301732 N chr6 14301815 N DUP 5
SRR1766476.9592062 chr6 14301732 N chr6 14301815 N DUP 5
SRR1766481.12218179 chr6 14301699 N chr6 14301828 N DEL 5
SRR1766473.970430 chr6 14301753 N chr6 14301838 N DEL 3
SRR1766472.6523051 chr13 19779565 N chr13 19779743 N DEL 10
SRR1766477.8344625 chr13 19779565 N chr13 19779743 N DEL 14
SRR1766471.1368981 chr13 19779635 N chr13 19779813 N DEL 3
SRR1766473.6852899 chr13 19779565 N chr13 19779743 N DEL 5
SRR1766482.1896685 chr13 19779635 N chr13 19779813 N DEL 5
SRR1766477.9576089 chr13 19779546 N chr13 19779673 N DUP 2
SRR1766476.1728858 chr13 19779673 N chr13 19779849 N DUP 5
SRR1766449.4358827 chr13 19779573 N chr13 19779827 N DUP 5
SRR1766473.6483208 chr13 19779546 N chr13 19779673 N DUP 2
SRR1766471.9752054 chr13 19779573 N chr13 19779827 N DUP 5
SRR1766477.1013284 chr13 19779518 N chr13 19779694 N DUP 3
SRR1766443.219929 chr13 19779673 N chr13 19779801 N DEL 10
SRR1766479.349534 chr13 19779673 N chr13 19779801 N DEL 10
SRR1766450.10350474 chr13 19779518 N chr13 19779694 N DUP 5
SRR1766479.2563372 chr13 19779654 N chr13 19779830 N DUP 5
SRR1766447.1361611 chr13 19779636 N chr13 19779734 N DUP 5
SRR1766486.10323399 chr13 19779560 N chr13 19779639 N DEL 5
SRR1766466.9703606 chr13 19779511 N chr13 19779687 N DUP 5
SRR1766449.6485307 chr13 19779511 N chr13 19779687 N DUP 5
SRR1766479.1947079 chr13 19779526 N chr13 19779704 N DEL 5
SRR1766473.6766822 chr13 19779565 N chr13 19779743 N DEL 12
SRR1766472.1382520 chr13 19779528 N chr13 19779706 N DEL 4
SRR1766460.926437 chr13 19779527 N chr13 19779705 N DEL 5
SRR1766485.6256624 chr13 19779528 N chr13 19779832 N DUP 7
SRR1766461.1353669 chr13 19779528 N chr13 19779832 N DUP 7
SRR1766450.7025100 chr13 19779511 N chr13 19779814 N DUP 2
SRR1766445.10374462 chr13 19779623 N chr13 19779848 N DUP 1
SRR1766462.969711 chr13 19779623 N chr13 19779848 N DUP 3
SRR1766479.4372203 chr13 19779511 N chr13 19779814 N DUP 3
SRR1766470.10349113 chr13 19779513 N chr13 19779865 N DUP 8
SRR1766480.3078961 chr8 138865587 N chr8 138865655 N DEL 9
SRR1766470.5637666 chr8 138865753 N chr8 138865864 N DEL 13
SRR1766454.6765661 chr8 138865768 N chr8 138865861 N DEL 10
SRR1766449.5068727 chr8 138865768 N chr8 138865943 N DEL 5
SRR1766478.1055589 chr8 138865740 N chr8 138865981 N DUP 6
SRR1766460.580617 chr8 138865872 N chr8 138865943 N DEL 7
SRR1766484.11026751 chr8 138865526 N chr8 138865762 N DEL 1
SRR1766481.1747106 chr8 138865547 N chr8 138865783 N DEL 5
SRR1766455.7834136 chr8 138865815 N chr8 138865984 N DUP 4
SRR1766472.11657813 chr8 138865828 N chr8 138865997 N DUP 7
SRR1766471.11954221 chr19 38364452 N chr19 38364567 N DUP 5
SRR1766448.170518 chr19 38364461 N chr19 38364654 N DEL 5
SRR1766452.4230313 chr12 132621012 N chr12 132621074 N DEL 2
SRR1766444.6803640 chr12 132621012 N chr12 132621074 N DEL 3
SRR1766486.11242618 chr12 132621012 N chr12 132621074 N DEL 10
SRR1766483.9079138 chr12 132621012 N chr12 132621074 N DEL 10
SRR1766444.871769 chr12 132621012 N chr12 132621074 N DEL 12
SRR1766472.7326404 chr12 132621012 N chr12 132621074 N DEL 6
SRR1766454.1314268 chr12 132621012 N chr12 132621074 N DEL 15
SRR1766447.11354775 chr12 132621012 N chr12 132621074 N DEL 24
SRR1766475.3235225 chr12 132621019 N chr12 132621081 N DEL 8
SRR1766479.1001112 chr12 132621024 N chr12 132621086 N DEL 3
SRR1766447.7367544 chr17 46243538 N chr17 46243633 N DEL 6
SRR1766473.6486702 chr17 46243542 N chr17 46243637 N DEL 2
SRR1766442.22978505 chr17 46243541 N chr17 46243636 N DEL 3
SRR1766442.41022465 chr17 46243541 N chr17 46243636 N DEL 3
SRR1766469.3929845 chr2 34043164 N chr2 34043476 N DEL 5
SRR1766446.6288199 chr2 34043164 N chr2 34043476 N DEL 5
SRR1766442.29395350 chr4 186694162 N chr4 186694229 N DUP 5
SRR1766471.5452198 chr4 186694141 N chr4 186694352 N DEL 1
SRR1766442.15115322 chr4 186694106 N chr4 186694385 N DEL 1
SRR1766483.3965841 chr6 69169652 N chr6 69169738 N DUP 5
SRR1766482.11550261 chr12 8625910 N chr12 8626086 N DUP 5
SRR1766464.8487326 chr12 8625910 N chr12 8626086 N DUP 5
SRR1766479.11222357 chr12 8625907 N chr12 8626132 N DUP 1
SRR1766483.10422334 chr12 8625911 N chr12 8626087 N DUP 5
SRR1766480.1154299 chr12 8625917 N chr12 8626142 N DUP 5
SRR1766454.7610910 chr12 8625928 N chr12 8626104 N DUP 9
SRR1766442.38615234 chr12 8625898 N chr12 8625949 N DEL 5
SRR1766471.411121 chr12 8626054 N chr12 8626105 N DEL 4
SRR1766475.8020788 chr12 8625968 N chr12 8626095 N DUP 3
SRR1766454.5758797 chr12 8625973 N chr12 8626149 N DUP 5
SRR1766442.1168332 chr12 8625912 N chr12 8626088 N DUP 5
SRR1766442.44968965 chr12 8625893 N chr12 8626118 N DUP 3
SRR1766459.11443440 chr12 8625963 N chr12 8626139 N DUP 2
SRR1766451.5136182 chr12 8625891 N chr12 8626070 N DEL 6
SRR1766476.4125421 chr12 8625891 N chr12 8626070 N DEL 6
SRR1766462.10574630 chr12 8625891 N chr12 8626070 N DEL 6
SRR1766442.30666157 chr12 8626070 N chr12 8626167 N DUP 7
SRR1766460.1902711 chr3 9788555 N chr3 9789146 N DEL 4
SRR1766455.9020130 chr3 9788457 N chr3 9789046 N DUP 5
SRR1766456.5769056 chr4 19288874 N chr4 19288965 N DUP 13
SRR1766444.5717475 chr4 19288931 N chr4 19289002 N DEL 9
SRR1766446.7500321 chr4 19288891 N chr4 19289002 N DEL 7
SRR1766442.35802503 chr4 19288895 N chr4 19289002 N DEL 9
SRR1766450.6952426 chr4 19288921 N chr4 19288998 N DEL 2
SRR1766472.5962005 chr4 19288891 N chr4 19289002 N DEL 7
SRR1766479.11150483 chr5 69515425 N chr5 69515551 N DUP 4
SRR1766454.3757606 chr5 69515400 N chr5 69515704 N DUP 5
SRR1766456.5248101 chr5 69515651 N chr5 69515701 N DUP 2
SRR1766452.3654544 chr5 69515568 N chr5 69515745 N DUP 5
SRR1766484.2753568 chr5 69515435 N chr5 69515738 N DUP 6
SRR1766444.2952751 chr5 69515568 N chr5 69515745 N DUP 5
SRR1766472.10154566 chr5 69515568 N chr5 69515745 N DUP 5
SRR1766442.10979661 chr5 69515568 N chr5 69515745 N DUP 12
SRR1766452.6884391 chr5 69515690 N chr5 69515739 N DUP 12
SRR1766477.7031888 chr5 69515689 N chr5 69515738 N DUP 15
SRR1766483.3791478 chr5 69515651 N chr5 69515750 N DUP 1
SRR1766450.5431747 chr5 69515678 N chr5 69515776 N DUP 7
SRR1766476.9013852 chr5 69515690 N chr5 69515788 N DUP 7
SRR1766445.351829 chr5 69515688 N chr5 69515789 N DUP 5
SRR1766463.5740455 chr5 69515678 N chr5 69515776 N DUP 16
SRR1766469.5327789 chr5 69515432 N chr5 69515688 N DEL 6
SRR1766459.4676687 chr5 69515438 N chr5 69515694 N DEL 5
SRR1766463.9509113 chr5 69515433 N chr5 69515689 N DEL 6
SRR1766458.3055678 chr19 14540166 N chr19 14540347 N DEL 5
SRR1766467.6679875 chr16 10702735 N chr16 10703253 N DUP 8
SRR1766485.253810 chr3 127154896 N chr3 127155032 N DUP 1
SRR1766469.4001365 chr3 127155141 N chr3 127155605 N DEL 3
SRR1766452.3597420 chr3 127155024 N chr3 127155190 N DUP 9
SRR1766442.18103555 chr3 127155045 N chr3 127155621 N DUP 1
SRR1766481.9682978 chr3 127155110 N chr3 127155184 N DUP 5
SRR1766479.6358088 chr3 127155110 N chr3 127155184 N DUP 7
SRR1766478.6919107 chr3 127155114 N chr3 127155216 N DUP 2
SRR1766442.21952003 chr3 127155225 N chr3 127155469 N DEL 12
SRR1766483.9189142 chr3 127155271 N chr3 127155601 N DEL 4
SRR1766485.3178873 chr3 127155131 N chr3 127155197 N DEL 9
SRR1766446.3799978 chr3 127155125 N chr3 127155199 N DEL 9
SRR1766451.3826749 chr3 127155096 N chr3 127155202 N DEL 6
SRR1766453.9507247 chr3 127155096 N chr3 127155202 N DEL 6
SRR1766486.2971203 chr3 127155436 N chr3 127155675 N DEL 9
SRR1766481.9682978 chr3 127155101 N chr3 127155465 N DUP 4
SRR1766485.10270276 chr3 127155101 N chr3 127155465 N DUP 4
SRR1766442.28404641 chr3 127155465 N chr3 127155702 N DEL 4
SRR1766472.6537879 chr3 127155465 N chr3 127155702 N DEL 4
SRR1766462.3972456 chr3 127155083 N chr3 127155517 N DUP 1
SRR1766485.7810432 chr3 127155310 N chr3 127155555 N DUP 12
SRR1766478.8704995 chr3 127155173 N chr3 127155508 N DEL 5
SRR1766448.7619888 chr3 127155099 N chr3 127155619 N DUP 8
SRR1766469.7798101 chr3 127155515 N chr3 127155660 N DUP 2
SRR1766446.5380723 chr3 127155036 N chr3 127155666 N DUP 5
SRR1766472.1748152 chr3 127155570 N chr3 127155715 N DUP 4
SRR1766482.817656 chr3 127155242 N chr3 127155598 N DEL 8
SRR1766476.6708643 chr3 127155026 N chr3 127155708 N DUP 4
SRR1766480.981493 chr3 127155047 N chr3 127155597 N DEL 11
SRR1766467.8649616 chr3 127155255 N chr3 127155601 N DEL 10
SRR1766455.1926442 chr3 127155489 N chr3 127155608 N DEL 8
SRR1766442.29960524 chr3 127155102 N chr3 127155688 N DEL 2
SRR1766471.6741755 chr3 127155048 N chr3 127155690 N DEL 4
SRR1766481.162558 chr19 480611 N chr19 481106 N DEL 1
SRR1766460.3921967 chr19 480611 N chr19 481056 N DEL 5
SRR1766442.1664899 chr19 480705 N chr19 481149 N DEL 5
SRR1766480.8608351 chr19 480747 N chr19 481594 N DEL 2
SRR1766463.10639667 chr19 480778 N chr19 481549 N DEL 18
SRR1766449.9175319 chr19 480733 N chr19 480819 N DUP 6
SRR1766470.8243208 chr19 480653 N chr19 480779 N DUP 4
SRR1766483.4717152 chr19 480830 N chr19 481562 N DEL 6
SRR1766455.3666255 chr19 480665 N chr19 480818 N DEL 5
SRR1766480.8608351 chr19 480704 N chr19 480805 N DEL 3
SRR1766483.4152223 chr19 480691 N chr19 480818 N DEL 14
SRR1766442.25929985 chr19 480906 N chr19 481059 N DEL 23
SRR1766464.10349951 chr19 480960 N chr19 481277 N DEL 5
SRR1766479.5614508 chr19 480604 N chr19 480983 N DUP 5
SRR1766475.3744517 chr19 480929 N chr19 481158 N DEL 10
SRR1766453.5503909 chr19 480898 N chr19 481100 N DUP 5
SRR1766450.4813774 chr19 480793 N chr19 481021 N DUP 9
SRR1766478.473554 chr19 481012 N chr19 481580 N DEL 8
SRR1766472.6534139 chr19 481005 N chr19 481057 N DEL 13
SRR1766479.4817102 chr19 480992 N chr19 481586 N DEL 17
SRR1766442.1664899 chr19 480988 N chr19 481088 N DUP 5
SRR1766442.30394899 chr19 480744 N chr19 480960 N DEL 5
SRR1766476.2176850 chr19 481056 N chr19 481586 N DEL 2
SRR1766443.6832162 chr19 481022 N chr19 481588 N DUP 15
SRR1766458.6012420 chr19 481097 N chr19 481311 N DUP 5
SRR1766445.10021108 chr19 480779 N chr19 481097 N DEL 5
SRR1766466.10721516 chr19 481073 N chr19 481211 N DUP 1
SRR1766442.46906939 chr19 480817 N chr19 481148 N DEL 5
SRR1766466.1868984 chr19 480966 N chr19 481195 N DEL 5
SRR1766473.4954154 chr19 481333 N chr19 481586 N DEL 5
SRR1766483.5298728 chr19 480660 N chr19 481257 N DEL 5
SRR1766459.8474506 chr19 480688 N chr19 481396 N DEL 4
SRR1766468.3313706 chr19 480688 N chr19 481396 N DEL 1
SRR1766459.11321447 chr19 480666 N chr19 481486 N DUP 9
SRR1766471.5598663 chr19 480663 N chr19 481533 N DUP 5
SRR1766464.9260921 chr19 481447 N chr19 481721 N DUP 5
SRR1766476.255577 chr19 481549 N chr19 481638 N DEL 5
SRR1766472.2297656 chr19 481509 N chr19 481610 N DUP 4
SRR1766459.10390478 chr19 480633 N chr19 481480 N DEL 5
SRR1766460.7260932 chr19 480631 N chr19 481516 N DEL 10
SRR1766461.4987839 chr19 480629 N chr19 481514 N DEL 5
SRR1766486.4514432 chr19 481591 N chr19 481665 N DUP 17
SRR1766454.1092975 chr19 480653 N chr19 481649 N DUP 6
SRR1766484.3248593 chr19 480653 N chr19 481649 N DUP 7
SRR1766453.9627248 chr19 480653 N chr19 481649 N DUP 9
SRR1766459.11167873 chr19 480653 N chr19 481649 N DUP 11
SRR1766459.10428478 chr19 480788 N chr19 481623 N DEL 20
SRR1766442.29871329 chr19 481321 N chr19 481648 N DEL 20
SRR1766475.3884818 chr19 481321 N chr19 481648 N DEL 18
SRR1766467.114115 chr19 480777 N chr19 481648 N DEL 7
SRR1766452.1581638 chr19 480631 N chr19 481654 N DEL 4
SRR1766483.9409280 chr19 480633 N chr19 481656 N DEL 7
SRR1766472.4536524 chr19 480678 N chr19 481689 N DEL 5
SRR1766484.10780905 chr19 481725 N chr19 481823 N DEL 10
SRR1766480.1931054 chr11 131680844 N chr11 131680925 N DUP 5
SRR1766457.1057925 chr11 131680982 N chr11 131681073 N DUP 14
SRR1766462.7397654 chr11 131680967 N chr11 131681348 N DUP 5
SRR1766470.6441119 chr11 131680966 N chr11 131681347 N DUP 6
SRR1766442.6059651 chr11 131680973 N chr11 131681746 N DUP 3
SRR1766454.7328645 chr11 131680976 N chr11 131681883 N DUP 4
SRR1766467.6577654 chr11 131680936 N chr11 131681081 N DUP 15
SRR1766476.4492416 chr11 131680937 N chr11 131681142 N DUP 9
SRR1766478.1188501 chr11 131681162 N chr11 131681457 N DEL 5
SRR1766455.7994078 chr11 131680951 N chr11 131681064 N DEL 9
SRR1766444.700229 chr11 131681184 N chr11 131681311 N DEL 14
SRR1766478.3782222 chr11 131681102 N chr11 131681481 N DUP 6
SRR1766451.24679 chr11 131681003 N chr11 131681170 N DUP 4
SRR1766465.1142782 chr11 131681142 N chr11 131681311 N DEL 19
SRR1766462.8258259 chr11 131680938 N chr11 131681267 N DUP 12
SRR1766449.1260167 chr11 131681128 N chr11 131681777 N DEL 7
SRR1766480.8202628 chr11 131681049 N chr11 131681176 N DEL 3
SRR1766454.2824306 chr11 131680952 N chr11 131681185 N DEL 11
SRR1766448.9822195 chr11 131681084 N chr11 131681293 N DUP 3
SRR1766484.5088782 chr11 131680938 N chr11 131681395 N DUP 14
SRR1766470.5143778 chr11 131681014 N chr11 131681395 N DUP 5
SRR1766467.3543878 chr11 131681012 N chr11 131681311 N DEL 5
SRR1766482.5509295 chr11 131681134 N chr11 131681345 N DEL 10
SRR1766447.7790093 chr11 131680952 N chr11 131681319 N DEL 12
SRR1766471.2917280 chr11 131680937 N chr11 131681450 N DUP 13
SRR1766443.11224912 chr11 131680936 N chr11 131681449 N DUP 5
SRR1766471.8583522 chr11 131681006 N chr11 131681347 N DEL 5
SRR1766467.1193630 chr11 131681014 N chr11 131681395 N DUP 8
SRR1766461.4282895 chr11 131681000 N chr11 131681465 N DUP 5
SRR1766477.4888951 chr11 131680998 N chr11 131681463 N DUP 5
SRR1766486.9741504 chr11 131681574 N chr11 131681745 N DEL 11
SRR1766480.4244510 chr11 131681024 N chr11 131681581 N DUP 14
SRR1766486.9812069 chr11 131680938 N chr11 131681523 N DUP 20
SRR1766448.3585115 chr11 131680963 N chr11 131681420 N DEL 5
SRR1766442.22272196 chr11 131680956 N chr11 131681431 N DEL 11
SRR1766472.5422475 chr11 131681127 N chr11 131681464 N DEL 13
SRR1766485.9659235 chr11 131680954 N chr11 131681449 N DEL 13
SRR1766475.10705296 chr11 131681127 N chr11 131681464 N DEL 13
SRR1766452.3067670 chr11 131681127 N chr11 131681464 N DEL 13
SRR1766442.34978219 chr11 131681268 N chr11 131681525 N DEL 5
SRR1766484.10828974 chr11 131681396 N chr11 131681525 N DUP 2
SRR1766468.106180 chr11 131681059 N chr11 131681396 N DEL 5
SRR1766476.7867569 chr11 131681016 N chr11 131681529 N DEL 5
SRR1766442.46337649 chr11 131681389 N chr11 131681646 N DUP 5
SRR1766463.3795159 chr11 131681389 N chr11 131681646 N DUP 5
SRR1766449.1260167 chr11 131681033 N chr11 131681592 N DEL 5
SRR1766451.8219698 chr11 131680952 N chr11 131681617 N DEL 5
SRR1766478.7370959 chr11 131680954 N chr11 131681631 N DEL 1
SRR1766443.7504084 chr11 131681691 N chr11 131681958 N DUP 13
SRR1766464.876466 chr11 131681002 N chr11 131681645 N DEL 5
SRR1766485.9168166 chr11 131681704 N chr11 131681881 N DEL 11
SRR1766482.4839095 chr11 131681398 N chr11 131681743 N DUP 10
SRR1766467.7049026 chr11 131681004 N chr11 131681691 N DEL 5
SRR1766445.2478786 chr11 131681391 N chr11 131681478 N DEL 16
SRR1766449.5389202 chr11 131681034 N chr11 131681763 N DEL 6
SRR1766482.446016 chr11 131681380 N chr11 131681861 N DUP 3
SRR1766480.4230284 chr11 131680951 N chr11 131681746 N DEL 14
SRR1766453.3738605 chr11 131680848 N chr11 131681761 N DEL 3
SRR1766446.106277 chr11 131680971 N chr11 131681836 N DUP 11
SRR1766471.9004494 chr11 131680960 N chr11 131681797 N DEL 20
SRR1766476.10535103 chr11 131681072 N chr11 131681801 N DEL 1
SRR1766461.3533903 chr11 131681398 N chr11 131681877 N DUP 5
SRR1766466.9379062 chr11 131681857 N chr11 131681944 N DUP 5
SRR1766477.5812676 chr11 131681857 N chr11 131681944 N DUP 5
SRR1766451.10582359 chr11 131681038 N chr11 131681859 N DEL 5
SRR1766458.9306513 chr6 29845661 N chr6 29845716 N DUP 1
SRR1766482.6897894 chr6 29845661 N chr6 29845716 N DUP 5
SRR1766476.8407240 chr6 29845613 N chr6 29845724 N DUP 5
SRR1766451.420466 chr6 29845613 N chr6 29845724 N DUP 5
SRR1766486.9776361 chr6 29845613 N chr6 29845724 N DUP 5
SRR1766481.3905344 chr6 29845679 N chr6 29845736 N DEL 5
SRR1766477.3761220 chr6 29845679 N chr6 29845736 N DEL 5
SRR1766452.10168761 chr6 29845679 N chr6 29845736 N DEL 5
SRR1766457.7149944 chr6 29845628 N chr6 29845741 N DEL 5
SRR1766463.7176843 chr6 29845629 N chr6 29845742 N DEL 5
SRR1766462.5304650 chr6 29845631 N chr6 29845744 N DEL 5
SRR1766462.10713797 chr6 29845631 N chr6 29845744 N DEL 5
SRR1766453.3161536 chr9 125780091 N chr9 125780217 N DUP 5
SRR1766486.8277557 chr9 125780243 N chr9 125780420 N DEL 5
SRR1766460.11013096 chr9 125780243 N chr9 125780420 N DEL 10
SRR1766457.6876832 chr9 125780243 N chr9 125780420 N DEL 15
SRR1766463.1836404 chr9 125780243 N chr9 125780420 N DEL 15
SRR1766469.3729991 chr9 125780032 N chr9 125780208 N DEL 5
SRR1766457.3100563 chr9 125780032 N chr9 125780208 N DEL 5
SRR1766473.1715817 chr9 125780032 N chr9 125780208 N DEL 5
SRR1766475.3195745 chr9 125780032 N chr9 125780208 N DEL 5
SRR1766448.1070765 chr9 125780065 N chr9 125780192 N DEL 3
SRR1766474.1213355 chr9 125780032 N chr9 125780208 N DEL 5
SRR1766466.8953459 chr9 125779983 N chr9 125780284 N DUP 15
SRR1766448.2256244 chr9 125779983 N chr9 125780284 N DUP 5
SRR1766442.17904595 chr9 125780243 N chr9 125780420 N DEL 3
SRR1766465.1996166 chr9 125780037 N chr9 125780340 N DEL 5
SRR1766457.4803259 chr5 558862 N chr5 559301 N DEL 1
SRR1766478.5310482 chr5 558862 N chr5 559301 N DEL 1
SRR1766442.3598853 chr5 558893 N chr5 559259 N DEL 4
SRR1766449.2096247 chr5 558910 N chr5 559130 N DEL 4
SRR1766449.2258755 chr5 558891 N chr5 559257 N DEL 5
SRR1766467.1351607 chr5 558891 N chr5 559257 N DEL 5
SRR1766461.1385920 chr5 558894 N chr5 559260 N DEL 2
SRR1766453.1613995 chr5 558831 N chr5 558903 N DUP 5
SRR1766448.4552331 chr5 558906 N chr5 559126 N DEL 5
SRR1766442.20597419 chr5 558961 N chr5 559254 N DEL 5
SRR1766475.5831005 chr5 558888 N chr5 559325 N DUP 5
SRR1766448.8373151 chr5 558979 N chr5 559126 N DEL 5
SRR1766484.12051404 chr5 558934 N chr5 559227 N DEL 5
SRR1766471.11038675 chr5 559049 N chr5 559269 N DEL 4
SRR1766447.5200106 chr5 559049 N chr5 559269 N DEL 5
SRR1766483.2122065 chr5 559049 N chr5 559269 N DEL 5
SRR1766471.1531709 chr5 558891 N chr5 559038 N DEL 5
SRR1766455.6755346 chr5 558891 N chr5 559038 N DEL 5
SRR1766442.8085411 chr5 558896 N chr5 559043 N DEL 5
SRR1766469.3798052 chr5 558940 N chr5 559233 N DEL 8
SRR1766465.2719337 chr5 558931 N chr5 559224 N DEL 5
SRR1766467.2516924 chr5 559157 N chr5 559231 N DEL 5
SRR1766445.9089361 chr5 559166 N chr5 559240 N DEL 2
SRR1766457.1090462 chr5 559162 N chr5 559236 N DEL 3
SRR1766449.2258755 chr5 558868 N chr5 559307 N DEL 5
SRR1766442.37200262 chr10 133121586 N chr10 133121732 N DUP 5
SRR1766476.6492879 chr10 133121747 N chr10 133121824 N DEL 5
SRR1766463.3716772 chr10 133121487 N chr10 133121775 N DUP 10
SRR1766479.9604286 chr10 133121682 N chr10 133121852 N DUP 5
SRR1766456.3853258 chr10 133121598 N chr10 133121805 N DEL 5
SRR1766455.7979304 chr7 100741765 N chr7 100742068 N DEL 5
SRR1766457.2160339 chr7 100741685 N chr7 100742135 N DUP 1
SRR1766471.11537251 chr7 100741645 N chr7 100741746 N DEL 2
SRR1766452.5085712 chr7 100741864 N chr7 100742089 N DEL 5
SRR1766461.8596346 chr7 100741864 N chr7 100741990 N DUP 5
SRR1766442.3770754 chr17 7176759 N chr17 7176886 N DUP 1
SRR1766464.6843283 chr17 7176736 N chr17 7176861 N DEL 7
SRR1766469.776599 chr17 7176740 N chr17 7176865 N DEL 6
SRR1766468.2865332 chr20 62451715 N chr20 62452064 N DEL 5
SRR1766445.10287398 chr20 62451728 N chr20 62452069 N DEL 7
SRR1766466.5977059 chr20 62451900 N chr20 62452000 N DUP 5
SRR1766462.10970962 chr20 62452080 N chr20 62452262 N DUP 10
SRR1766480.7115752 chr20 62452070 N chr20 62452272 N DUP 9
SRR1766484.6447295 chr20 62451883 N chr20 62452319 N DEL 5
SRR1766460.6861771 chr20 3785326 N chr20 3785390 N DEL 5
SRR1766465.9045589 chr7 147396163 N chr7 147396342 N DEL 9
SRR1766481.7251598 chr1 143262470 N chr1 143262771 N DUP 5
SRR1766465.9009945 chr1 143262478 N chr1 143262779 N DUP 4
SRR1766478.5899883 chr1 143262461 N chr1 143262762 N DUP 1
SRR1766463.8450677 chr1 143262455 N chr1 143262756 N DUP 6
SRR1766475.2324720 chr1 143262478 N chr1 143262779 N DUP 5
SRR1766446.8272106 chr1 143262459 N chr1 143262737 N DUP 3
SRR1766450.7563119 chr1 143262470 N chr1 143262771 N DUP 5
SRR1766484.3408005 chr1 143262479 N chr1 143262780 N DUP 5
SRR1766455.4215534 chr1 143262458 N chr1 143262759 N DUP 4
SRR1766454.4975628 chr1 143262475 N chr1 143262776 N DUP 5
SRR1766461.9215315 chr1 143262478 N chr1 143262779 N DUP 5
SRR1766448.9957486 chr1 143262456 N chr1 143262507 N DUP 3
SRR1766449.247594 chr1 143262472 N chr1 143262773 N DUP 5
SRR1766454.10619763 chr1 143262478 N chr1 143262779 N DUP 5
SRR1766447.5522415 chr1 143262478 N chr1 143262779 N DUP 3
SRR1766481.2841439 chr1 143262495 N chr1 143262595 N DUP 5
SRR1766456.5366011 chr1 143262480 N chr1 143262781 N DUP 5
SRR1766454.3478782 chr1 143262472 N chr1 143262773 N DUP 3
SRR1766474.11038714 chr1 143262452 N chr1 143262503 N DUP 1
SRR1766479.9285635 chr1 143262470 N chr1 143262570 N DUP 5
SRR1766478.1427738 chr1 143262478 N chr1 143262779 N DUP 5
SRR1766449.4927109 chr1 143262457 N chr1 143262758 N DUP 5
SRR1766471.11866583 chr1 143262467 N chr1 143262696 N DUP 5
SRR1766442.19650328 chr1 143262473 N chr1 143262774 N DUP 2
SRR1766481.8501839 chr1 143262470 N chr1 143262771 N DUP 5
SRR1766454.10619763 chr1 143262471 N chr1 143262772 N DUP 5
SRR1766453.9316181 chr1 143262478 N chr1 143262779 N DUP 5
SRR1766467.8439593 chr20 18022093 N chr20 18022993 N DEL 5
SRR1766448.4643441 chr20 18022093 N chr20 18022993 N DEL 5
SRR1766479.9930182 chr20 18022172 N chr20 18022478 N DEL 3
SRR1766462.8629128 chr20 18022169 N chr20 18022475 N DEL 5
SRR1766470.3524798 chr20 18022148 N chr20 18022512 N DEL 5
SRR1766455.3391460 chr20 18022168 N chr20 18022474 N DEL 5
SRR1766465.652876 chr20 18022168 N chr20 18022474 N DEL 5
SRR1766456.5901476 chr20 18022168 N chr20 18022474 N DEL 5
SRR1766472.10233955 chr20 18022168 N chr20 18022474 N DEL 5
SRR1766445.2606449 chr20 18022168 N chr20 18022474 N DEL 5
SRR1766471.974741 chr20 18022110 N chr20 18022314 N DUP 5
SRR1766442.22632508 chr20 18022114 N chr20 18023012 N DUP 2
SRR1766460.11014805 chr20 18022266 N chr20 18022702 N DEL 10
SRR1766462.1631439 chr20 18022195 N chr20 18022499 N DUP 5
SRR1766442.30880696 chr20 18022267 N chr20 18023122 N DEL 1
SRR1766472.7175497 chr20 18022421 N chr20 18022754 N DEL 5
SRR1766472.8465826 chr20 18022180 N chr20 18022484 N DUP 5
SRR1766467.8439593 chr20 18022222 N chr20 18022396 N DEL 5
SRR1766479.9930182 chr20 18022337 N chr20 18022394 N DEL 10
SRR1766483.1002366 chr20 18022498 N chr20 18022859 N DEL 10
SRR1766470.4745316 chr20 18022411 N chr20 18023429 N DUP 4
SRR1766485.7988599 chr20 18022413 N chr20 18023107 N DUP 2
SRR1766444.7293689 chr20 18022169 N chr20 18022473 N DUP 11
SRR1766461.595106 chr20 18022556 N chr20 18022859 N DEL 5
SRR1766470.306636 chr20 18022239 N chr20 18022587 N DUP 3
SRR1766465.2628934 chr20 18022214 N chr20 18022520 N DEL 4
SRR1766481.6623817 chr20 18022361 N chr20 18022507 N DEL 9
SRR1766445.10054169 chr20 18022252 N chr20 18022515 N DEL 1
SRR1766442.1739994 chr20 18022232 N chr20 18022610 N DEL 19
SRR1766458.8738183 chr20 18022224 N chr20 18022602 N DEL 19
SRR1766475.5806936 chr20 18022233 N chr20 18022611 N DEL 19
SRR1766452.2423012 chr20 18022166 N chr20 18022602 N DEL 17
SRR1766470.4803338 chr20 18022756 N chr20 18023456 N DUP 5
SRR1766464.251462 chr20 18022243 N chr20 18022893 N DUP 5
SRR1766470.7086420 chr20 18022243 N chr20 18022893 N DUP 5
SRR1766484.7050357 chr20 18022243 N chr20 18022893 N DUP 5
SRR1766466.9299810 chr20 18022243 N chr20 18022893 N DUP 5
SRR1766484.7050357 chr20 18022243 N chr20 18022893 N DUP 5
SRR1766442.21459205 chr20 18022243 N chr20 18022893 N DUP 5
SRR1766484.9461607 chr20 18022243 N chr20 18022893 N DUP 5
SRR1766446.3629899 chr20 18022348 N chr20 18022826 N DEL 5
SRR1766443.9866989 chr20 18022352 N chr20 18022830 N DEL 5
SRR1766481.5395403 chr20 18022352 N chr20 18022830 N DEL 5
SRR1766449.3501766 chr20 18022721 N chr20 18022836 N DEL 10
SRR1766473.2436685 chr20 18022230 N chr20 18022896 N DEL 10
SRR1766473.8286337 chr20 18022715 N chr20 18022902 N DEL 5
SRR1766465.8939666 chr20 18022781 N chr20 18022897 N DEL 11
SRR1766473.7278593 chr20 18022234 N chr20 18022900 N DEL 5
SRR1766483.391723 chr20 18022903 N chr20 18022990 N DUP 5
SRR1766461.2824127 chr20 18022258 N chr20 18022910 N DEL 1
SRR1766480.6378122 chr20 18022779 N chr20 18023012 N DEL 9
SRR1766457.4923504 chr20 18022213 N chr20 18023039 N DEL 10
SRR1766464.10273931 chr20 18022721 N chr20 18023068 N DEL 14
SRR1766470.306636 chr20 18022352 N chr20 18023047 N DEL 4
SRR1766482.2098656 chr20 18022708 N chr20 18023055 N DEL 5
SRR1766443.9264102 chr20 18022368 N chr20 18023063 N DEL 3
SRR1766459.434951 chr20 18022865 N chr20 18023069 N DEL 7
SRR1766444.7058870 chr20 18022697 N chr20 18023217 N DUP 1
SRR1766473.10015669 chr20 18023117 N chr20 18023233 N DUP 1
SRR1766442.36073307 chr20 18022305 N chr20 18023175 N DEL 6
SRR1766473.10484335 chr20 18023340 N chr20 18023487 N DEL 13
SRR1766470.1795646 chr20 18022317 N chr20 18023334 N DEL 10
SRR1766468.5036645 chr20 18022288 N chr20 18023408 N DEL 5
SRR1766443.2736729 chr20 18023106 N chr20 18023460 N DEL 20
SRR1766466.3391961 chr6 9162872 N chr6 9163014 N DUP 8
SRR1766443.698099 chr6 9162872 N chr6 9163014 N DUP 9
SRR1766469.1243811 chr6 9162872 N chr6 9163014 N DUP 9
SRR1766485.9082321 chr6 9162886 N chr6 9163027 N DEL 7
SRR1766442.34298947 chr6 9163024 N chr6 9163077 N DUP 10
SRR1766460.11236143 chr11 17764211 N chr11 17764341 N DUP 13
SRR1766442.43461976 chrX 82073193 N chrX 82073260 N DEL 2
SRR1766450.1297426 chrX 82073193 N chrX 82073260 N DEL 2
SRR1766455.3685489 chrX 82073193 N chrX 82073260 N DEL 2
SRR1766442.7312799 chrX 82073193 N chrX 82073260 N DEL 3
SRR1766469.8044231 chrX 82073193 N chrX 82073260 N DEL 8
SRR1766478.10901455 chrX 82073193 N chrX 82073260 N DEL 9
SRR1766468.742747 chrX 82073193 N chrX 82073286 N DEL 12
SRR1766460.1876172 chr19 16379857 N chr19 16380041 N DEL 1
SRR1766442.21135648 chr19 16379857 N chr19 16380300 N DEL 5
SRR1766445.7258264 chr19 16379742 N chr19 16379926 N DUP 5
SRR1766473.1053484 chr19 16379742 N chr19 16379926 N DUP 5
SRR1766453.10092310 chr19 16379956 N chr19 16380251 N DEL 2
SRR1766479.13149448 chr19 16379964 N chr19 16380370 N DEL 10
SRR1766469.8867015 chr19 16379957 N chr19 16380289 N DEL 20
SRR1766459.10379201 chr19 16379938 N chr19 16380157 N DUP 5
SRR1766483.12187897 chr19 16379938 N chr19 16380157 N DUP 5
SRR1766468.1424378 chr19 16379938 N chr19 16380157 N DUP 5
SRR1766443.5770032 chr19 16379759 N chr19 16379945 N DEL 2
SRR1766473.5105499 chr19 16379759 N chr19 16379945 N DEL 2
SRR1766486.1132901 chr19 16380087 N chr19 16380199 N DEL 1
SRR1766444.4134240 chr19 16379926 N chr19 16380036 N DEL 18
SRR1766442.35771538 chr19 16380192 N chr19 16380378 N DEL 5
SRR1766486.10551009 chr19 16380192 N chr19 16380378 N DEL 5
SRR1766455.4096884 chr19 16380209 N chr19 16380393 N DUP 4
SRR1766460.1876172 chr19 16380211 N chr19 16380395 N DUP 2
SRR1766467.1893155 chr19 16380212 N chr19 16380396 N DUP 1
SRR1766442.31304083 chr19 16379738 N chr19 16380255 N DEL 1
SRR1766484.8151235 chr19 16379850 N chr19 16380293 N DEL 25
SRR1766447.1111851 chr19 16379807 N chr19 16380470 N DUP 1
SRR1766450.7206543 chr19 16379741 N chr19 16380369 N DEL 5
SRR1766460.7979433 chr19 16380399 N chr19 16380620 N DUP 10
SRR1766469.8867015 chr19 16379891 N chr19 16380630 N DEL 5
SRR1766455.2311870 chr19 16379891 N chr19 16380630 N DEL 5
SRR1766469.526719 chr19 16379905 N chr19 16380644 N DEL 5
SRR1766461.4552057 chr19 16380511 N chr19 16380697 N DEL 5
SRR1766479.12977883 chr3 134701420 N chr3 134701481 N DEL 7
SRR1766478.6165479 chr3 134701349 N chr3 134701446 N DUP 3
SRR1766443.654935 chr3 134701349 N chr3 134701446 N DUP 8
SRR1766446.5244203 chr3 134701397 N chr3 134701472 N DUP 6
SRR1766465.6388849 chr3 134701374 N chr3 134701449 N DUP 6
SRR1766471.5202884 chr3 134701378 N chr3 134701453 N DUP 3
SRR1766466.6781506 chr3 134701429 N chr3 134701482 N DUP 19
SRR1766458.332714 chr3 134701429 N chr3 134701482 N DUP 22
SRR1766483.5989940 chr3 134701429 N chr3 134701482 N DUP 22
SRR1766473.3623053 chr3 134701427 N chr3 134701504 N DUP 34
SRR1766457.7995779 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766477.7775706 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766459.4379318 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766470.6180568 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766474.10151694 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766471.9587337 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766452.1432668 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766442.41086000 chr3 134701427 N chr3 134701504 N DUP 35
SRR1766445.5422077 chr3 134701427 N chr3 134701504 N DUP 36
SRR1766486.3719446 chr3 134701427 N chr3 134701504 N DUP 41
SRR1766447.5094949 chr3 134701427 N chr3 134701504 N DUP 44
SRR1766449.9176559 chr3 134701384 N chr3 134701441 N DEL 1
SRR1766449.9298248 chr3 134701447 N chr3 134701522 N DUP 8
SRR1766462.793001 chr3 134701368 N chr3 134701427 N DEL 18
SRR1766482.12756642 chr3 134701446 N chr3 134701521 N DUP 14
SRR1766485.5117594 chr3 134701351 N chr3 134701552 N DUP 10
SRR1766448.2380883 chr3 134701351 N chr3 134701552 N DUP 10
SRR1766481.556751 chr12 105392911 N chr12 105392986 N DEL 3
SRR1766460.3131267 chr12 105392911 N chr12 105392986 N DEL 4
SRR1766480.1314780 chr1 4939639 N chr1 4939744 N DEL 1
SRR1766480.2346701 chr1 4939626 N chr1 4939729 N DUP 15
SRR1766481.2051429 chr1 4939626 N chr1 4939729 N DUP 14
SRR1766457.8085612 chr1 4939626 N chr1 4939729 N DUP 13
SRR1766481.8133118 chr20 60500422 N chr20 60500985 N DEL 5
SRR1766485.8511816 chr20 60500445 N chr20 60500870 N DEL 5
SRR1766450.5091368 chr20 60500447 N chr20 60500985 N DEL 5
SRR1766450.4553644 chr20 60500444 N chr20 60501426 N DEL 6
SRR1766453.6249867 chr20 60500457 N chr20 60500807 N DEL 4
SRR1766483.547354 chr20 60500378 N chr20 60500501 N DUP 1
SRR1766466.9328090 chr20 60500434 N chr20 60500551 N DUP 5
SRR1766460.3772926 chr20 60500659 N chr20 60501004 N DEL 5
SRR1766460.878317 chr20 60500735 N chr20 60501080 N DEL 15
SRR1766470.2244504 chr20 60500397 N chr20 60500653 N DEL 5
SRR1766462.2874078 chr20 60500821 N chr20 60501191 N DEL 5
SRR1766449.4284463 chr20 60500906 N chr20 60501395 N DEL 4
SRR1766442.18288483 chr20 60500511 N chr20 60500837 N DEL 5
SRR1766460.8051837 chr20 60500396 N chr20 60500846 N DEL 10
SRR1766451.2555662 chr20 60500410 N chr20 60500902 N DUP 2
SRR1766462.5980356 chr20 60501006 N chr20 60501395 N DEL 4
SRR1766477.10646060 chr20 60500665 N chr20 60501010 N DEL 9
SRR1766483.547354 chr20 60500395 N chr20 60501189 N DEL 10
SRR1766464.6782220 chr20 60501214 N chr20 60501476 N DUP 5
SRR1766457.8805986 chr20 60500814 N chr20 60501370 N DUP 5
SRR1766451.2555662 chr20 60500505 N chr20 60501275 N DEL 5
SRR1766477.9609591 chr20 60501378 N chr20 60501454 N DEL 5
SRR1766462.3890879 chr20 60501363 N chr20 60501462 N DUP 7
SRR1766446.5126123 chr20 60500445 N chr20 60501452 N DEL 15
SRR1766480.293217 chr20 60501332 N chr20 60501533 N DEL 20
SRR1766446.5579418 chr20 60500426 N chr20 60501533 N DEL 14
SRR1766442.25071003 chr20 60500491 N chr20 60501725 N DEL 5
SRR1766457.4689944 chr20 60500394 N chr20 60501749 N DEL 7
SRR1766473.2232274 chr15 28105157 N chr15 28105424 N DUP 1
SRR1766471.791223 chr15 28105215 N chr15 28105609 N DUP 5
SRR1766456.3202608 chr15 28105413 N chr15 28106176 N DEL 3
SRR1766466.3431373 chr15 28105413 N chr15 28105880 N DEL 5
SRR1766450.8669449 chr15 28105299 N chr15 28105601 N DUP 5
SRR1766474.4644442 chr15 28105296 N chr15 28105598 N DUP 8
SRR1766464.8668271 chr15 28105375 N chr15 28105713 N DUP 6
SRR1766444.695734 chr15 28105713 N chr15 28106014 N DEL 5
SRR1766468.2056319 chr15 28105675 N chr15 28105808 N DEL 5
SRR1766482.9438526 chr15 28105750 N chr15 28105907 N DEL 5
SRR1766471.5446562 chr15 28105606 N chr15 28105979 N DEL 1
SRR1766462.5804078 chr15 28105152 N chr15 28105998 N DEL 10
SRR1766449.1065763 chr19 55508787 N chr19 55508936 N DEL 6
SRR1766483.7452266 chr19 55508787 N chr19 55508936 N DEL 6
SRR1766448.6568680 chr19 55508787 N chr19 55508936 N DEL 6
SRR1766481.7470619 chr19 55508787 N chr19 55508936 N DEL 6
SRR1766479.11341466 chr19 55508787 N chr19 55508936 N DEL 6
SRR1766442.4916245 chr19 55508787 N chr19 55508936 N DEL 6
SRR1766465.3831852 chr19 55508787 N chr19 55508862 N DEL 6
SRR1766476.143455 chr19 55508787 N chr19 55508862 N DEL 6
SRR1766485.3964972 chr19 55508787 N chr19 55508862 N DEL 6
SRR1766485.3733811 chr19 55508787 N chr19 55508936 N DEL 6
SRR1766455.2105709 chr19 55508787 N chr19 55508862 N DEL 6
SRR1766458.9377222 chr19 55508787 N chr19 55508862 N DEL 6
SRR1766462.284810 chr19 55508788 N chr19 55508863 N DEL 6
SRR1766468.782086 chr19 55508790 N chr19 55508865 N DEL 6
SRR1766473.1638037 chr19 55508799 N chr19 55508874 N DEL 3
SRR1766473.2672765 chr19 55508799 N chr19 55508874 N DEL 3
SRR1766480.6644725 chr19 55508798 N chr19 55508947 N DEL 4
SRR1766474.2741729 chr19 55508797 N chr19 55508946 N DEL 5
SRR1766458.3874377 chr19 55508817 N chr19 55508963 N DUP 5
SRR1766455.1707828 chr2 193502265 N chr2 193502346 N DUP 5
SRR1766472.7300658 chr2 193502273 N chr2 193502354 N DUP 4
SRR1766479.7237960 chr3 88436027 N chr3 88436086 N DEL 2
SRR1766484.6932937 chr3 88436022 N chr3 88436081 N DEL 4
SRR1766447.8968805 chr3 88436022 N chr3 88436081 N DEL 14
SRR1766454.8687322 chr3 88436032 N chr3 88436091 N DEL 5
