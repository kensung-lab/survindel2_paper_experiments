A00297:158:HT275DSXX:4:1556:1723:9956 chr4 179312099 N chr4 179312164 N DUP 5
A00297:158:HT275DSXX:2:2651:15872:9846 chr1 105595547 N chr1 105595634 N DEL 11
A00404:155:HV27LDSXX:1:2503:23999:12837 chr1 105595644 N chr1 105595722 N DUP 2
A00297:158:HT275DSXX:3:2304:18475:35524 chr7 158164367 N chr7 158164557 N DEL 5
A00297:158:HT275DSXX:3:1329:17680:34616 chr7 158164367 N chr7 158164557 N DEL 5
A00404:156:HV37TDSXX:3:2306:30752:13416 chr7 158164367 N chr7 158164557 N DEL 5
A00404:156:HV37TDSXX:1:2458:29695:4131 chr7 158164385 N chr7 158164573 N DUP 4
A00404:156:HV37TDSXX:2:2551:6470:10848 chr7 158164388 N chr7 158164576 N DUP 1
A00297:158:HT275DSXX:1:1212:21793:26897 chr7 158164376 N chr7 158164502 N DUP 5
A00404:156:HV37TDSXX:2:2560:19578:27038 chr7 158164502 N chr7 158164565 N DEL 5
A00404:155:HV27LDSXX:3:1609:11270:1658 chr7 158164502 N chr7 158164565 N DEL 5
A00404:156:HV37TDSXX:3:2426:7410:13698 chr7 158164502 N chr7 158164565 N DEL 5
A00404:155:HV27LDSXX:2:1238:7301:22717 chr7 158164502 N chr7 158164565 N DEL 5
A00404:155:HV27LDSXX:2:2239:9525:24158 chr7 158164502 N chr7 158164565 N DEL 5
A00297:158:HT275DSXX:3:2230:15772:18443 chr7 158164502 N chr7 158164565 N DEL 5
A00404:156:HV37TDSXX:1:2274:22254:35368 chr7 158164502 N chr7 158164565 N DEL 5
A00404:155:HV27LDSXX:4:2301:25003:2112 chr7 158164502 N chr7 158164565 N DEL 5
A00404:156:HV37TDSXX:4:2328:3929:11553 chr7 158164502 N chr7 158164565 N DEL 5
A00404:155:HV27LDSXX:2:1105:12599:22561 chr7 158164502 N chr7 158164565 N DEL 5
A00404:156:HV37TDSXX:1:2328:20555:29731 chr7 158164502 N chr7 158164565 N DEL 5
A00404:156:HV37TDSXX:2:2669:26377:1297 chr7 158164502 N chr7 158164565 N DEL 8
A00297:158:HT275DSXX:2:2209:6262:36636 chr7 158164502 N chr7 158164565 N DEL 11
A00404:155:HV27LDSXX:3:1269:9860:31219 chr7 158164502 N chr7 158164565 N DEL 26
A00404:156:HV37TDSXX:2:1209:8757:24486 chr7 158164502 N chr7 158164565 N DEL 25
A00404:155:HV27LDSXX:2:2471:13440:18850 chr7 158164502 N chr7 158164565 N DEL 24
A00297:158:HT275DSXX:4:2271:26648:3771 chr10 17629677 N chr10 17629756 N DUP 5
A00297:158:HT275DSXX:2:1105:25012:20509 chr10 17629665 N chr10 17629822 N DEL 8
A00404:155:HV27LDSXX:2:1434:29695:20134 chr16 83657986 N chr16 83658116 N DEL 15
A00297:158:HT275DSXX:3:2645:32416:5055 chr16 83658678 N chr16 83659494 N DUP 9
A00404:156:HV37TDSXX:3:2334:4327:15248 chr16 83658138 N chr16 83658678 N DEL 8
A00404:156:HV37TDSXX:1:2161:28610:9612 chr16 83658055 N chr16 83658681 N DEL 5
A00297:158:HT275DSXX:1:1446:24948:25316 chr16 83658367 N chr16 83658476 N DEL 3
A00404:156:HV37TDSXX:2:1313:19985:26177 chr16 83658367 N chr16 83658476 N DEL 3
A00404:156:HV37TDSXX:2:2513:21368:9690 chr16 83658130 N chr16 83658476 N DEL 5
A00404:155:HV27LDSXX:4:1552:8721:18317 chr16 83658101 N chr16 83658339 N DEL 5
A00404:156:HV37TDSXX:3:2334:4327:15248 chr16 83658137 N chr16 83658483 N DEL 5
A00297:158:HT275DSXX:1:2247:17155:32456 chr16 83658210 N chr16 83658556 N DEL 15
A00297:158:HT275DSXX:2:1501:28980:27070 chr16 83658135 N chr16 83658481 N DEL 5
A00404:155:HV27LDSXX:1:2546:1190:29481 chr16 83658044 N chr16 83658476 N DEL 14
A00404:155:HV27LDSXX:3:1620:28113:8030 chr16 83658404 N chr16 83658619 N DUP 2
A00404:156:HV37TDSXX:1:1605:27896:9189 chr16 83658611 N chr16 83659429 N DEL 7
A00404:156:HV37TDSXX:1:1531:23122:20369 chr16 83658096 N chr16 83658634 N DUP 10
A00404:155:HV27LDSXX:1:1376:27932:13322 chr16 83658096 N chr16 83658634 N DUP 10
A00404:156:HV37TDSXX:1:1605:27896:9189 chr16 83658096 N chr16 83658634 N DUP 10
A00404:156:HV37TDSXX:3:2436:28574:25708 chr16 83658138 N chr16 83658678 N DEL 10
A00404:155:HV27LDSXX:3:1409:8395:17002 chr16 83658138 N chr16 83658678 N DEL 7
A00404:155:HV27LDSXX:4:2442:32371:14152 chr16 83658054 N chr16 83658680 N DEL 5
A00297:158:HT275DSXX:2:2434:23041:17409 chr16 83658057 N chr16 83658683 N DEL 5
A00404:156:HV37TDSXX:2:2513:21368:9690 chr16 83658059 N chr16 83658685 N DEL 5
A00404:155:HV27LDSXX:1:1376:27932:13322 chr16 83658017 N chr16 83658686 N DEL 5
A00404:155:HV27LDSXX:1:1609:24777:29778 chr16 83658420 N chr16 83658723 N DEL 10
A00404:155:HV27LDSXX:2:2536:3613:24220 chr16 83658423 N chr16 83658769 N DEL 10
A00404:156:HV37TDSXX:2:1230:8594:8609 chr16 83658181 N chr16 83658635 N DEL 20
A00404:155:HV27LDSXX:4:2668:8287:25520 chr16 83658464 N chr16 83658894 N DUP 4
A00297:158:HT275DSXX:1:2261:12002:25034 chr16 83658409 N chr16 83658841 N DEL 5
A00297:158:HT275DSXX:1:2110:21902:8923 chr16 83658044 N chr16 83658842 N DEL 2
A00404:156:HV37TDSXX:2:2225:16369:9204 chr16 83658428 N chr16 83658492 N DUP 5
A00404:156:HV37TDSXX:3:2127:11568:28354 chr16 83658934 N chr16 83659129 N DEL 23
A00297:158:HT275DSXX:1:1608:20238:1470 chr16 83658474 N chr16 83658947 N DUP 5
A00404:155:HV27LDSXX:3:2254:22137:12524 chr16 83658167 N chr16 83658599 N DEL 5
A00297:158:HT275DSXX:3:2152:20528:11584 chr16 83658069 N chr16 83658501 N DEL 4
A00404:156:HV37TDSXX:1:1674:24587:31015 chr16 83658120 N chr16 83659303 N DUP 5
A00404:156:HV37TDSXX:1:2525:1651:6261 chr16 83659172 N chr16 83659323 N DEL 3
A00404:155:HV27LDSXX:3:1255:7636:23296 chr16 83658784 N chr16 83659299 N DUP 5
A00404:155:HV27LDSXX:3:1360:12608:35978 chr16 83659067 N chr16 83659497 N DEL 36
A00404:156:HV37TDSXX:3:2258:21224:20055 chr16 83659428 N chr16 83659515 N DEL 5
A00297:158:HT275DSXX:2:1454:31901:6042 chr16 3235758 N chr16 3235851 N DEL 10
A00297:158:HT275DSXX:3:2355:9489:15483 chr16 3235727 N chr16 3235960 N DEL 6
A00404:156:HV37TDSXX:1:2477:24270:18004 chr8 2371603 N chr8 2371822 N DUP 2
A00297:158:HT275DSXX:2:2413:11424:9064 chr8 2371698 N chr8 2371811 N DUP 7
A00404:156:HV37TDSXX:3:2447:19633:17738 chr8 2371713 N chr8 2371852 N DEL 3
A00297:158:HT275DSXX:2:1170:17662:31203 chr8 2371727 N chr8 2371866 N DEL 8
A00297:158:HT275DSXX:2:2410:25789:28620 chr6 169233631 N chr6 169233783 N DEL 5
A00297:158:HT275DSXX:3:2164:10827:7028 chr6 169233782 N chr6 169233962 N DUP 5
A00404:156:HV37TDSXX:3:2318:5077:35211 chr6 169233782 N chr6 169233962 N DUP 5
A00404:156:HV37TDSXX:2:2127:32714:34695 chr6 169233782 N chr6 169233962 N DUP 5
A00404:156:HV37TDSXX:3:2360:12943:11537 chr6 169233782 N chr6 169233962 N DUP 5
A00404:156:HV37TDSXX:3:2566:24460:24784 chr6 169233782 N chr6 169233962 N DUP 5
A00404:155:HV27LDSXX:2:1366:14696:4805 chr6 169233844 N chr6 169233968 N DEL 6
A00404:155:HV27LDSXX:2:1366:14696:4805 chr6 169233886 N chr6 169233979 N DEL 5
A00404:155:HV27LDSXX:4:1246:30969:36338 chr6 169233974 N chr6 169234097 N DUP 5
A00404:156:HV37TDSXX:4:1640:6027:8923 chr6 169233797 N chr6 169233979 N DEL 5
A00404:155:HV27LDSXX:1:2301:9679:34507 chr6 169233803 N chr6 169233985 N DEL 2
A00404:155:HV27LDSXX:3:1128:20708:33567 chr6 169233812 N chr6 169233994 N DEL 2
A00297:158:HT275DSXX:4:1262:4562:7795 chr12 20764292 N chr12 20764377 N DEL 5
A00404:156:HV37TDSXX:3:2514:19768:15875 chr12 20764292 N chr12 20764377 N DEL 15
A00404:155:HV27LDSXX:3:2666:3866:4586 chr12 20764292 N chr12 20764377 N DEL 20
A00297:158:HT275DSXX:2:1474:32786:10144 chr12 20764292 N chr12 20764377 N DEL 15
A00404:155:HV27LDSXX:4:2114:14389:31986 chr12 20764292 N chr12 20764377 N DEL 7
A00404:156:HV37TDSXX:1:1404:24722:18317 chr12 20764292 N chr12 20764377 N DEL 5
A00404:156:HV37TDSXX:4:2553:27263:19899 chr12 20764292 N chr12 20764377 N DEL 5
A00404:156:HV37TDSXX:4:2262:3947:24330 chr12 20764295 N chr12 20764380 N DEL 5
A00297:158:HT275DSXX:4:2320:28049:7983 chr12 20764377 N chr12 20764502 N DUP 5
A00297:158:HT275DSXX:1:1425:20735:7279 chr12 20764245 N chr12 20764537 N DUP 5
A00404:155:HV27LDSXX:2:1173:29098:21512 chr12 20764245 N chr12 20764537 N DUP 5
A00404:155:HV27LDSXX:3:1324:8314:14481 chr12 20764245 N chr12 20764537 N DUP 5
A00297:158:HT275DSXX:1:2251:18457:11506 chr12 20764245 N chr12 20764537 N DUP 5
A00404:156:HV37TDSXX:1:2171:22019:14325 chr12 20764245 N chr12 20764537 N DUP 5
A00404:155:HV27LDSXX:2:2649:12952:21637 chr12 20764245 N chr12 20764537 N DUP 5
A00404:155:HV27LDSXX:3:2110:30734:6120 chr12 20764245 N chr12 20764537 N DUP 5
A00297:158:HT275DSXX:3:1133:23348:33379 chr12 20764251 N chr12 20764629 N DEL 25
A00297:158:HT275DSXX:3:1655:18222:7748 chr12 20764293 N chr12 20764629 N DEL 25
A00297:158:HT275DSXX:3:2655:16333:13714 chr12 20764293 N chr12 20764629 N DEL 25
A00404:156:HV37TDSXX:4:2347:23538:32049 chr12 20764293 N chr12 20764629 N DEL 23
A00297:158:HT275DSXX:1:1540:7346:20572 chr7 156428800 N chr7 156429193 N DEL 9
A00404:155:HV27LDSXX:3:1258:2862:7138 chr7 156428877 N chr7 156429270 N DEL 5
A00404:156:HV37TDSXX:1:2145:21920:24925 chr7 156429002 N chr7 156429169 N DUP 5
A00404:156:HV37TDSXX:4:1325:4652:4163 chr7 156429151 N chr7 156429208 N DEL 15
A00404:156:HV37TDSXX:3:2133:31801:26819 chr7 156429013 N chr7 156429238 N DEL 15
A00297:158:HT275DSXX:4:1452:28953:9392 chr7 156428853 N chr7 156429246 N DEL 3
A00404:155:HV27LDSXX:1:1573:2835:29011 chr7 156429094 N chr7 156429319 N DEL 1
A00404:155:HV27LDSXX:4:2635:31222:11631 chr7 156429192 N chr7 156429417 N DEL 15
A00404:156:HV37TDSXX:2:2655:7012:13416 chr7 156428837 N chr7 156429398 N DEL 5
A00404:156:HV37TDSXX:4:1550:21287:22608 chr1 125179302 N chr1 125179424 N DEL 5
A00297:158:HT275DSXX:4:1348:6858:12399 chr1 125179356 N chr1 125179409 N DEL 10
A00404:155:HV27LDSXX:2:1308:25229:17754 chr1 125179251 N chr1 125179397 N DUP 4
A00404:156:HV37TDSXX:1:2274:23556:36526 chr1 125179351 N chr1 125179404 N DEL 56
A00404:155:HV27LDSXX:1:2367:15817:3803 chr1 125179360 N chr1 125179413 N DEL 4
A00297:158:HT275DSXX:4:2653:25726:8656 chr1 125179355 N chr1 125179408 N DEL 11
A00404:156:HV37TDSXX:2:1278:25789:18255 chr1 125179365 N chr1 125179418 N DEL 1
A00404:156:HV37TDSXX:4:1413:4607:25191 chr1 125179351 N chr1 125179404 N DEL 57
A00297:158:HT275DSXX:4:2367:12879:17347 chr9 134992321 N chr9 134992468 N DEL 10
A00404:156:HV37TDSXX:1:1521:20076:20729 chr9 134992363 N chr9 134992565 N DEL 11
A00404:155:HV27LDSXX:1:1169:17770:14231 chr9 134992291 N chr9 134992396 N DUP 1
A00404:155:HV27LDSXX:4:1140:23068:3615 chr9 134992291 N chr9 134992396 N DUP 3
A00297:158:HT275DSXX:1:1664:11993:24893 chr9 134992403 N chr9 134992605 N DUP 17
A00404:156:HV37TDSXX:4:2607:9670:19554 chr9 134992380 N chr9 134992453 N DEL 11
A00297:158:HT275DSXX:1:1543:21576:27586 chr9 134992474 N chr9 134992564 N DUP 19
A00404:155:HV27LDSXX:2:2325:5014:30624 chr9 134992496 N chr9 134992587 N DUP 10
A00404:156:HV37TDSXX:2:2214:22634:3458 chr9 134992496 N chr9 134992587 N DUP 17
A00297:158:HT275DSXX:2:2311:14498:15358 chr9 134992496 N chr9 134992587 N DUP 18
A00297:158:HT275DSXX:2:2311:14507:15374 chr9 134992496 N chr9 134992587 N DUP 18
A00297:158:HT275DSXX:1:1625:2410:34569 chr9 134992496 N chr9 134992587 N DUP 18
A00297:158:HT275DSXX:1:1625:2600:34397 chr9 134992496 N chr9 134992587 N DUP 18
A00404:156:HV37TDSXX:1:2257:32262:31939 chr9 134992515 N chr9 134992611 N DEL 13
A00404:156:HV37TDSXX:1:2257:32461:32002 chr9 134992515 N chr9 134992611 N DEL 13
A00297:158:HT275DSXX:2:1371:32425:29997 chr9 134992427 N chr9 134992536 N DEL 5
A00297:158:HT275DSXX:2:2263:4508:19820 chr16 89196407 N chr16 89196489 N DEL 1
A00404:155:HV27LDSXX:2:2256:19596:25817 chr16 89196407 N chr16 89196489 N DEL 5
A00404:156:HV37TDSXX:2:1336:14606:1391 chr16 89196407 N chr16 89196489 N DEL 5
A00404:156:HV37TDSXX:1:1115:27218:21230 chr16 89196407 N chr16 89196489 N DEL 5
A00404:155:HV27LDSXX:2:2302:8549:17644 chr16 89196407 N chr16 89196489 N DEL 5
A00404:155:HV27LDSXX:4:1412:15167:22122 chr16 89196407 N chr16 89196489 N DEL 5
A00404:155:HV27LDSXX:2:2436:29396:12947 chr16 89196414 N chr16 89196496 N DEL 8
A00404:156:HV37TDSXX:1:1161:32136:11490 chr16 89196414 N chr16 89196496 N DEL 8
A00404:156:HV37TDSXX:4:1529:8910:24721 chr16 89196414 N chr16 89196496 N DEL 8
A00297:158:HT275DSXX:3:2546:26449:26506 chr3 114303654 N chr3 114303749 N DEL 12
A00297:158:HT275DSXX:4:2333:13955:12101 chr3 114303657 N chr3 114303752 N DEL 10
A00404:156:HV37TDSXX:2:1612:11360:7983 chr3 114303654 N chr3 114303749 N DEL 18
A00404:156:HV37TDSXX:2:1617:10556:13604 chr3 114303655 N chr3 114303750 N DEL 12
A00297:158:HT275DSXX:1:2227:22327:20932 chr3 114303654 N chr3 114303749 N DEL 13
A00404:155:HV27LDSXX:1:1169:20934:26913 chr3 114303656 N chr3 114303751 N DEL 11
A00404:155:HV27LDSXX:3:2565:28013:30154 chr3 114303654 N chr3 114303749 N DEL 14
A00404:156:HV37TDSXX:1:2205:4083:25003 chr3 114303654 N chr3 114303749 N DEL 14
A00404:156:HV37TDSXX:1:2205:4173:25097 chr3 114303654 N chr3 114303749 N DEL 14
A00297:158:HT275DSXX:3:2436:13042:15405 chr3 114303722 N chr3 114303773 N DEL 5
A00404:155:HV27LDSXX:3:1463:16721:21245 chr3 114303722 N chr3 114303773 N DEL 5
A00404:155:HV27LDSXX:2:1475:20057:29778 chr3 153646744 N chr3 153646832 N DEL 10
A00404:156:HV37TDSXX:4:1510:17653:7106 chr3 153646744 N chr3 153646832 N DEL 12
A00404:155:HV27LDSXX:3:2506:13711:21543 chr3 153646744 N chr3 153646832 N DEL 14
A00297:158:HT275DSXX:2:2316:21576:1939 chr3 153646689 N chr3 153646846 N DEL 1
A00297:158:HT275DSXX:4:2115:9326:10222 chr3 153646753 N chr3 153646841 N DEL 6
A00404:156:HV37TDSXX:2:1250:19144:19085 chr3 153646747 N chr3 153646835 N DEL 12
A00404:155:HV27LDSXX:2:2537:30879:13103 chr3 153646753 N chr3 153646841 N DEL 9
A00404:155:HV27LDSXX:3:1554:17987:1423 chr22 44732996 N chr22 44733174 N DEL 10
A00404:155:HV27LDSXX:3:2374:27534:15139 chr6 147616281 N chr6 147616330 N DUP 10
A00297:158:HT275DSXX:1:1636:25852:30827 chr6 147616287 N chr6 147616361 N DUP 10
A00404:156:HV37TDSXX:3:2149:4933:36839 chr6 147616287 N chr6 147616361 N DUP 10
A00404:156:HV37TDSXX:4:1636:27281:36245 chr6 147616287 N chr6 147616361 N DUP 10
A00297:158:HT275DSXX:3:2577:11966:9596 chr6 147616287 N chr6 147616361 N DUP 10
A00297:158:HT275DSXX:4:1461:21287:30060 chr6 147616287 N chr6 147616361 N DUP 10
A00404:156:HV37TDSXX:3:2109:17273:23516 chr6 147616287 N chr6 147616386 N DUP 6
A00404:156:HV37TDSXX:2:1434:9869:28855 chr6 147616287 N chr6 147616386 N DUP 8
A00404:156:HV37TDSXX:4:2272:14696:19429 chr6 147616376 N chr6 147616438 N DEL 13
A00297:158:HT275DSXX:3:1140:32922:32612 chr6 147616287 N chr6 147616386 N DUP 9
A00404:155:HV27LDSXX:2:2504:12653:34147 chr6 147616287 N chr6 147616361 N DUP 10
A00404:155:HV27LDSXX:4:1420:15609:13182 chr6 147616412 N chr6 147616474 N DEL 21
A00404:155:HV27LDSXX:4:1578:6976:17550 chr6 147616326 N chr6 147616438 N DEL 16
A00404:155:HV27LDSXX:2:1541:18376:36479 chr6 147616337 N chr6 147616474 N DEL 19
A00297:158:HT275DSXX:3:1255:11831:6261 chr6 147616337 N chr6 147616474 N DEL 12
A00297:158:HT275DSXX:3:2635:16758:16423 chr6 147616337 N chr6 147616474 N DEL 5
A00297:158:HT275DSXX:4:2625:7663:20400 chr6 147616312 N chr6 147616474 N DEL 5
A00404:156:HV37TDSXX:3:2617:7374:34209 chr6 147616312 N chr6 147616474 N DEL 5
A00404:155:HV27LDSXX:4:1443:19714:9612 chr6 147616312 N chr6 147616474 N DEL 5
A00297:158:HT275DSXX:2:1560:23321:5776 chr6 147616299 N chr6 147616486 N DEL 3
A00404:156:HV37TDSXX:1:2501:15872:14418 chr1 234247696 N chr1 234248145 N DEL 2
A00404:156:HV37TDSXX:1:1623:24316:21026 chr1 234247696 N chr1 234248145 N DEL 2
A00404:155:HV27LDSXX:1:2170:15447:31062 chr1 234247696 N chr1 234248145 N DEL 5
A00404:156:HV37TDSXX:1:1201:25934:20666 chr1 234247696 N chr1 234248145 N DEL 5
A00404:156:HV37TDSXX:1:1201:26612:21277 chr1 234247696 N chr1 234248145 N DEL 5
A00404:156:HV37TDSXX:4:2569:3314:3192 chr1 234247696 N chr1 234248145 N DEL 5
A00297:158:HT275DSXX:1:1431:25003:11976 chr1 234247696 N chr1 234248145 N DEL 5
A00297:158:HT275DSXX:2:2236:20030:22341 chr1 234247696 N chr1 234248145 N DEL 5
A00297:158:HT275DSXX:4:2165:21585:12508 chr1 234247696 N chr1 234248145 N DEL 5
A00297:158:HT275DSXX:4:2165:26530:31344 chr1 234247696 N chr1 234248145 N DEL 5
A00297:158:HT275DSXX:1:1110:21224:9752 chr1 234247709 N chr1 234248158 N DEL 5
A00297:158:HT275DSXX:4:2454:18674:9283 chr1 234247696 N chr1 234248145 N DEL 5
A00404:155:HV27LDSXX:1:1427:11360:24205 chr1 234247720 N chr1 234248167 N DUP 5
A00297:158:HT275DSXX:4:1268:11487:25582 chr1 234247721 N chr1 234248168 N DUP 5
A00404:155:HV27LDSXX:4:1276:21784:10629 chr1 234247725 N chr1 234248172 N DUP 2
A00404:156:HV37TDSXX:3:2423:8657:9283 chr1 234247838 N chr1 234248511 N DEL 5
A00404:156:HV37TDSXX:1:2501:15872:14418 chr1 234247569 N chr1 234247798 N DEL 5
A00297:158:HT275DSXX:1:2663:27172:5212 chr1 234247843 N chr1 234247926 N DUP 1
A00297:158:HT275DSXX:2:2308:10113:4100 chr1 234247843 N chr1 234247926 N DUP 1
A00404:155:HV27LDSXX:1:1640:9851:5024 chr1 234247843 N chr1 234247926 N DUP 1
A00297:158:HT275DSXX:2:2159:1895:15076 chr1 234247926 N chr1 234248291 N DEL 5
A00404:155:HV27LDSXX:4:1623:28519:33317 chr1 234247926 N chr1 234248515 N DEL 5
A00404:155:HV27LDSXX:1:1275:22733:10739 chr1 234247514 N chr1 234247939 N DEL 35
A00404:156:HV37TDSXX:4:1567:20862:36119 chr1 234247964 N chr1 234248579 N DUP 35
A00297:158:HT275DSXX:1:2609:1461:21590 chr1 234247964 N chr1 234248579 N DUP 40
A00297:158:HT275DSXX:1:2609:1506:21386 chr1 234247964 N chr1 234248579 N DUP 40
A00404:156:HV37TDSXX:1:1442:13015:36432 chr1 234247964 N chr1 234248579 N DUP 40
A00297:158:HT275DSXX:4:1654:26973:9032 chr1 234247964 N chr1 234248579 N DUP 37
A00297:158:HT275DSXX:1:1320:20329:9925 chr1 234248055 N chr1 234248474 N DUP 49
A00404:155:HV27LDSXX:1:1204:11840:33144 chr1 234248055 N chr1 234248474 N DUP 43
A00404:155:HV27LDSXX:1:1205:14850:2628 chr1 234248055 N chr1 234248474 N DUP 43
A00404:155:HV27LDSXX:1:1355:24858:29450 chr1 234248055 N chr1 234248474 N DUP 35
A00404:155:HV27LDSXX:1:1444:1054:26459 chr1 234248055 N chr1 234248474 N DUP 35
A00297:158:HT275DSXX:4:2508:21414:31501 chr1 234248055 N chr1 234248474 N DUP 35
A00297:158:HT275DSXX:2:2543:18439:2581 chr1 234248055 N chr1 234248474 N DUP 35
A00297:158:HT275DSXX:2:1416:24758:33786 chr1 234247602 N chr1 234248055 N DEL 25
A00404:156:HV37TDSXX:4:2156:12246:14810 chr1 234247602 N chr1 234248055 N DEL 35
A00404:155:HV27LDSXX:3:1150:21838:35806 chr1 234247602 N chr1 234248055 N DEL 22
A00297:158:HT275DSXX:1:2641:9896:12712 chr1 234247602 N chr1 234248055 N DEL 15
A00404:155:HV27LDSXX:1:2331:19235:17049 chr1 234247602 N chr1 234248055 N DEL 23
A00297:158:HT275DSXX:1:2523:29243:33004 chr1 234247602 N chr1 234248055 N DEL 15
A00404:156:HV37TDSXX:1:1343:5285:14278 chr1 234247602 N chr1 234248055 N DEL 15
A00404:155:HV27LDSXX:1:1632:6668:5055 chr1 234247712 N chr1 234248159 N DUP 3
A00404:156:HV37TDSXX:2:2250:3821:28995 chr1 234247589 N chr1 234248070 N DEL 5
A00404:156:HV37TDSXX:3:1624:5638:8531 chr1 234247589 N chr1 234248070 N DEL 5
A00404:156:HV37TDSXX:3:2423:8657:9283 chr1 234247626 N chr1 234248075 N DEL 2
A00297:158:HT275DSXX:2:1276:17400:19883 chr1 234247712 N chr1 234248159 N DUP 5
A00297:158:HT275DSXX:1:2510:29758:9220 chr1 234247712 N chr1 234248159 N DUP 5
A00297:158:HT275DSXX:3:1265:21667:28995 chr1 234247712 N chr1 234248159 N DUP 5
A00297:158:HT275DSXX:1:2418:26006:26177 chr1 234247712 N chr1 234248159 N DUP 5
A00404:156:HV37TDSXX:2:2365:7789:30107 chr1 234247712 N chr1 234248159 N DUP 5
A00404:155:HV27LDSXX:2:1353:30092:30686 chr1 234247712 N chr1 234248159 N DUP 5
A00404:155:HV27LDSXX:1:2249:18710:7874 chr1 234247712 N chr1 234248159 N DUP 5
A00404:155:HV27LDSXX:4:1157:8052:30405 chr1 234247712 N chr1 234248159 N DUP 5
A00404:155:HV27LDSXX:2:2355:10646:36182 chr1 234247712 N chr1 234248159 N DUP 5
A00297:158:HT275DSXX:1:1411:28076:24752 chr1 234247712 N chr1 234248159 N DUP 5
A00404:156:HV37TDSXX:1:2128:9326:31955 chr1 234247712 N chr1 234248159 N DUP 5
A00404:156:HV37TDSXX:4:2172:13395:19241 chr1 234247712 N chr1 234248159 N DUP 5
A00297:158:HT275DSXX:1:1207:22670:14669 chr1 234247712 N chr1 234248159 N DUP 5
A00297:158:HT275DSXX:1:1221:23348:27148 chr1 234247712 N chr1 234248159 N DUP 5
A00297:158:HT275DSXX:4:1654:26973:9032 chr1 234247712 N chr1 234248159 N DUP 5
A00404:156:HV37TDSXX:2:2244:27859:4993 chr1 234247712 N chr1 234248159 N DUP 5
A00404:156:HV37TDSXX:2:2644:24108:9518 chr1 234247712 N chr1 234248159 N DUP 5
A00404:155:HV27LDSXX:4:1608:14733:5118 chr1 234247712 N chr1 234248159 N DUP 5
A00404:156:HV37TDSXX:2:1332:29894:14653 chr1 234247712 N chr1 234248159 N DUP 5
A00297:158:HT275DSXX:3:2560:18394:2973 chr1 234247712 N chr1 234248159 N DUP 5
A00404:156:HV37TDSXX:1:1441:16269:1767 chr1 234247972 N chr1 234248279 N DUP 5
A00404:155:HV27LDSXX:2:1615:28818:20369 chr1 234247647 N chr1 234248180 N DEL 4
A00404:156:HV37TDSXX:3:1161:31629:8422 chr1 234247831 N chr1 234248560 N DEL 5
A00404:156:HV37TDSXX:1:1441:16269:1767 chr1 234247831 N chr1 234248560 N DEL 5
A00297:158:HT275DSXX:1:1320:20329:9925 chr1 234247831 N chr1 234248560 N DEL 5
A00404:155:HV27LDSXX:4:1540:3341:3208 chr1 234247831 N chr1 234248560 N DEL 5
A00297:158:HT275DSXX:2:2420:17734:19179 chr1 234247831 N chr1 234248560 N DEL 6
A00404:155:HV27LDSXX:2:1354:18493:24064 chr1 234247838 N chr1 234248511 N DEL 1
A00404:155:HV27LDSXX:2:2142:11605:8093 chr1 234247838 N chr1 234248511 N DEL 5
A00404:155:HV27LDSXX:2:2651:24053:9361 chr1 234247838 N chr1 234248511 N DEL 5
A00297:158:HT275DSXX:1:2609:1506:21386 chr1 234247838 N chr1 234248511 N DEL 5
A00297:158:HT275DSXX:4:2268:5339:25739 chr1 234247831 N chr1 234248560 N DEL 10
A00404:155:HV27LDSXX:4:2429:30725:33223 chr1 234247831 N chr1 234248560 N DEL 10
A00404:156:HV37TDSXX:2:2421:23800:12587 chr1 234247905 N chr1 234248270 N DEL 10
A00297:158:HT275DSXX:4:2508:21414:31501 chr1 234247831 N chr1 234248560 N DEL 19
A00404:156:HV37TDSXX:2:2250:3821:28995 chr1 234247831 N chr1 234248560 N DEL 19
A00404:156:HV37TDSXX:1:2366:13991:2331 chr1 234248011 N chr1 234248402 N DUP 2
A00404:155:HV27LDSXX:2:2251:13774:29324 chr1 234248011 N chr1 234248402 N DUP 4
A00404:156:HV37TDSXX:1:1178:7880:10003 chr1 234248347 N chr1 234248570 N DUP 5
A00404:155:HV27LDSXX:4:1540:3341:3208 chr1 234247982 N chr1 234248347 N DEL 5
A00297:158:HT275DSXX:2:1169:13141:5118 chr1 234248073 N chr1 234248464 N DUP 9
A00297:158:HT275DSXX:3:2428:1244:4272 chr1 234248073 N chr1 234248464 N DUP 13
A00297:158:HT275DSXX:1:1207:22670:14669 chr1 234248459 N chr1 234248626 N DUP 27
A00404:156:HV37TDSXX:1:2235:20745:7169 chr1 234248459 N chr1 234248682 N DUP 30
A00297:158:HT275DSXX:4:1363:7681:12132 chr1 234248459 N chr1 234248570 N DUP 25
A00404:156:HV37TDSXX:3:2356:5990:7701 chr1 234248010 N chr1 234248459 N DEL 23
A00404:155:HV27LDSXX:1:1136:19307:17049 chr1 234247982 N chr1 234248459 N DEL 16
A00404:156:HV37TDSXX:3:2669:15383:23970 chr1 234247991 N chr1 234248468 N DEL 6
A00404:155:HV27LDSXX:4:2656:1588:19867 chr1 234248473 N chr1 234248584 N DUP 1
A00404:156:HV37TDSXX:2:1332:29894:14653 chr1 234248518 N chr1 234248629 N DUP 10
A00404:155:HV27LDSXX:1:2354:27633:12680 chr1 234248528 N chr1 234248583 N DUP 4
A00297:158:HT275DSXX:1:1221:23348:27148 chr1 234248528 N chr1 234248583 N DUP 4
A00404:156:HV37TDSXX:2:1632:7545:31876 chr1 234247574 N chr1 234248531 N DEL 3
A00297:158:HT275DSXX:3:1248:31412:3912 chr1 234248540 N chr1 234248651 N DUP 11
A00404:156:HV37TDSXX:4:2672:13051:15640 chr1 234248484 N chr1 234248651 N DUP 11
A00404:155:HV27LDSXX:2:2523:11822:36558 chr1 234248459 N chr1 234248682 N DUP 32
A00404:156:HV37TDSXX:4:2508:11035:4257 chr1 234248459 N chr1 234248682 N DUP 30
A00297:158:HT275DSXX:3:1427:3052:7185 chr1 234248459 N chr1 234248682 N DUP 26
A00297:158:HT275DSXX:3:2428:1244:4272 chr1 234248459 N chr1 234248682 N DUP 16
A00404:155:HV27LDSXX:4:1608:14733:5118 chr1 234248466 N chr1 234248689 N DUP 20
A00404:155:HV27LDSXX:1:2331:19235:17049 chr1 234247856 N chr1 234248529 N DEL 6
A00404:156:HV37TDSXX:3:1407:18810:19570 chr1 234247832 N chr1 234248561 N DEL 12
A00404:156:HV37TDSXX:1:2128:9326:31955 chr1 234247836 N chr1 234248565 N DEL 8
A00297:158:HT275DSXX:1:2641:9896:12712 chr1 234248540 N chr1 234248651 N DUP 1
A00404:155:HV27LDSXX:4:1513:5683:36417 chr1 234248540 N chr1 234248651 N DUP 3
A00297:158:HT275DSXX:4:1476:27742:31344 chr1 234248540 N chr1 234248651 N DUP 6
A00404:155:HV27LDSXX:4:2429:30725:33223 chr1 234248540 N chr1 234248651 N DUP 9
A00404:155:HV27LDSXX:2:1353:30092:30686 chr1 234247836 N chr1 234248621 N DEL 15
A00404:156:HV37TDSXX:3:1407:18810:19570 chr1 234248595 N chr1 234248652 N DEL 5
A00404:156:HV37TDSXX:4:2672:13051:15640 chr1 234248539 N chr1 234248652 N DEL 15
A00404:156:HV37TDSXX:1:1224:30237:19539 chr1 234248595 N chr1 234248652 N DEL 5
A00404:156:HV37TDSXX:3:1464:14009:11224 chr1 234247556 N chr1 234248653 N DEL 5
A00404:156:HV37TDSXX:1:2236:25238:20932 chr5 1212110 N chr5 1212170 N DEL 2
A00297:158:HT275DSXX:4:2652:7952:34115 chr5 1211956 N chr5 1212119 N DEL 7
A00404:156:HV37TDSXX:4:2469:1127:33505 chr5 1211956 N chr5 1212119 N DEL 7
A00404:156:HV37TDSXX:1:2460:27073:3881 chr5 1211959 N chr5 1212122 N DEL 7
A00404:156:HV37TDSXX:4:1354:18367:34397 chr10 12276933 N chr10 12277159 N DEL 2
A00404:155:HV27LDSXX:2:2306:12897:16720 chr10 12276933 N chr10 12277159 N DEL 4
A00404:155:HV27LDSXX:3:2318:26485:13135 chr10 12276933 N chr10 12277159 N DEL 4
A00404:156:HV37TDSXX:3:2444:14995:12399 chr10 12276933 N chr10 12277159 N DEL 4
A00404:155:HV27LDSXX:3:1604:2058:34334 chr10 12277112 N chr10 12277339 N DUP 2
A00404:155:HV27LDSXX:1:2131:3179:27164 chr10 12277116 N chr10 12277343 N DUP 3
A00297:158:HT275DSXX:3:2349:27001:8641 chr15 82703481 N chr15 82703546 N DUP 21
A00297:158:HT275DSXX:2:2574:32154:35697 chr11 69324721 N chr11 69325111 N DEL 5
A00404:155:HV27LDSXX:1:2577:4336:17456 chr11 69324608 N chr11 69324686 N DEL 2
A00297:158:HT275DSXX:3:1204:5936:16031 chr11 69324502 N chr11 69324808 N DUP 5
A00297:158:HT275DSXX:1:1272:31973:1157 chr11 69324850 N chr11 69325144 N DEL 2
A00404:155:HV27LDSXX:3:1243:1262:15640 chr11 69324868 N chr11 69325160 N DUP 5
A00297:158:HT275DSXX:3:2547:5122:5916 chr11 69324499 N chr11 69324870 N DEL 5
A00297:158:HT275DSXX:2:2471:7491:25081 chr11 69324703 N chr11 69325093 N DEL 15
A00404:156:HV37TDSXX:4:1101:8458:7905 chr11 69324457 N chr11 69325199 N DEL 5
A00404:155:HV27LDSXX:4:1333:22571:10426 chr5 152698319 N chr5 152698387 N DEL 9
A00297:158:HT275DSXX:2:2606:32542:6308 chr2 61848953 N chr2 61849066 N DEL 1
A00404:156:HV37TDSXX:3:1258:2871:1767 chr2 61848951 N chr2 61849024 N DEL 5
A00404:156:HV37TDSXX:3:1258:2899:1846 chr2 61848951 N chr2 61849024 N DEL 5
A00404:155:HV27LDSXX:1:2439:27733:1423 chr2 61848951 N chr2 61849078 N DEL 12
A00404:156:HV37TDSXX:2:2571:23339:16423 chr2 61848953 N chr2 61849066 N DEL 5
A00297:158:HT275DSXX:4:2277:30987:16110 chr2 61848953 N chr2 61849066 N DEL 5
A00404:155:HV27LDSXX:1:2439:27733:1423 chr2 61849032 N chr2 61849125 N DEL 8
A00404:155:HV27LDSXX:2:2127:8024:13009 chr2 61849011 N chr2 61849168 N DEL 17
A00297:158:HT275DSXX:4:2417:22254:27477 chr2 61849190 N chr2 61849245 N DEL 24
A00404:155:HV27LDSXX:4:2267:28058:3834 chr2 61849192 N chr2 61849247 N DEL 23
A00404:155:HV27LDSXX:4:2267:28248:3724 chr2 61849192 N chr2 61849247 N DEL 23
A00404:156:HV37TDSXX:3:2161:11424:15295 chr2 61849003 N chr2 61849164 N DEL 7
A00297:158:HT275DSXX:3:2332:30318:24377 chr2 61849065 N chr2 61849220 N DEL 28
A00404:155:HV27LDSXX:1:2140:8097:29543 chr2 61849065 N chr2 61849220 N DEL 17
A00297:158:HT275DSXX:3:1326:3269:11005 chr2 61849065 N chr2 61849220 N DEL 17
A00297:158:HT275DSXX:4:1655:2682:25520 chr2 61849165 N chr2 61849220 N DEL 16
A00404:156:HV37TDSXX:4:2546:14163:10770 chr2 61849190 N chr2 61849245 N DEL 25
A00404:156:HV37TDSXX:4:1119:2031:35321 chr2 61849190 N chr2 61849245 N DEL 24
A00404:156:HV37TDSXX:3:2370:20708:13870 chr2 61849160 N chr2 61849245 N DEL 20
A00404:156:HV37TDSXX:1:2354:11035:7138 chr2 61849160 N chr2 61849245 N DEL 19
A00404:156:HV37TDSXX:4:2225:29631:16266 chr2 61849066 N chr2 61849221 N DEL 14
A00297:158:HT275DSXX:1:1528:16658:28776 chr2 61849047 N chr2 61849232 N DEL 3
A00297:158:HT275DSXX:1:1528:17119:30577 chr2 61849047 N chr2 61849232 N DEL 3
A00297:158:HT275DSXX:3:2275:14859:28980 chr2 61849060 N chr2 61849245 N DEL 7
A00404:155:HV27LDSXX:2:2134:24325:33880 chr2 61849060 N chr2 61849245 N DEL 8
A00404:156:HV37TDSXX:3:2231:24569:8218 chr2 61849060 N chr2 61849245 N DEL 10
A00297:158:HT275DSXX:3:1211:9751:35289 chr2 61848974 N chr2 61849253 N DEL 5
A00297:158:HT275DSXX:1:2526:10547:10614 chr20 35084697 N chr20 35084794 N DEL 3
A00297:158:HT275DSXX:4:1544:32850:23062 chr20 35084697 N chr20 35084794 N DEL 3
A00297:158:HT275DSXX:2:2116:6244:19820 chr20 35084697 N chr20 35084794 N DEL 5
A00404:156:HV37TDSXX:1:2573:17915:22122 chr20 35084697 N chr20 35084794 N DEL 5
A00404:155:HV27LDSXX:2:2177:20672:8891 chr20 35084697 N chr20 35084794 N DEL 5
A00404:156:HV37TDSXX:1:1314:15817:7059 chr20 35084697 N chr20 35084794 N DEL 5
A00297:158:HT275DSXX:2:1317:2672:36307 chr20 35084697 N chr20 35084794 N DEL 5
A00297:158:HT275DSXX:3:2327:7048:4836 chr20 35084697 N chr20 35084794 N DEL 5
A00404:156:HV37TDSXX:4:1129:9299:30812 chr20 35084729 N chr20 35084794 N DEL 5
A00297:158:HT275DSXX:3:1123:3504:3615 chr20 35084729 N chr20 35084794 N DEL 5
A00404:155:HV27LDSXX:2:1136:26693:13620 chr20 35084729 N chr20 35084794 N DEL 5
A00297:158:HT275DSXX:1:1251:26883:11757 chr20 35084729 N chr20 35084794 N DEL 5
A00404:155:HV27LDSXX:1:2271:2980:20588 chr20 35084729 N chr20 35084794 N DEL 5
A00404:155:HV27LDSXX:2:2450:2474:30639 chr20 35084686 N chr20 35084749 N DUP 5
A00404:155:HV27LDSXX:4:1466:7527:35258 chr20 35084686 N chr20 35084749 N DUP 5
A00404:155:HV27LDSXX:2:2450:3495:31125 chr20 35084686 N chr20 35084749 N DUP 5
A00297:158:HT275DSXX:2:2303:1389:7748 chr20 35084686 N chr20 35084749 N DUP 5
A00404:155:HV27LDSXX:4:1348:15673:18458 chr20 35084729 N chr20 35084794 N DEL 5
A00404:155:HV27LDSXX:4:1348:15682:18474 chr20 35084729 N chr20 35084794 N DEL 5
A00404:155:HV27LDSXX:2:1330:20148:9111 chr20 35084729 N chr20 35084794 N DEL 5
A00404:155:HV27LDSXX:4:2605:5746:29293 chr20 35084729 N chr20 35084794 N DEL 5
A00297:158:HT275DSXX:1:2649:3893:27555 chr20 35084729 N chr20 35084794 N DEL 5
A00404:155:HV27LDSXX:1:1647:17490:18004 chr20 35084729 N chr20 35084794 N DEL 5
A00404:156:HV37TDSXX:1:1547:13675:1094 chr20 35084729 N chr20 35084794 N DEL 5
A00297:158:HT275DSXX:3:1134:5339:19789 chr20 35084732 N chr20 35084797 N DEL 5
A00404:155:HV27LDSXX:1:2568:5945:8187 chr20 35084700 N chr20 35084797 N DEL 5
A00297:158:HT275DSXX:1:1272:28565:24377 chr20 35084703 N chr20 35084800 N DEL 5
A00404:155:HV27LDSXX:3:1374:4372:28667 chr20 35084704 N chr20 35084801 N DEL 5
A00297:158:HT275DSXX:4:2551:12409:16501 chr20 35084705 N chr20 35084802 N DEL 5
A00404:156:HV37TDSXX:4:1658:1334:27853 chr20 35084707 N chr20 35084804 N DEL 5
A00404:156:HV37TDSXX:4:2521:27208:22216 chr4 60510652 N chr4 60510707 N DEL 20
A00404:156:HV37TDSXX:1:1217:16477:34194 chr16 57569789 N chr16 57569857 N DUP 5
A00404:155:HV27LDSXX:4:1153:20618:9017 chr16 57569701 N chr16 57569999 N DEL 4
A00404:156:HV37TDSXX:1:2546:22679:22357 chrX 87465994 N chrX 87466186 N DUP 5
A00297:158:HT275DSXX:1:1655:9778:32925 chr19 2991048 N chr19 2991405 N DUP 10
A00404:155:HV27LDSXX:2:1353:23927:30123 chr19 2991190 N chr19 2991535 N DEL 5
A00404:156:HV37TDSXX:3:2468:29451:2895 chr19 2991190 N chr19 2991535 N DEL 5
A00404:155:HV27LDSXX:2:1526:6596:27320 chr19 2991207 N chr19 2991550 N DUP 5
A00404:155:HV27LDSXX:2:2526:7202:5509 chr19 2991207 N chr19 2991550 N DUP 5
A00404:156:HV37TDSXX:2:1676:27335:35681 chr19 2991211 N chr19 2991554 N DUP 2
A00404:155:HV27LDSXX:2:2349:30689:6198 chr11 62656120 N chr11 62656286 N DEL 16
A00404:156:HV37TDSXX:1:2416:29631:22561 chrX 108141075 N chrX 108141168 N DUP 3
A00404:155:HV27LDSXX:4:2131:17770:21465 chr15 89746816 N chr15 89747065 N DEL 5
A00404:155:HV27LDSXX:4:2131:17960:21073 chr15 89746830 N chr15 89747005 N DEL 5
A00297:158:HT275DSXX:2:1206:5972:10864 chr15 89746657 N chr15 89746988 N DUP 1
A00297:158:HT275DSXX:2:1550:24478:21371 chr15 89746717 N chr15 89746872 N DEL 7
A00404:155:HV27LDSXX:4:1319:23421:32471 chr10 51393162 N chr10 51393594 N DEL 5
A00404:155:HV27LDSXX:3:1138:22390:5040 chr1 9155321 N chr1 9155650 N DEL 2
A00404:156:HV37TDSXX:3:1666:14597:1971 chr1 9155123 N chr1 9155327 N DEL 3
A00404:156:HV37TDSXX:3:2526:21739:23923 chr1 9155125 N chr1 9155329 N DEL 2
A00404:156:HV37TDSXX:4:1470:25238:24126 chr1 9155378 N chr1 9155705 N DUP 5
A00404:155:HV27LDSXX:1:2659:19976:22435 chr1 9155459 N chr1 9155788 N DEL 5
A00404:155:HV27LDSXX:2:1175:16134:18505 chr1 9155627 N chr1 9155792 N DEL 5
A00404:156:HV37TDSXX:3:1302:13512:8516 chr1 9155773 N chr1 9155854 N DUP 10
A00297:158:HT275DSXX:3:2542:12527:33051 chr1 9155362 N chr1 9155650 N DEL 5
A00297:158:HT275DSXX:4:1615:32642:4225 chr1 9155123 N chr1 9155655 N DEL 5
A00297:158:HT275DSXX:4:1547:19750:22921 chr1 9155377 N chr1 9155706 N DEL 5
A00297:158:HT275DSXX:1:1357:5041:10254 chr1 9155125 N chr1 9155739 N DEL 5
A00297:158:HT275DSXX:1:1502:15329:17143 chr1 9155828 N chr1 9156034 N DEL 2
A00297:158:HT275DSXX:1:2209:1949:16360 chr1 9155828 N chr1 9156034 N DEL 2
A00297:158:HT275DSXX:1:1202:2636:19648 chr1 9155837 N chr1 9155920 N DEL 5
A00404:155:HV27LDSXX:3:2164:27814:32377 chr1 9155303 N chr1 9155919 N DEL 5
A00297:158:HT275DSXX:1:2626:26187:18662 chr1 9155303 N chr1 9155919 N DEL 5
A00404:156:HV37TDSXX:2:2359:12373:15468 chr1 9155133 N chr1 9155870 N DEL 5
A00404:155:HV27LDSXX:2:1269:23375:27445 chr1 9155468 N chr1 9155797 N DEL 15
A00404:155:HV27LDSXX:2:1175:16134:18505 chr1 9155302 N chr1 9155959 N DEL 5
A00297:158:HT275DSXX:2:2643:18584:6464 chr1 9155388 N chr1 9155963 N DEL 5
A00297:158:HT275DSXX:3:2538:25192:19820 chr1 9155837 N chr1 9156043 N DEL 10
A00404:156:HV37TDSXX:4:1553:4960:36699 chr19 41432855 N chr19 41432941 N DEL 7
A00404:156:HV37TDSXX:1:2533:17644:3333 chr19 41432824 N chr19 41432967 N DUP 19
A00404:156:HV37TDSXX:1:2533:17743:6386 chr19 41432824 N chr19 41432967 N DUP 9
A00297:158:HT275DSXX:3:1141:4517:23093 chr19 41432731 N chr19 41432868 N DEL 3
A00404:156:HV37TDSXX:4:1553:4960:36699 chr19 41432800 N chr19 41432933 N DEL 11
A00404:155:HV27LDSXX:3:2227:20491:35822 chr3 169378535 N chr3 169378665 N DEL 4
A00297:158:HT275DSXX:2:2501:19804:21042 chr3 169378568 N chr3 169378637 N DEL 27
A00404:155:HV27LDSXX:1:1574:25111:26569 chr3 169378672 N chr3 169378735 N DUP 21
A00404:156:HV37TDSXX:2:1547:15411:35070 chr3 169378595 N chr3 169378663 N DEL 27
A00404:155:HV27LDSXX:3:2227:20482:35806 chr3 169378599 N chr3 169378741 N DEL 10
A00404:155:HV27LDSXX:3:2227:20491:35822 chr3 169378599 N chr3 169378741 N DEL 10
A00297:158:HT275DSXX:3:2367:3088:3646 chr3 169378591 N chr3 169378741 N DEL 10
A00404:155:HV27LDSXX:3:1261:1163:33442 chr3 169378587 N chr3 169378741 N DEL 10
A00404:155:HV27LDSXX:3:1261:1787:32142 chr3 169378587 N chr3 169378741 N DEL 10
A00297:158:HT275DSXX:4:2276:21983:24189 chr3 169378587 N chr3 169378741 N DEL 10
A00404:155:HV27LDSXX:1:2528:29107:2988 chr3 169378571 N chr3 169378737 N DEL 5
A00297:158:HT275DSXX:1:2457:24912:5776 chr3 169378575 N chr3 169378741 N DEL 10
A00404:155:HV27LDSXX:1:2541:31828:17660 chr3 169378571 N chr3 169378737 N DEL 5
A00404:155:HV27LDSXX:1:2161:20166:26428 chr3 169378563 N chr3 169378741 N DEL 10
A00297:158:HT275DSXX:4:2360:25563:2957 chr3 169378559 N chr3 169378741 N DEL 10
A00297:158:HT275DSXX:4:2667:27534:20870 chr3 169378555 N chr3 169378741 N DEL 10
A00404:156:HV37TDSXX:2:1252:13720:33739 chr3 169378551 N chr3 169378741 N DEL 10
A00404:156:HV37TDSXX:3:2338:29206:10019 chr9 134714628 N chr9 134714757 N DUP 4
A00404:156:HV37TDSXX:1:2230:16866:29825 chr9 134714811 N chr9 134715057 N DEL 5
A00404:156:HV37TDSXX:2:2271:27697:2769 chr9 134714787 N chr9 134714949 N DEL 8
A00404:155:HV27LDSXX:1:2460:27172:17300 chr9 134714775 N chr9 134714888 N DUP 17
A00404:156:HV37TDSXX:1:2464:20410:29731 chr9 134714750 N chr9 134714904 N DUP 2
A00404:155:HV27LDSXX:4:1552:9182:22028 chr9 134714422 N chr9 134714788 N DEL 8
A00404:156:HV37TDSXX:2:2271:27697:2769 chr9 134714702 N chr9 134714949 N DEL 16
A00404:156:HV37TDSXX:4:2364:22688:20462 chr9 134714827 N chr9 134714986 N DEL 5
A00404:155:HV27LDSXX:4:2522:2022:17080 chr9 134714794 N chr9 134715067 N DEL 5
A00297:158:HT275DSXX:1:1527:30047:36965 chr13 110558529 N chr13 110558844 N DEL 1
A00297:158:HT275DSXX:1:1528:30653:6198 chr13 110558529 N chr13 110558844 N DEL 1
A00404:155:HV27LDSXX:2:1166:11189:21652 chr13 110558529 N chr13 110558845 N DEL 9
A00297:158:HT275DSXX:1:2569:14100:33332 chr13 110558529 N chr13 110558845 N DEL 9
A00297:158:HT275DSXX:4:1372:9995:6057 chr3 196164723 N chr3 196164950 N DEL 2
A00404:155:HV27LDSXX:2:2612:15682:6167 chr3 196165158 N chr3 196165280 N DUP 15
A00297:158:HT275DSXX:2:2427:8820:5118 chr3 196165147 N chr3 196165269 N DUP 5
A00297:158:HT275DSXX:2:2664:17861:11694 chr3 196165048 N chr3 196165150 N DEL 1
A00297:158:HT275DSXX:3:2514:11324:24205 chr3 196165151 N chr3 196165273 N DUP 2
A00404:155:HV27LDSXX:3:2631:12029:25113 chr8 82370476 N chr8 82370670 N DUP 5
A00404:155:HV27LDSXX:4:1645:31910:17613 chr8 82370476 N chr8 82370670 N DUP 5
A00404:155:HV27LDSXX:4:1265:31141:19883 chr8 82370476 N chr8 82370670 N DUP 5
A00404:155:HV27LDSXX:4:1543:15890:6151 chr8 82370476 N chr8 82370670 N DUP 5
A00404:156:HV37TDSXX:4:1477:18602:28040 chr8 82370476 N chr8 82370670 N DUP 5
A00404:155:HV27LDSXX:3:2558:14326:33317 chr8 82370476 N chr8 82370670 N DUP 5
A00297:158:HT275DSXX:1:2167:2546:16141 chr8 82370476 N chr8 82370670 N DUP 5
A00404:155:HV27LDSXX:1:1233:28763:27915 chr8 82370476 N chr8 82370670 N DUP 5
A00404:155:HV27LDSXX:2:2404:27968:3865 chr8 82370476 N chr8 82370670 N DUP 5
A00404:156:HV37TDSXX:1:2358:28610:7952 chr8 82370478 N chr8 82370672 N DUP 5
A00404:156:HV37TDSXX:2:1276:1669:5415 chr8 82370483 N chr8 82370677 N DUP 5
A00404:155:HV27LDSXX:2:2662:8838:5337 chr8 82370484 N chr8 82370678 N DUP 5
A00404:156:HV37TDSXX:3:2523:24542:4413 chr8 82370476 N chr8 82370670 N DUP 3
A00404:155:HV27LDSXX:3:2148:22914:35978 chr7 735202 N chr7 735503 N DEL 5
A00297:158:HT275DSXX:1:2325:8567:13886 chr7 735139 N chr7 735440 N DEL 5
A00404:155:HV27LDSXX:3:2148:22914:35978 chr7 735166 N chr7 735596 N DEL 35
A00404:156:HV37TDSXX:2:1447:26838:17628 chr7 735215 N chr7 735372 N DEL 26
A00404:156:HV37TDSXX:4:1216:25138:30029 chr7 735440 N chr7 735709 N DUP 5
A00297:158:HT275DSXX:2:2629:3857:7388 chr12 10526290 N chr12 10526342 N DEL 55
A00297:158:HT275DSXX:3:1514:11749:10191 chr12 10526290 N chr12 10526342 N DEL 56
A00404:155:HV27LDSXX:2:1116:22345:35055 chr12 10526290 N chr12 10526342 N DEL 56
A00297:158:HT275DSXX:2:1460:13838:33786 chr12 10526290 N chr12 10526342 N DEL 56
A00404:155:HV27LDSXX:1:1461:23059:8641 chr12 10526290 N chr12 10526342 N DEL 56
A00404:155:HV27LDSXX:3:1617:11279:27164 chr10 678764 N chr10 678888 N DEL 14
A00404:155:HV27LDSXX:1:1516:8070:11992 chr10 678764 N chr10 678888 N DEL 14
A00404:155:HV27LDSXX:4:2673:28917:11459 chr10 678764 N chr10 678888 N DEL 14
A00404:156:HV37TDSXX:2:1607:7093:34726 chr10 678764 N chr10 678888 N DEL 21
A00404:156:HV37TDSXX:4:2360:16197:3208 chr10 678764 N chr10 678888 N DEL 16
A00297:158:HT275DSXX:2:2130:14353:25097 chr10 678764 N chr10 678888 N DEL 20
A00404:156:HV37TDSXX:4:2352:21441:24846 chr10 679229 N chr10 679416 N DUP 17
A00404:156:HV37TDSXX:4:1676:5520:32095 chr10 679015 N chr10 679482 N DEL 14
A00297:158:HT275DSXX:2:1270:6171:32127 chr10 678953 N chr10 679696 N DUP 16
A00297:158:HT275DSXX:3:1413:4182:32189 chr10 678731 N chr10 679708 N DEL 2
A00404:156:HV37TDSXX:2:2147:29586:19946 chr10 678731 N chr10 679708 N DEL 1
A00297:158:HT275DSXX:2:1550:3215:33990 chr1 213151334 N chr1 213151843 N DEL 10
A00297:158:HT275DSXX:2:2451:31476:30796 chr1 213151334 N chr1 213151843 N DEL 10
A00404:155:HV27LDSXX:3:2547:18430:35790 chr1 213151301 N chr1 213151398 N DUP 12
A00297:158:HT275DSXX:2:2523:15112:30107 chr1 213151296 N chr1 213151393 N DUP 5
A00404:156:HV37TDSXX:2:1175:26069:21872 chr1 213151370 N chr1 213151498 N DEL 5
A00297:158:HT275DSXX:1:1164:18177:23735 chr1 213151424 N chr1 213151552 N DEL 2
A00404:155:HV27LDSXX:2:2245:17219:30906 chr1 213151471 N chr1 213151599 N DEL 5
A00404:155:HV27LDSXX:4:2506:2998:33270 chr1 213151471 N chr1 213151599 N DEL 5
A00404:156:HV37TDSXX:2:2155:18557:26522 chr1 213151359 N chr1 213151485 N DUP 5
A00297:158:HT275DSXX:2:2513:18258:2362 chr1 213151345 N chr1 213151471 N DUP 5
A00297:158:HT275DSXX:4:2310:7500:18991 chr1 213151370 N chr1 213151498 N DEL 10
A00404:155:HV27LDSXX:3:1603:25464:16564 chr1 213151396 N chr1 213151524 N DEL 5
A00404:155:HV27LDSXX:1:2222:26395:3333 chr1 213151578 N chr1 213151833 N DEL 12
A00404:155:HV27LDSXX:4:2277:4182:23015 chr1 213151578 N chr1 213151833 N DEL 18
A00404:155:HV27LDSXX:3:1638:24713:30545 chr1 213151199 N chr1 213151552 N DEL 5
A00297:158:HT275DSXX:1:2246:20247:19492 chr1 213151359 N chr1 213151612 N DUP 10
A00404:156:HV37TDSXX:4:1434:7039:2785 chr1 213151201 N chr1 213151554 N DEL 5
A00404:156:HV37TDSXX:4:1434:7039:2785 chr1 213151205 N chr1 213151558 N DEL 5
A00404:155:HV27LDSXX:4:1369:27082:13135 chr1 213151206 N chr1 213151559 N DEL 5
A00404:155:HV27LDSXX:3:1638:24713:30545 chr1 213151539 N chr1 213151665 N DUP 5
A00404:156:HV37TDSXX:1:2520:19208:29371 chr1 213151539 N chr1 213151665 N DUP 5
A00297:158:HT275DSXX:4:1227:27742:27555 chr1 213151471 N chr1 213151599 N DEL 5
A00297:158:HT275DSXX:4:1227:27796:27993 chr1 213151539 N chr1 213151665 N DUP 5
A00404:155:HV27LDSXX:4:1164:3170:23860 chr1 213151300 N chr1 213151477 N DEL 2
A00404:156:HV37TDSXX:3:2210:29749:1251 chr1 213151358 N chr1 213151613 N DEL 7
A00404:155:HV27LDSXX:3:2125:26395:27665 chr1 213151570 N chr1 213151698 N DEL 5
A00404:156:HV37TDSXX:3:1103:4237:25426 chr1 213151770 N chr1 213152050 N DEL 2
A00404:156:HV37TDSXX:2:1251:23421:20008 chr1 213151469 N chr1 213151771 N DUP 9
A00404:156:HV37TDSXX:3:2236:4390:30577 chr1 213151391 N chr1 213151771 N DUP 5
A00404:156:HV37TDSXX:3:2236:4652:31000 chr1 213151391 N chr1 213151771 N DUP 5
A00297:158:HT275DSXX:3:2355:25482:3693 chr1 213151570 N chr1 213151698 N DEL 5
A00404:155:HV27LDSXX:3:2362:27697:25254 chr1 213151570 N chr1 213151698 N DEL 5
A00297:158:HT275DSXX:3:1301:25192:3912 chr1 213151570 N chr1 213151698 N DEL 5
A00297:158:HT275DSXX:2:1207:27724:6480 chr1 213151570 N chr1 213151698 N DEL 5
A00404:156:HV37TDSXX:4:2240:15429:6950 chr1 213151391 N chr1 213151771 N DUP 8
A00404:155:HV27LDSXX:3:1645:6189:18223 chr1 213151232 N chr1 213151712 N DEL 1
A00404:155:HV27LDSXX:4:2553:21242:14418 chr1 213151232 N chr1 213151712 N DEL 1
A00404:156:HV37TDSXX:4:1624:23647:2644 chr1 213151391 N chr1 213151771 N DUP 10
A00404:155:HV27LDSXX:1:2129:26585:1407 chr1 213151391 N chr1 213151771 N DUP 10
A00404:155:HV27LDSXX:4:1166:29089:15045 chr1 213151391 N chr1 213151771 N DUP 10
A00404:155:HV27LDSXX:4:2277:4300:20619 chr1 213151391 N chr1 213151771 N DUP 10
A00404:156:HV37TDSXX:2:2451:15429:26240 chr1 213151451 N chr1 213151833 N DEL 11
A00404:156:HV37TDSXX:4:2261:7889:24142 chr1 213151407 N chr1 213151789 N DEL 5
A00297:158:HT275DSXX:3:2355:25482:3693 chr1 213151226 N chr1 213151833 N DEL 5
A00404:155:HV27LDSXX:3:1509:27082:18051 chr1 213151228 N chr1 213151835 N DEL 5
A00404:156:HV37TDSXX:3:2236:4390:30577 chr1 213151226 N chr1 213151833 N DEL 5
A00404:156:HV37TDSXX:3:2236:4652:31000 chr1 213151230 N chr1 213151837 N DEL 5
A00404:156:HV37TDSXX:3:2236:4661:30984 chr1 213151226 N chr1 213151833 N DEL 5
A00404:155:HV27LDSXX:4:2277:4182:23015 chr1 213151232 N chr1 213151839 N DEL 5
A00404:156:HV37TDSXX:2:2642:18638:9189 chr1 213151399 N chr1 213151962 N DEL 5
A00297:158:HT275DSXX:3:2603:16676:30843 chr1 213151466 N chr1 213151949 N DUP 13
A00297:158:HT275DSXX:3:1348:27100:22623 chr1 213151263 N chr1 213151971 N DUP 10
A00297:158:HT275DSXX:1:1432:2474:28228 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:1:1633:12680:11522 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:1:2364:30273:21699 chr6 154481281 N chr6 154481553 N DUP 7
A00404:155:HV27LDSXX:3:2609:31177:13933 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:2:1449:4083:18521 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:4:2329:11767:10473 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:3:2260:31250:18192 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:3:2264:32009:16720 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:2:1429:31340:17628 chr6 154481281 N chr6 154481553 N DUP 7
A00404:155:HV27LDSXX:3:1133:26096:15217 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:4:1360:20193:1360 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:4:1618:5104:17848 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:2:1562:29631:7560 chr5 5677737 N chr5 5678187 N DEL 12
A00297:158:HT275DSXX:2:2319:15926:7091 chr5 5677783 N chr5 5677967 N DEL 5
A00404:156:HV37TDSXX:3:2658:4444:14700 chr5 5677847 N chr5 5678031 N DEL 5
A00297:158:HT275DSXX:4:1575:28944:25535 chr5 5677942 N chr5 5678209 N DEL 5
A00404:156:HV37TDSXX:3:2611:13756:9157 chr15 32778286 N chr15 32778341 N DEL 15
A00404:155:HV27LDSXX:3:1259:2989:32095 chr15 32778286 N chr15 32778341 N DEL 12
A00404:156:HV37TDSXX:2:1542:11062:14168 chr9 137380489 N chr9 137380599 N DEL 5
A00297:158:HT275DSXX:2:2401:11180:17785 chr9 137380621 N chr9 137380673 N DUP 10
A00297:158:HT275DSXX:4:2323:22480:16376 chr21 42140468 N chr21 42140559 N DEL 5
A00297:158:HT275DSXX:1:1654:3170:3223 chr21 42140496 N chr21 42140587 N DEL 1
A00297:158:HT275DSXX:3:1656:5394:18349 chr21 42140451 N chr21 42140586 N DUP 5
A00404:155:HV27LDSXX:1:1652:6578:8500 chr21 42140451 N chr21 42140586 N DUP 5
A00297:158:HT275DSXX:1:1654:3170:3223 chr21 42140508 N chr21 42140599 N DEL 13
A00297:158:HT275DSXX:1:1464:12961:21840 chr21 42140481 N chr21 42140572 N DEL 2
A00404:156:HV37TDSXX:4:2410:16740:21527 chr15 48435831 N chr15 48435962 N DEL 5
A00404:155:HV27LDSXX:2:2113:11369:7654 chr8 1330830 N chr8 1330916 N DEL 5
A00297:158:HT275DSXX:2:1611:17083:10191 chr20 62014067 N chr20 62014167 N DUP 10
A00404:156:HV37TDSXX:2:2344:26585:6073 chr20 62014080 N chr20 62014196 N DEL 5
A00404:155:HV27LDSXX:4:2537:26449:20932 chr20 62014069 N chr20 62014203 N DEL 6
A00404:156:HV37TDSXX:2:1175:10140:28197 chr20 62014071 N chr20 62014207 N DEL 4
A00297:158:HT275DSXX:1:2515:21368:27633 chr20 62014071 N chr20 62014209 N DEL 2
A00297:158:HT275DSXX:2:1551:23231:13542 chr20 62014071 N chr20 62014209 N DEL 2
A00297:158:HT275DSXX:3:2168:10700:22968 chr13 112981245 N chr13 112981341 N DEL 11
A00297:158:HT275DSXX:2:2476:11858:5212 chr6 170157785 N chr6 170158533 N DEL 1
A00297:158:HT275DSXX:3:2313:31476:13823 chr6 170157785 N chr6 170158533 N DEL 3
A00297:158:HT275DSXX:3:2313:31720:13620 chr6 170157785 N chr6 170158533 N DEL 3
A00404:155:HV27LDSXX:3:1430:9995:28604 chr6 170157785 N chr6 170158533 N DEL 5
A00297:158:HT275DSXX:3:1113:26594:5368 chr6 170157812 N chr6 170157935 N DEL 3
A00404:156:HV37TDSXX:2:1361:15212:32628 chr6 170157812 N chr6 170157935 N DEL 5
A00297:158:HT275DSXX:2:2668:25012:16689 chr6 170157812 N chr6 170157935 N DEL 6
A00404:155:HV27LDSXX:2:1529:6659:9017 chr6 170157812 N chr6 170157935 N DEL 7
A00404:156:HV37TDSXX:4:2601:14353:2738 chr6 170157812 N chr6 170157935 N DEL 7
A00404:155:HV27LDSXX:4:2215:11360:9298 chr6 170157812 N chr6 170157935 N DEL 7
A00297:158:HT275DSXX:3:1112:9399:34929 chr6 170157842 N chr6 170158215 N DEL 7
A00297:158:HT275DSXX:1:1352:8006:27696 chr6 170157842 N chr6 170158215 N DEL 7
A00297:158:HT275DSXX:2:2644:4237:5509 chr6 170157806 N chr6 170158552 N DUP 10
A00297:158:HT275DSXX:4:2267:16107:23844 chr6 170157898 N chr6 170158190 N DEL 5
A00297:158:HT275DSXX:3:1627:7907:8296 chr6 170157898 N chr6 170158190 N DEL 5
A00297:158:HT275DSXX:4:2231:19226:18129 chr6 170157898 N chr6 170158190 N DEL 5
A00404:156:HV37TDSXX:3:2118:32172:25708 chr6 170157845 N chr6 170157967 N DUP 7
A00404:156:HV37TDSXX:3:2118:32199:25786 chr6 170157845 N chr6 170157967 N DUP 7
A00404:156:HV37TDSXX:3:2609:31485:3850 chr6 170157845 N chr6 170157967 N DUP 7
A00404:155:HV27LDSXX:1:2658:23014:34585 chr6 170157845 N chr6 170157967 N DUP 7
A00404:156:HV37TDSXX:3:1178:17797:33473 chr6 170157845 N chr6 170157967 N DUP 7
A00297:158:HT275DSXX:3:2138:28962:27070 chr6 170157845 N chr6 170157967 N DUP 7
A00297:158:HT275DSXX:3:2313:31476:13823 chr6 170157852 N chr6 170157974 N DUP 7
A00297:158:HT275DSXX:3:2313:31720:13620 chr6 170157852 N chr6 170157974 N DUP 7
A00297:158:HT275DSXX:2:2158:8006:10598 chr6 170157856 N chr6 170157978 N DUP 4
A00297:158:HT275DSXX:2:2158:8386:12164 chr6 170157856 N chr6 170157978 N DUP 4
A00404:155:HV27LDSXX:1:1213:14100:25942 chr6 170157912 N chr6 170158368 N DUP 5
A00404:155:HV27LDSXX:1:1349:6705:3615 chr6 170157912 N chr6 170158368 N DUP 5
A00297:158:HT275DSXX:2:2636:24505:36135 chr6 170157912 N chr6 170158368 N DUP 5
A00404:156:HV37TDSXX:2:2562:20672:8985 chr6 170157912 N chr6 170158035 N DUP 5
A00404:156:HV37TDSXX:4:2563:7093:30906 chr6 170158027 N chr6 170158445 N DEL 8
A00404:156:HV37TDSXX:2:1361:15212:32628 chr6 170158027 N chr6 170158445 N DEL 5
A00404:156:HV37TDSXX:3:2524:13512:36793 chr6 170157968 N chr6 170158258 N DUP 1
A00297:158:HT275DSXX:1:2225:26087:22404 chr6 170158059 N chr6 170158266 N DUP 31
A00297:158:HT275DSXX:2:2668:25012:16689 chr6 170158055 N chr6 170158387 N DUP 5
A00404:155:HV27LDSXX:4:2215:11360:9298 chr6 170158055 N chr6 170158387 N DUP 5
A00297:158:HT275DSXX:3:1627:7907:8296 chr6 170157970 N chr6 170158054 N DEL 5
A00404:156:HV37TDSXX:4:1246:20717:35806 chr6 170158050 N chr6 170158424 N DUP 10
A00297:158:HT275DSXX:2:1338:20455:3129 chr6 170158050 N chr6 170158424 N DUP 10
A00404:156:HV37TDSXX:2:1265:32669:28573 chr6 170157981 N chr6 170158065 N DEL 5
A00297:158:HT275DSXX:4:2557:21206:8876 chr6 170157985 N chr6 170158069 N DEL 5
A00404:156:HV37TDSXX:2:1277:18096:14168 chr6 170157811 N chr6 170158182 N DUP 7
A00404:155:HV27LDSXX:2:2306:24795:20854 chr6 170158134 N chr6 170158299 N DUP 5
A00404:155:HV27LDSXX:3:2172:8549:32612 chr6 170158147 N chr6 170158229 N DUP 4
A00404:155:HV27LDSXX:3:1446:10393:23688 chr6 170158286 N chr6 170158580 N DEL 5
A00404:156:HV37TDSXX:4:2325:17354:6934 chr6 170157975 N chr6 170158059 N DEL 6
A00404:155:HV27LDSXX:4:2456:4869:20259 chr6 170157955 N chr6 170158414 N DEL 9
A00404:156:HV37TDSXX:2:1644:13720:9752 chr6 170157975 N chr6 170158059 N DEL 5
A00404:155:HV27LDSXX:1:1213:14100:25942 chr6 170157975 N chr6 170158059 N DEL 13
A00297:158:HT275DSXX:1:1474:12771:19038 chr6 170158349 N chr6 170158643 N DEL 13
A00297:158:HT275DSXX:3:1462:31873:18991 chr6 170158360 N chr6 170158445 N DEL 3
A00404:155:HV27LDSXX:1:2362:2935:35289 chr6 170158360 N chr6 170158445 N DEL 5
A00404:155:HV27LDSXX:3:1312:23267:8656 chr6 170158360 N chr6 170158445 N DEL 5
A00297:158:HT275DSXX:2:1237:24795:30624 chr6 170158329 N chr6 170158621 N DUP 5
A00404:156:HV37TDSXX:3:1130:3730:14309 chr6 170158320 N chr6 170158612 N DUP 5
A00297:158:HT275DSXX:4:1474:4770:6872 chr6 170158153 N chr6 170158320 N DEL 5
A00404:155:HV27LDSXX:1:1668:10339:11350 chr6 170158115 N chr6 170158407 N DEL 17
A00297:158:HT275DSXX:3:2232:15899:29966 chr6 170158383 N chr6 170158466 N DUP 5
A00297:158:HT275DSXX:3:2232:15908:29919 chr6 170158383 N chr6 170158466 N DUP 5
A00404:155:HV27LDSXX:2:2306:24795:20854 chr6 170157973 N chr6 170158390 N DEL 5
A00404:155:HV27LDSXX:1:1668:10339:11350 chr6 170157995 N chr6 170158412 N DEL 5
A00404:155:HV27LDSXX:1:2362:2935:35289 chr6 170158423 N chr6 170158550 N DEL 5
A00297:158:HT275DSXX:1:2339:26214:14231 chr7 60911830 N chr7 60912015 N DUP 3
A00404:155:HV27LDSXX:1:1514:15374:17660 chr7 60911855 N chr7 60912042 N DEL 5
A00404:155:HV27LDSXX:3:1151:14895:18865 chr4 19226462 N chr4 19226547 N DEL 30
A00297:158:HT275DSXX:2:2160:23547:8234 chr4 19226439 N chr4 19226547 N DEL 25
A00404:156:HV37TDSXX:3:2171:5810:14434 chr4 19226416 N chr4 19226547 N DEL 16
A00404:155:HV27LDSXX:2:2248:24876:35149 chr4 19226691 N chr4 19226744 N DEL 2
A00297:158:HT275DSXX:4:1405:27444:29387 chr6 165749331 N chr6 165749567 N DEL 13
A00404:155:HV27LDSXX:3:1628:16432:19304 chr6 165749331 N chr6 165749435 N DEL 15
A00404:156:HV37TDSXX:1:1257:20157:14481 chr6 165749331 N chr6 165749435 N DEL 17
A00404:156:HV37TDSXX:2:1271:16740:7467 chr6 165749331 N chr6 165749435 N DEL 19
A00297:158:HT275DSXX:1:1350:3685:12414 chr6 165749331 N chr6 165749435 N DEL 20
A00404:155:HV27LDSXX:2:2113:7898:2425 chr6 165749331 N chr6 165749435 N DEL 22
A00404:156:HV37TDSXX:3:1464:9290:14700 chr6 165749331 N chr6 165749435 N DEL 32
A00404:156:HV37TDSXX:1:2515:22345:7905 chr6 165749334 N chr6 165749508 N DUP 10
A00404:156:HV37TDSXX:3:1277:13096:12242 chr6 165749334 N chr6 165749508 N DUP 9
A00404:155:HV27LDSXX:4:1456:13006:7764 chr6 165749334 N chr6 165749508 N DUP 8
A00404:156:HV37TDSXX:4:1176:6768:23328 chr6 165749556 N chr6 165749625 N DEL 5
A00297:158:HT275DSXX:2:2578:20229:31704 chr6 165749392 N chr6 165749482 N DEL 10
A00404:155:HV27LDSXX:3:1420:25102:14998 chr6 165749476 N chr6 165749564 N DEL 16
A00404:155:HV27LDSXX:4:1244:12138:32878 chr6 165749474 N chr6 165749562 N DEL 25
A00404:155:HV27LDSXX:3:1118:13557:21026 chr6 165749418 N chr6 165749506 N DEL 13
A00404:156:HV37TDSXX:1:1170:1353:31109 chr6 165749418 N chr6 165749506 N DEL 12
A00404:156:HV37TDSXX:1:1539:11822:2769 chr6 165749447 N chr6 165749565 N DEL 21
A00297:158:HT275DSXX:4:1665:3658:33724 chr6 165749405 N chr6 165749639 N DEL 4
A00404:156:HV37TDSXX:2:1362:17680:17331 chr7 17112872 N chr7 17113102 N DUP 9
A00404:155:HV27LDSXX:4:1175:3179:21496 chr14 19023367 N chr14 19023516 N DEL 7
A00297:158:HT275DSXX:2:1304:9019:11193 chr5 33626707 N chr5 33626795 N DUP 2
A00297:158:HT275DSXX:4:1272:29161:19147 chr5 33626707 N chr5 33626795 N DUP 3
A00404:156:HV37TDSXX:1:2104:32497:29778 chr5 33626707 N chr5 33626795 N DUP 3
A00404:156:HV37TDSXX:2:1224:29188:1783 chr16 46414835 N chr16 46414977 N DUP 2
A00404:156:HV37TDSXX:4:2537:14570:5807 chrX 647735 N chrX 648472 N DUP 5
A00404:156:HV37TDSXX:2:1639:8784:5149 chrX 647432 N chrX 648417 N DEL 5
A00404:155:HV27LDSXX:3:2669:10230:36182 chrX 647650 N chrX 648469 N DUP 5
A00404:155:HV27LDSXX:4:2450:4426:17018 chrX 647678 N chrX 648417 N DEL 5
A00404:156:HV37TDSXX:2:2534:14868:5509 chrX 647650 N chrX 648469 N DUP 5
A00404:156:HV37TDSXX:4:2537:14751:6245 chrX 647653 N chrX 648472 N DUP 5
A00404:156:HV37TDSXX:4:1414:18313:33552 chrX 647412 N chrX 648397 N DEL 5
A00404:155:HV27LDSXX:3:1560:2998:12383 chrX 647671 N chrX 648328 N DEL 5
A00404:155:HV27LDSXX:4:2510:21549:11381 chrX 647671 N chrX 648328 N DEL 5
A00404:156:HV37TDSXX:1:1525:11532:2769 chrX 647412 N chrX 648397 N DEL 5
A00404:155:HV27LDSXX:4:1607:16776:15264 chrX 647732 N chrX 648469 N DUP 5
A00404:156:HV37TDSXX:4:2537:14570:5807 chrX 647404 N chrX 648469 N DUP 5
A00404:156:HV37TDSXX:4:2537:14751:6245 chrX 647404 N chrX 648469 N DUP 5
A00404:155:HV27LDSXX:1:2564:1551:9565 chrX 647404 N chrX 648469 N DUP 5
A00404:156:HV37TDSXX:4:1350:18023:28447 chrX 648159 N chrX 648486 N DUP 5
A00297:158:HT275DSXX:2:1315:25997:5149 chrX 648306 N chrX 648469 N DUP 5
A00297:158:HT275DSXX:4:2526:16378:6089 chrX 647671 N chrX 648328 N DEL 5
A00404:155:HV27LDSXX:1:1111:24731:36902 chrX 647671 N chrX 648328 N DEL 5
A00404:155:HV27LDSXX:3:1560:2998:12383 chrX 647671 N chrX 648328 N DEL 5
A00404:155:HV27LDSXX:1:2542:25373:29183 chrX 647674 N chrX 648331 N DEL 5
A00404:156:HV37TDSXX:4:1350:18023:28447 chrX 647685 N chrX 648342 N DEL 1
A00404:156:HV37TDSXX:1:1260:30689:4413 chrX 648305 N chrX 648470 N DEL 5
A00404:156:HV37TDSXX:3:1229:18945:27915 chrX 647403 N chrX 648470 N DEL 8
A00404:156:HV37TDSXX:3:1229:18945:27915 chrX 647403 N chrX 648470 N DEL 5
A00404:155:HV27LDSXX:2:2659:9851:23844 chr16 55023161 N chr16 55023225 N DUP 17
A00404:156:HV37TDSXX:3:2341:24008:8093 chr16 55023161 N chr16 55023225 N DUP 16
A00404:155:HV27LDSXX:1:1354:17544:34976 chr16 55023165 N chr16 55023229 N DUP 11
A00404:156:HV37TDSXX:1:1547:29360:6965 chr1 222689644 N chr1 222689731 N DEL 3
A00404:156:HV37TDSXX:1:1547:32841:7513 chr1 222689644 N chr1 222689731 N DEL 3
A00297:158:HT275DSXX:1:1316:24505:32878 chr16 85346346 N chr16 85346447 N DEL 10
A00404:155:HV27LDSXX:3:2118:30101:36714 chr16 85346573 N chr16 85346847 N DEL 12
A00404:155:HV27LDSXX:3:1355:31204:11631 chr16 85346573 N chr16 85346847 N DEL 13
A00404:156:HV37TDSXX:4:1550:32199:14168 chr16 85346594 N chr16 85346870 N DUP 1
A00404:155:HV27LDSXX:1:2353:26955:20337 chr16 85346502 N chr16 85346590 N DEL 5
A00404:156:HV37TDSXX:1:2528:27163:29340 chr16 85346270 N chr16 85346764 N DEL 7
A00404:155:HV27LDSXX:3:1639:6795:25347 chr18 9886993 N chr18 9887397 N DUP 5
A00404:156:HV37TDSXX:4:2655:11704:14497 chr18 9887070 N chr18 9887386 N DEL 5
A00404:156:HV37TDSXX:3:2654:14796:13745 chr18 9887121 N chr18 9887302 N DEL 2
A00297:158:HT275DSXX:3:2369:25337:28056 chr18 9887121 N chr18 9887302 N DEL 20
A00404:156:HV37TDSXX:2:1118:29297:35947 chr18 9887243 N chr18 9887604 N DEL 13
A00404:156:HV37TDSXX:2:1129:13304:17769 chr18 9887046 N chr18 9887227 N DEL 8
A00297:158:HT275DSXX:1:1237:26756:24283 chr18 9887028 N chr18 9887344 N DEL 30
A00404:156:HV37TDSXX:2:2458:22670:11130 chr18 9887127 N chr18 9887308 N DEL 12
A00404:156:HV37TDSXX:2:2312:32570:15687 chr18 9887248 N chr18 9887384 N DEL 4
A00404:156:HV37TDSXX:4:2655:11704:14497 chr18 9887070 N chr18 9887386 N DEL 15
A00297:158:HT275DSXX:2:2227:29234:4398 chr18 9887093 N chr18 9887409 N DEL 16
A00297:158:HT275DSXX:2:1117:32244:31814 chr18 9887458 N chr18 9887549 N DEL 5
A00297:158:HT275DSXX:2:2227:29234:4398 chr18 9887093 N chr18 9887409 N DEL 5
A00404:156:HV37TDSXX:3:2107:4878:17112 chr18 9887172 N chr18 9887488 N DEL 10
A00404:155:HV27LDSXX:1:2206:12897:6073 chr18 9887524 N chr18 9887613 N DUP 5
A00297:158:HT275DSXX:4:1556:19090:15859 chr18 9887523 N chr18 9887614 N DEL 5
A00297:158:HT275DSXX:4:2161:11948:9784 chr18 9887265 N chr18 9887671 N DEL 31
A00297:158:HT275DSXX:4:2161:11948:9784 chr18 9887265 N chr18 9887671 N DEL 21
A00404:155:HV27LDSXX:2:2609:20889:18349 chr18 9887550 N chr18 9887686 N DEL 9
A00297:158:HT275DSXX:2:1401:11496:18082 chr18 9887238 N chr18 9887779 N DEL 3
A00297:158:HT275DSXX:4:1169:10429:20744 chr18 9887589 N chr18 9887860 N DEL 12
A00297:158:HT275DSXX:1:2455:19777:21621 chr20 14955047 N chr20 14955191 N DEL 3
A00297:158:HT275DSXX:2:1208:19633:1172 chr2 146697005 N chr2 146697072 N DEL 5
A00404:155:HV27LDSXX:2:1359:30029:16705 chr2 146697005 N chr2 146697072 N DEL 5
A00404:156:HV37TDSXX:2:2620:27950:19930 chr13 34540649 N chr13 34540845 N DUP 5
A00404:155:HV27LDSXX:3:2633:29089:16799 chr13 34540945 N chr13 34540994 N DUP 10
A00404:155:HV27LDSXX:2:2447:24243:27289 chr13 34540945 N chr13 34540994 N DUP 12
A00404:155:HV27LDSXX:3:1463:18819:13479 chr13 34541009 N chr13 34541286 N DEL 5
A00297:158:HT275DSXX:1:2530:29071:3552 chr13 34541009 N chr13 34541286 N DEL 11
A00297:158:HT275DSXX:4:2641:25156:23234 chr13 34541009 N chr13 34541286 N DEL 11
A00404:155:HV27LDSXX:2:1259:1859:19836 chr13 34541009 N chr13 34541286 N DEL 11
A00404:155:HV27LDSXX:1:2252:26187:4883 chr13 34541009 N chr13 34541286 N DEL 11
A00404:155:HV27LDSXX:2:1578:4399:24330 chr13 34541046 N chr13 34541321 N DUP 5
A00297:158:HT275DSXX:4:2150:18403:23312 chr13 34540906 N chr13 34541004 N DEL 7
A00404:155:HV27LDSXX:4:2631:9941:31579 chr13 34541054 N chr13 34541506 N DUP 12
A00404:155:HV27LDSXX:1:2131:14832:32471 chr13 34540917 N chr13 34541016 N DEL 5
A00404:155:HV27LDSXX:1:1311:31024:24283 chr13 34541151 N chr13 34541200 N DUP 6
A00404:156:HV37TDSXX:1:2343:17544:32033 chr13 34541226 N chr13 34541504 N DEL 12
A00404:155:HV27LDSXX:1:1616:3830:12038 chr13 34541156 N chr13 34541430 N DUP 5
A00297:158:HT275DSXX:3:2158:18665:31939 chr13 34541151 N chr13 34541200 N DUP 18
A00404:155:HV27LDSXX:1:2252:26187:4883 chr13 34541075 N chr13 34541154 N DEL 9
A00297:158:HT275DSXX:1:1254:10013:11287 chr13 34541156 N chr13 34541205 N DUP 10
A00404:155:HV27LDSXX:3:1303:22670:21245 chr13 34541156 N chr13 34541205 N DUP 10
A00404:155:HV27LDSXX:1:1138:14796:1658 chr13 34541172 N chr13 34541270 N DUP 11
A00404:156:HV37TDSXX:4:2445:15845:30185 chr13 34541263 N chr13 34541441 N DEL 10
A00404:155:HV27LDSXX:3:1229:20781:22420 chr13 34541330 N chr13 34541511 N DEL 9
A00404:156:HV37TDSXX:1:1504:10194:4085 chr13 34540918 N chr13 34541244 N DEL 5
A00404:156:HV37TDSXX:2:1577:20464:26757 chr13 34541009 N chr13 34541286 N DEL 5
A00404:155:HV27LDSXX:4:1553:30165:22639 chr13 34541406 N chr13 34541509 N DEL 3
A00404:155:HV27LDSXX:4:2563:9480:10426 chr13 34541425 N chr13 34541476 N DEL 9
A00404:156:HV37TDSXX:1:1136:14443:28823 chr13 34541425 N chr13 34541476 N DEL 10
A00297:158:HT275DSXX:2:2175:31006:14387 chr13 34541425 N chr13 34541476 N DEL 13
A00404:155:HV27LDSXX:3:2620:31891:8155 chr13 34541010 N chr13 34541464 N DEL 11
A00297:158:HT275DSXX:4:2232:17020:30624 chr13 34541430 N chr13 34541481 N DEL 5
A00404:155:HV27LDSXX:4:1654:1362:25989 chr13 34541430 N chr13 34541481 N DEL 5
A00404:155:HV27LDSXX:4:1654:2510:12007 chr13 34541430 N chr13 34541481 N DEL 5
A00297:158:HT275DSXX:2:1406:25183:19116 chr13 34541356 N chr13 34541537 N DEL 13
A00404:155:HV27LDSXX:3:1303:22670:21245 chr13 34541025 N chr13 34541531 N DEL 5
A00404:156:HV37TDSXX:4:1428:15664:16407 chr13 34541026 N chr13 34541532 N DEL 5
A00404:156:HV37TDSXX:4:1428:16016:15953 chr13 34541026 N chr13 34541532 N DEL 5
A00404:156:HV37TDSXX:2:1348:31304:16971 chr13 34541028 N chr13 34541534 N DEL 5
A00404:155:HV27LDSXX:1:1335:10755:10504 chr19 32058451 N chr19 32058553 N DEL 4
A00297:158:HT275DSXX:4:2457:14633:28119 chr5 131579821 N chr5 131579900 N DEL 4
A00404:156:HV37TDSXX:4:2676:7943:20885 chr15 26893285 N chr15 26893539 N DEL 5
A00404:155:HV27LDSXX:4:1636:4824:11412 chr15 26893346 N chr15 26893400 N DEL 5
A00404:155:HV27LDSXX:4:1218:23059:3129 chr15 26893346 N chr15 26893400 N DEL 5
A00404:155:HV27LDSXX:3:2516:22209:9799 chr15 26893404 N chr15 26893496 N DEL 5
A00297:158:HT275DSXX:3:2671:7003:6261 chr15 26893356 N chr15 26893557 N DUP 5
A00404:155:HV27LDSXX:2:2323:28565:8750 chr9 35913696 N chr9 35914153 N DEL 7
A00404:156:HV37TDSXX:4:2145:24994:21010 chr9 35913676 N chr9 35913777 N DUP 25
A00404:155:HV27LDSXX:2:1418:17011:33051 chr9 35913697 N chr9 35914522 N DUP 10
A00404:155:HV27LDSXX:2:2430:10447:11694 chr9 35913670 N chr9 35914391 N DUP 12
A00404:155:HV27LDSXX:2:1565:28637:2018 chr9 35913730 N chr9 35914555 N DUP 15
A00404:156:HV37TDSXX:3:1368:7428:21621 chr9 35913714 N chr9 35913767 N DUP 5
A00404:155:HV27LDSXX:4:2172:6488:33082 chr9 35913762 N chr9 35914385 N DEL 15
A00404:156:HV37TDSXX:4:2104:23791:30358 chr9 35913775 N chr9 35914500 N DEL 15
A00404:156:HV37TDSXX:4:2664:28483:2503 chr9 35913764 N chr9 35913965 N DUP 5
A00404:155:HV27LDSXX:4:1231:5864:19382 chr9 35913778 N chr9 35914347 N DEL 17
A00404:156:HV37TDSXX:1:1232:23457:28902 chr9 35913777 N chr9 35914346 N DEL 20
A00297:158:HT275DSXX:3:2569:9688:23437 chr9 35913784 N chr9 35914139 N DEL 17
A00297:158:HT275DSXX:3:2569:9688:23437 chr9 35913809 N chr9 35914484 N DEL 8
A00404:156:HV37TDSXX:1:1412:28167:22811 chr9 35913848 N chr9 35914469 N DEL 5
A00404:155:HV27LDSXX:2:2276:1506:11271 chr9 35913655 N chr9 35914068 N DEL 5
A00404:155:HV27LDSXX:3:2313:8504:20509 chr9 35913658 N chr9 35914065 N DEL 13
A00404:156:HV37TDSXX:1:1374:12066:6918 chr9 35913774 N chr9 35914079 N DEL 8
A00297:158:HT275DSXX:2:2347:1940:6324 chr9 35913799 N chr9 35914420 N DUP 8
A00404:155:HV27LDSXX:2:1309:22444:28494 chr9 35913799 N chr9 35914420 N DUP 5
A00297:158:HT275DSXX:1:2369:20772:23688 chr9 35913784 N chr9 35913835 N DEL 22
A00404:156:HV37TDSXX:4:2366:7925:22294 chr9 35913835 N chr9 35913938 N DUP 5
A00297:158:HT275DSXX:2:2347:1940:6324 chr9 35913835 N chr9 35914038 N DUP 10
A00404:155:HV27LDSXX:3:2169:31819:17926 chr9 35913835 N chr9 35913938 N DUP 5
A00404:156:HV37TDSXX:3:1339:8061:4460 chr9 35913919 N chr9 35914436 N DUP 16
A00404:156:HV37TDSXX:4:2274:32796:36808 chr9 35913964 N chr9 35914435 N DUP 15
A00297:158:HT275DSXX:3:1608:4526:13401 chr9 35913730 N chr9 35914555 N DUP 15
A00297:158:HT275DSXX:4:1262:3766:10739 chr9 35914217 N chr9 35914382 N DEL 10
A00404:155:HV27LDSXX:3:2142:9896:21637 chr9 35914346 N chr9 35914555 N DUP 11
A00404:156:HV37TDSXX:1:1421:29857:21198 chr9 35914346 N chr9 35914555 N DUP 15
A00404:155:HV27LDSXX:3:2377:17635:24987 chr9 35914217 N chr9 35914484 N DEL 15
A00404:155:HV27LDSXX:3:2234:21486:34225 chr9 35913914 N chr9 35914221 N DUP 10
A00404:155:HV27LDSXX:1:1524:12924:18521 chr9 35914217 N chr9 35914484 N DEL 17
A00404:155:HV27LDSXX:1:1524:16758:16360 chr9 35914217 N chr9 35914484 N DEL 17
A00297:158:HT275DSXX:4:2565:11125:15280 chr9 35913914 N chr9 35914221 N DUP 8
A00297:158:HT275DSXX:1:1362:5936:25739 chr9 35913914 N chr9 35914435 N DUP 19
A00404:155:HV27LDSXX:3:2142:9896:21637 chr9 35913863 N chr9 35913914 N DEL 5
A00404:155:HV27LDSXX:3:2656:21314:15890 chr9 35913863 N chr9 35913914 N DEL 5
A00404:155:HV27LDSXX:4:2657:1298:9220 chr9 35914206 N chr9 35914469 N DEL 14
A00404:155:HV27LDSXX:4:2547:16523:35493 chr9 35913863 N chr9 35913914 N DEL 7
A00404:155:HV27LDSXX:2:1418:17011:33051 chr9 35913863 N chr9 35913914 N DEL 10
A00404:155:HV27LDSXX:1:2370:22761:14794 chr9 35914271 N chr9 35914384 N DEL 4
A00404:156:HV37TDSXX:3:1514:15492:25066 chr9 35913964 N chr9 35914275 N DEL 5
A00297:158:HT275DSXX:2:2417:28736:26584 chr9 35913690 N chr9 35913997 N DEL 5
A00297:158:HT275DSXX:3:2453:8458:35430 chr9 35913694 N chr9 35914001 N DEL 3
A00297:158:HT275DSXX:1:2344:11035:27179 chr9 35914013 N chr9 35914382 N DEL 1
A00404:155:HV27LDSXX:2:1232:2799:31015 chr9 35913938 N chr9 35913989 N DEL 5
A00297:158:HT275DSXX:2:1156:22516:10645 chr9 35913938 N chr9 35913989 N DEL 1
A00404:155:HV27LDSXX:2:2555:9598:36902 chr9 35913784 N chr9 35913835 N DEL 23
A00404:155:HV27LDSXX:4:1625:29243:12273 chr9 35913938 N chr9 35913989 N DEL 5
A00404:155:HV27LDSXX:2:1144:4020:35540 chr9 35913989 N chr9 35914038 N DUP 7
A00404:155:HV27LDSXX:3:1560:16315:20447 chr9 35913989 N chr9 35914406 N DUP 20
A00297:158:HT275DSXX:4:1530:21395:28087 chr9 35913989 N chr9 35914406 N DUP 8
A00404:155:HV27LDSXX:2:1144:4020:35540 chr9 35914032 N chr9 35914187 N DEL 4
A00404:156:HV37TDSXX:1:2263:20781:20760 chr9 35914328 N chr9 35914431 N DUP 6
A00404:155:HV27LDSXX:3:1102:30337:36057 chr9 35914382 N chr9 35914431 N DUP 13
A00404:155:HV27LDSXX:4:2151:10257:29434 chr9 35913938 N chr9 35913989 N DEL 5
A00404:155:HV27LDSXX:2:1224:21414:14841 chr9 35913940 N chr9 35913991 N DEL 5
A00404:155:HV27LDSXX:1:2370:22761:14794 chr9 35913943 N chr9 35913994 N DEL 5
A00404:155:HV27LDSXX:1:2476:4318:5932 chr9 35913989 N chr9 35914038 N DUP 10
A00404:156:HV37TDSXX:4:2330:25446:36260 chr9 35913989 N chr9 35914038 N DUP 10
A00404:155:HV27LDSXX:4:2657:1298:9220 chr9 35914331 N chr9 35914536 N DUP 11
A00404:156:HV37TDSXX:4:2274:32796:36808 chr9 35913938 N chr9 35913989 N DEL 5
A00404:156:HV37TDSXX:1:2436:4472:16250 chr9 35913967 N chr9 35914114 N DUP 10
A00404:156:HV37TDSXX:4:1315:4734:15389 chr9 35913914 N chr9 35914435 N DUP 10
A00404:155:HV27LDSXX:2:2306:8892:35712 chr9 35914063 N chr9 35914484 N DEL 10
A00297:158:HT275DSXX:2:2563:16378:10097 chr9 35914113 N chr9 35914222 N DEL 12
A00297:158:HT275DSXX:2:2257:17463:31673 chr9 35914113 N chr9 35914222 N DEL 12
A00404:155:HV27LDSXX:3:1102:30337:36057 chr9 35914053 N chr9 35914206 N DUP 5
A00404:156:HV37TDSXX:4:2101:16893:9204 chr9 35914221 N chr9 35914488 N DEL 10
A00404:156:HV37TDSXX:4:2105:10456:16000 chr9 35914431 N chr9 35914484 N DEL 6
A00297:158:HT275DSXX:1:2630:2953:3505 chr9 35913913 N chr9 35914016 N DUP 10
A00404:155:HV27LDSXX:1:2521:19614:17049 chr9 35913708 N chr9 35913813 N DEL 10
A00297:158:HT275DSXX:1:2344:11035:27179 chr9 35913981 N chr9 35914346 N DEL 5
A00297:158:HT275DSXX:3:1524:8983:12383 chr9 35913708 N chr9 35914117 N DEL 10
A00297:158:HT275DSXX:3:2605:5113:12007 chr9 35914103 N chr9 35914420 N DUP 5
A00404:155:HV27LDSXX:4:2159:14579:11898 chr9 35914103 N chr9 35914420 N DUP 5
A00297:158:HT275DSXX:3:2453:8458:35430 chr9 35914103 N chr9 35914420 N DUP 5
A00404:155:HV27LDSXX:3:2313:8504:20509 chr9 35914103 N chr9 35914420 N DUP 7
A00404:155:HV27LDSXX:2:1232:2799:31015 chr9 35914103 N chr9 35914420 N DUP 5
A00297:158:HT275DSXX:1:1272:28357:26866 chr9 35914328 N chr9 35914431 N DUP 8
A00404:155:HV27LDSXX:2:2675:19334:28839 chr9 35913799 N chr9 35914420 N DUP 5
A00404:155:HV27LDSXX:4:1232:15718:33974 chr9 35914185 N chr9 35914502 N DEL 2
A00404:156:HV37TDSXX:1:2526:14778:4288 chr9 35913914 N chr9 35914435 N DUP 6
A00404:156:HV37TDSXX:1:2436:4472:16250 chr9 35913707 N chr9 35913812 N DEL 7
A00404:156:HV37TDSXX:1:2263:20781:20760 chr9 35914057 N chr9 35914474 N DEL 19
A00404:155:HV27LDSXX:2:2428:16098:17816 chr9 35913916 N chr9 35914223 N DUP 14
A00404:156:HV37TDSXX:2:2209:13367:12837 chr9 35913939 N chr9 35914456 N DEL 16
A00404:155:HV27LDSXX:2:1565:28637:2018 chr9 35914206 N chr9 35914469 N DEL 14
A00404:155:HV27LDSXX:2:2542:22941:33959 chr9 35913914 N chr9 35914435 N DUP 19
A00297:158:HT275DSXX:4:2529:11505:10770 chr9 35913914 N chr9 35914435 N DUP 14
A00404:156:HV37TDSXX:4:1315:4734:15389 chr9 35914206 N chr9 35914469 N DEL 19
A00404:155:HV27LDSXX:3:2234:21486:34225 chr9 35914217 N chr9 35914484 N DEL 17
A00404:155:HV27LDSXX:2:1533:24740:17347 chr9 35914217 N chr9 35914484 N DEL 17
A00404:155:HV27LDSXX:2:1237:5104:16094 chr9 35914215 N chr9 35914478 N DEL 19
A00297:158:HT275DSXX:4:1564:32542:36025 chr9 35913863 N chr9 35914064 N DEL 10
A00404:156:HV37TDSXX:1:1454:26829:28917 chr9 35913962 N chr9 35914479 N DEL 8
A00404:155:HV27LDSXX:4:1121:6397:27978 chr9 35913775 N chr9 35914236 N DEL 19
A00297:158:HT275DSXX:3:2605:5113:12007 chr9 35914346 N chr9 35914555 N DUP 15
A00404:156:HV37TDSXX:2:1360:12210:2127 chr9 35913676 N chr9 35914291 N DUP 10
A00404:156:HV37TDSXX:1:1527:21088:11741 chr9 35913634 N chr9 35913789 N DUP 9
A00297:158:HT275DSXX:1:2277:25626:23766 chr9 35913829 N chr9 35914265 N DEL 5
A00297:158:HT275DSXX:4:1646:1488:35916 chr9 35913938 N chr9 35914299 N DEL 14
A00297:158:HT275DSXX:4:2215:16504:36839 chr9 35913682 N chr9 35914299 N DEL 10
A00297:158:HT275DSXX:4:2215:16504:36839 chr9 35913675 N chr9 35914292 N DEL 5
A00297:158:HT275DSXX:3:2544:2591:22294 chr9 35913938 N chr9 35914299 N DEL 14
A00404:155:HV27LDSXX:1:2455:5963:6183 chr9 35913621 N chr9 35914292 N DEL 5
A00297:158:HT275DSXX:3:2544:2591:22294 chr9 35913968 N chr9 35914329 N DEL 15
A00404:155:HV27LDSXX:3:1329:4300:32268 chr9 35914346 N chr9 35914555 N DUP 15
A00404:155:HV27LDSXX:4:1257:6533:16000 chr9 35914346 N chr9 35914555 N DUP 15
A00404:155:HV27LDSXX:4:1258:8133:4711 chr9 35914346 N chr9 35914555 N DUP 15
A00404:156:HV37TDSXX:1:2440:14181:12148 chr9 35914346 N chr9 35914555 N DUP 15
A00297:158:HT275DSXX:4:1340:26838:32753 chr9 35914217 N chr9 35914382 N DEL 10
A00404:155:HV27LDSXX:4:2128:20202:17973 chr9 35914064 N chr9 35914435 N DUP 11
A00297:158:HT275DSXX:3:2302:20808:16391 chr9 35914064 N chr9 35914435 N DUP 14
A00297:158:HT275DSXX:3:1514:25644:29309 chr9 35913914 N chr9 35914221 N DUP 9
A00297:158:HT275DSXX:2:1166:1931:25629 chr9 35913989 N chr9 35914406 N DUP 5
A00297:158:HT275DSXX:2:2563:16378:10097 chr9 35913762 N chr9 35913917 N DEL 10
A00297:158:HT275DSXX:4:1646:1488:35916 chr9 35913989 N chr9 35914406 N DUP 19
A00404:156:HV37TDSXX:1:2303:25337:20729 chr9 35914379 N chr9 35914534 N DUP 10
A00404:155:HV27LDSXX:1:1438:26892:18944 chr9 35914379 N chr9 35914432 N DUP 10
A00297:158:HT275DSXX:4:1622:23258:27743 chr9 35914379 N chr9 35914432 N DUP 10
A00404:155:HV27LDSXX:3:2229:1750:7247 chr9 35914379 N chr9 35914432 N DUP 8
A00404:156:HV37TDSXX:1:2469:3378:29857 chr9 35913767 N chr9 35914384 N DEL 5
A00404:156:HV37TDSXX:4:1552:6768:20572 chr9 35914218 N chr9 35914379 N DEL 5
A00297:158:HT275DSXX:4:1262:3766:10739 chr9 35914218 N chr9 35914379 N DEL 5
A00404:156:HV37TDSXX:4:2175:5077:29575 chr9 35914431 N chr9 35914484 N DEL 22
A00404:155:HV27LDSXX:1:1405:21350:31516 chr9 35914217 N chr9 35914484 N DEL 17
A00404:156:HV37TDSXX:4:2455:21251:16877 chr9 35914217 N chr9 35914484 N DEL 17
A00297:158:HT275DSXX:4:1564:32542:36025 chr9 35914217 N chr9 35914484 N DEL 17
A00404:155:HV27LDSXX:3:2509:12084:9017 chr9 35913658 N chr9 35914383 N DEL 4
A00297:158:HT275DSXX:3:1359:10592:2425 chr9 35914484 N chr9 35914533 N DUP 22
A00404:155:HV27LDSXX:3:2113:2618:4178 chr9 35914328 N chr9 35914431 N DUP 7
A00404:155:HV27LDSXX:3:2113:3034:2863 chr9 35914328 N chr9 35914431 N DUP 7
A00404:155:HV27LDSXX:1:2219:25238:10473 chr9 35913999 N chr9 35914518 N DUP 8
A00297:158:HT275DSXX:1:2616:30228:17425 chr9 35914469 N chr9 35914522 N DUP 4
A00297:158:HT275DSXX:1:1158:25256:11819 chr9 35914206 N chr9 35914469 N DEL 14
A00404:156:HV37TDSXX:1:1454:26829:28917 chr9 35914469 N chr9 35914522 N DUP 20
A00404:156:HV37TDSXX:3:2661:9616:32174 chr9 35914508 N chr9 35914563 N DEL 5
A00404:156:HV37TDSXX:3:2126:5556:34100 chr9 35914406 N chr9 35914563 N DEL 5
A00404:156:HV37TDSXX:3:2135:19361:25003 chr9 35913938 N chr9 35914563 N DEL 5
A00404:156:HV37TDSXX:2:2403:20103:18082 chr7 61286934 N chr7 61287423 N DUP 10
A00297:158:HT275DSXX:2:2412:18683:2409 chr4 188755236 N chr4 188755438 N DEL 24
A00297:158:HT275DSXX:1:1618:13765:26647 chr2 89264431 N chr2 89264589 N DEL 3
A00404:155:HV27LDSXX:4:1109:8847:8609 chr2 89264467 N chr2 89264568 N DEL 30
A00404:156:HV37TDSXX:4:2356:2862:8609 chr2 89264467 N chr2 89264568 N DEL 15
A00297:158:HT275DSXX:4:2436:28809:5729 chr2 89264493 N chr2 89264566 N DUP 12
A00404:156:HV37TDSXX:1:2369:14778:28056 chr2 89264482 N chr2 89264535 N DEL 7
A00404:155:HV27LDSXX:3:1233:1344:27680 chr2 89264490 N chr2 89264543 N DEL 9
A00404:155:HV27LDSXX:4:2656:14326:10895 chr2 89264467 N chr2 89264544 N DEL 7
A00297:158:HT275DSXX:1:2533:23981:29496 chr2 89264544 N chr2 89264610 N DUP 12
A00404:156:HV37TDSXX:4:1410:2401:3082 chr2 89264508 N chr2 89264746 N DUP 2
A00404:156:HV37TDSXX:4:1338:12979:26663 chr10 70999618 N chr10 70999689 N DUP 6
A00404:156:HV37TDSXX:1:2231:24560:27242 chr6 102816457 N chr6 102816514 N DEL 61
A00404:156:HV37TDSXX:4:2421:25861:35102 chr4 114207444 N chr4 114207499 N DUP 14
A00404:156:HV37TDSXX:3:2603:1687:22576 chr4 114207481 N chr4 114207558 N DEL 17
A00404:156:HV37TDSXX:3:2603:1687:22733 chr4 114207481 N chr4 114207558 N DEL 17
A00404:156:HV37TDSXX:2:1377:25048:20760 chr4 114207481 N chr4 114207558 N DEL 14
A00404:156:HV37TDSXX:3:1564:25699:5071 chr4 114207465 N chr4 114207558 N DEL 15
A00404:155:HV27LDSXX:3:2321:32036:20212 chr4 114207469 N chr4 114207562 N DEL 10
A00404:156:HV37TDSXX:2:2459:1931:26819 chr4 114207470 N chr4 114207563 N DEL 9
A00297:158:HT275DSXX:1:1312:24578:24330 chr7 656718 N chr7 657132 N DEL 8
A00404:156:HV37TDSXX:4:1204:2329:8594 chr7 656967 N chr7 657092 N DEL 5
A00297:158:HT275DSXX:3:2319:13322:8187 chr7 656948 N chr7 657253 N DEL 2
A00404:156:HV37TDSXX:3:1426:11026:1642 chr7 657137 N chr7 657388 N DUP 5
A00404:155:HV27LDSXX:3:2636:6903:30201 chr7 657056 N chr7 657411 N DUP 5
A00297:158:HT275DSXX:1:2154:32181:21308 chr15 101095928 N chr15 101096447 N DEL 5
A00404:156:HV37TDSXX:2:1407:8214:20948 chr15 101095963 N chr15 101096297 N DEL 10
A00297:158:HT275DSXX:2:1513:11496:9533 chr15 101095965 N chr15 101096114 N DEL 5
A00297:158:HT275DSXX:2:2512:6759:21590 chr15 101095965 N chr15 101096114 N DEL 5
A00404:155:HV27LDSXX:3:1229:25635:33583 chr15 101095965 N chr15 101096114 N DEL 5
A00404:155:HV27LDSXX:1:2402:3007:13025 chr15 101095965 N chr15 101096114 N DEL 5
A00297:158:HT275DSXX:4:1131:7952:11851 chr15 101095931 N chr15 101096376 N DEL 5
A00404:155:HV27LDSXX:2:1357:12337:12868 chr15 101095901 N chr15 101096235 N DEL 5
A00404:156:HV37TDSXX:4:1115:1777:4601 chr15 101095974 N chr15 101096049 N DEL 5
A00404:155:HV27LDSXX:3:2628:10836:7921 chr15 101095974 N chr15 101096049 N DEL 5
A00404:155:HV27LDSXX:1:2610:15438:23688 chr15 101095974 N chr15 101096049 N DEL 5
A00404:156:HV37TDSXX:2:2654:5104:4852 chr15 101095974 N chr15 101096049 N DEL 5
A00404:155:HV27LDSXX:1:1141:11695:27414 chr15 101095974 N chr15 101096049 N DEL 6
A00404:155:HV27LDSXX:2:1316:18340:17347 chr15 101095974 N chr15 101096049 N DEL 9
A00404:156:HV37TDSXX:2:2344:22363:13573 chr15 101095938 N chr15 101096307 N DUP 11
A00404:156:HV37TDSXX:1:2324:26485:32205 chr15 101095938 N chr15 101096307 N DUP 10
A00404:155:HV27LDSXX:3:1469:20735:9251 chr15 101095938 N chr15 101096307 N DUP 10
A00297:158:HT275DSXX:3:2160:6072:17550 chr15 101095938 N chr15 101096048 N DUP 10
A00297:158:HT275DSXX:3:2160:6949:17534 chr15 101095938 N chr15 101096307 N DUP 10
A00297:158:HT275DSXX:4:1634:6207:21230 chr15 101095974 N chr15 101096049 N DEL 15
A00297:158:HT275DSXX:3:1430:25536:34820 chr15 101095938 N chr15 101096307 N DUP 10
A00404:156:HV37TDSXX:3:2441:26910:24549 chr15 101095974 N chr15 101096049 N DEL 15
A00297:158:HT275DSXX:2:1336:1145:13683 chr15 101095938 N chr15 101096307 N DUP 10
A00404:156:HV37TDSXX:3:2131:15628:27618 chr15 101095938 N chr15 101096011 N DUP 5
A00404:156:HV37TDSXX:3:2131:15646:27618 chr15 101095938 N chr15 101096307 N DUP 10
A00404:156:HV37TDSXX:2:2651:25907:29606 chr15 101095938 N chr15 101096307 N DUP 10
A00404:155:HV27LDSXX:4:1308:11234:7701 chr15 101095938 N chr15 101096307 N DUP 10
A00404:156:HV37TDSXX:2:1660:8359:31657 chr15 101096113 N chr15 101096225 N DEL 15
A00404:155:HV27LDSXX:3:2466:18132:15452 chr15 101095938 N chr15 101096307 N DUP 10
A00297:158:HT275DSXX:2:1145:16957:32111 chr15 101095927 N chr15 101096037 N DUP 10
A00404:155:HV27LDSXX:3:2236:10999:25927 chr15 101095945 N chr15 101096018 N DUP 5
A00404:156:HV37TDSXX:2:2675:15917:27179 chr15 101096447 N chr15 101096557 N DUP 5
A00297:158:HT275DSXX:1:1314:3070:36620 chr15 101096043 N chr15 101096414 N DEL 4
A00297:158:HT275DSXX:1:2214:32362:34522 chr15 101096011 N chr15 101096382 N DEL 10
A00404:156:HV37TDSXX:3:2235:21775:20697 chr15 101096079 N chr15 101096228 N DEL 5
A00404:156:HV37TDSXX:2:2630:28311:5431 chr15 101096037 N chr15 101096445 N DEL 10
A00404:155:HV27LDSXX:2:1678:21187:13510 chr15 101096076 N chr15 101096447 N DEL 5
A00404:156:HV37TDSXX:3:2632:28393:11365 chr15 101095938 N chr15 101096307 N DUP 10
A00404:155:HV27LDSXX:4:2328:8305:15436 chr15 101095938 N chr15 101096307 N DUP 10
A00404:155:HV27LDSXX:4:2328:9164:9784 chr15 101095938 N chr15 101096307 N DUP 10
A00404:156:HV37TDSXX:1:2541:13223:17597 chr15 101096076 N chr15 101096447 N DEL 5
A00404:156:HV37TDSXX:4:1456:6768:18850 chr15 101096037 N chr15 101096445 N DEL 10
A00404:155:HV27LDSXX:2:1263:26160:20087 chr15 101095938 N chr15 101096085 N DUP 5
A00404:156:HV37TDSXX:3:2359:2383:25598 chr15 101095929 N chr15 101096113 N DUP 1
A00404:155:HV27LDSXX:1:2402:3007:13025 chr15 101095929 N chr15 101096113 N DUP 5
A00404:155:HV27LDSXX:4:2566:17716:24001 chr15 101095937 N chr15 101096049 N DEL 10
A00404:155:HV27LDSXX:3:2657:30915:26882 chr15 101096085 N chr15 101096382 N DEL 5
A00404:155:HV27LDSXX:4:1339:11369:14011 chr15 101095966 N chr15 101096113 N DUP 5
A00404:156:HV37TDSXX:2:2137:26232:36871 chr15 101096111 N chr15 101096297 N DEL 10
A00404:156:HV37TDSXX:1:2324:26485:32205 chr15 101095966 N chr15 101096113 N DUP 5
A00404:156:HV37TDSXX:2:2344:22363:13573 chr15 101095966 N chr15 101096113 N DUP 5
A00404:156:HV37TDSXX:2:1269:20989:7842 chr15 101095938 N chr15 101096085 N DUP 5
A00297:158:HT275DSXX:1:2524:32181:27884 chr15 101096085 N chr15 101096197 N DEL 8
A00404:155:HV27LDSXX:1:2342:9100:11303 chr15 101096225 N chr15 101096372 N DUP 10
A00404:155:HV27LDSXX:2:2202:8585:18427 chr15 101095949 N chr15 101096022 N DUP 5
A00404:156:HV37TDSXX:1:2275:25934:22326 chr15 101095949 N chr15 101096022 N DUP 5
A00297:158:HT275DSXX:3:1308:10655:7138 chr15 101095966 N chr15 101096076 N DUP 5
A00297:158:HT275DSXX:3:1308:11505:6856 chr15 101095966 N chr15 101096076 N DUP 5
A00404:156:HV37TDSXX:3:2374:17716:36432 chr15 101096085 N chr15 101096197 N DEL 9
A00404:155:HV27LDSXX:1:2174:30716:7216 chr15 101096114 N chr15 101096446 N DUP 5
A00297:158:HT275DSXX:3:1226:24921:17127 chr15 101095965 N chr15 101096151 N DEL 5
A00297:158:HT275DSXX:2:2401:20356:24345 chr15 101095965 N chr15 101096151 N DEL 5
A00404:155:HV27LDSXX:3:2142:27688:16313 chr15 101095928 N chr15 101096151 N DEL 5
A00404:156:HV37TDSXX:2:2675:15917:27179 chr15 101095928 N chr15 101096151 N DEL 5
A00297:158:HT275DSXX:1:2362:13539:32769 chr15 101095933 N chr15 101096156 N DEL 5
A00404:155:HV27LDSXX:4:2328:8305:15436 chr15 101095933 N chr15 101096156 N DEL 5
A00404:155:HV27LDSXX:4:2328:9164:9784 chr15 101096188 N chr15 101096335 N DUP 10
A00404:156:HV37TDSXX:2:2568:22227:31187 chr15 101095936 N chr15 101096194 N DUP 5
A00404:155:HV27LDSXX:4:1554:18548:31454 chr15 101095936 N chr15 101096194 N DUP 5
A00404:155:HV27LDSXX:2:1409:5312:36119 chr15 101095936 N chr15 101096194 N DUP 5
A00404:156:HV37TDSXX:1:2471:16378:16705 chr15 101095936 N chr15 101096194 N DUP 5
A00404:155:HV27LDSXX:4:2417:31584:2675 chr15 101095942 N chr15 101096200 N DUP 5
A00404:155:HV27LDSXX:4:2417:31602:2675 chr15 101095936 N chr15 101096194 N DUP 5
A00404:156:HV37TDSXX:4:1672:17454:7012 chr15 101095929 N chr15 101096076 N DUP 5
A00404:156:HV37TDSXX:2:1350:27633:3693 chr15 101095941 N chr15 101096125 N DUP 5
A00404:156:HV37TDSXX:3:1305:19895:24298 chr15 101096259 N chr15 101096593 N DEL 10
A00297:158:HT275DSXX:2:2231:1371:24032 chr15 101095941 N chr15 101096125 N DUP 5
A00404:155:HV27LDSXX:1:1669:31241:13416 chr15 101096447 N chr15 101096557 N DUP 5
A00297:158:HT275DSXX:3:2554:6198:12790 chr15 101095964 N chr15 101096222 N DUP 2
A00404:156:HV37TDSXX:1:2468:30047:10817 chr15 101096076 N chr15 101096225 N DEL 7
A00404:155:HV27LDSXX:3:2473:6180:9032 chr15 101096076 N chr15 101096225 N DEL 10
A00297:158:HT275DSXX:4:1116:22046:35509 chr15 101095963 N chr15 101096556 N DEL 5
A00404:156:HV37TDSXX:4:1244:2266:35196 chr15 101096080 N chr15 101096229 N DEL 5
A00404:155:HV27LDSXX:2:1454:32660:23015 chr15 101095937 N chr15 101096049 N DEL 5
A00297:158:HT275DSXX:3:2366:32262:17315 chr15 101095904 N chr15 101096051 N DUP 4
A00404:155:HV27LDSXX:2:1454:32660:23015 chr15 101096447 N chr15 101096557 N DUP 5
A00404:155:HV27LDSXX:3:2551:16297:24236 chr15 101096007 N chr15 101096526 N DEL 6
A00297:158:HT275DSXX:1:2374:13467:2644 chr15 101095938 N chr15 101096011 N DUP 5
A00297:158:HT275DSXX:3:1226:24921:17127 chr15 101096085 N chr15 101096197 N DEL 11
A00404:156:HV37TDSXX:3:2178:4282:7153 chr15 101095938 N chr15 101096085 N DUP 12
A00297:158:HT275DSXX:3:1472:2853:36933 chr15 101096085 N chr15 101096197 N DEL 11
A00297:158:HT275DSXX:4:2551:30255:34350 chr15 101096085 N chr15 101096197 N DEL 10
A00404:155:HV27LDSXX:2:2219:14118:24377 chr15 101096150 N chr15 101096521 N DEL 10
A00297:158:HT275DSXX:3:2329:25780:2832 chr15 101096085 N chr15 101096197 N DEL 10
A00297:158:HT275DSXX:1:2441:18701:16720 chr15 101096085 N chr15 101096197 N DEL 10
A00297:158:HT275DSXX:1:2441:18719:16720 chr15 101096077 N chr15 101096448 N DEL 5
A00297:158:HT275DSXX:2:1307:8079:7717 chr15 101096085 N chr15 101096197 N DEL 10
A00404:155:HV27LDSXX:4:2615:13340:24439 chr15 101096085 N chr15 101096197 N DEL 10
A00404:156:HV37TDSXX:2:1350:27633:3693 chr15 101096085 N chr15 101096197 N DEL 10
A00404:155:HV27LDSXX:4:2503:20112:20603 chr15 101096198 N chr15 101096456 N DUP 5
A00297:158:HT275DSXX:3:1404:26892:10864 chr15 101096152 N chr15 101096523 N DEL 5
A00404:156:HV37TDSXX:2:2158:29243:20008 chr15 101096152 N chr15 101096523 N DEL 5
A00404:156:HV37TDSXX:4:1323:7527:27211 chr15 101096042 N chr15 101096524 N DEL 14
A00404:156:HV37TDSXX:3:1553:11180:33254 chr15 101096152 N chr15 101096523 N DEL 5
A00297:158:HT275DSXX:4:1128:16911:3443 chr15 101096234 N chr15 101096603 N DUP 15
A00404:155:HV27LDSXX:2:2420:1253:35383 chr15 101095970 N chr15 101096526 N DEL 5
A00404:156:HV37TDSXX:4:1124:14244:30765 chr15 101096076 N chr15 101096521 N DEL 10
A00404:156:HV37TDSXX:1:2504:32814:5431 chr15 101095970 N chr15 101096526 N DEL 5
A00404:155:HV27LDSXX:3:2551:16297:24236 chr15 101095970 N chr15 101096526 N DEL 5
A00404:155:HV27LDSXX:3:2106:14859:32330 chr15 101096076 N chr15 101096521 N DEL 10
A00404:155:HV27LDSXX:3:2154:2899:16752 chr15 101096234 N chr15 101096566 N DUP 15
A00404:155:HV27LDSXX:1:2334:16758:16016 chr15 101095970 N chr15 101096526 N DEL 5
A00404:156:HV37TDSXX:3:2210:10646:23437 chr15 101096080 N chr15 101096525 N DEL 10
A00297:158:HT275DSXX:3:2450:10908:35070 chr15 101096234 N chr15 101096566 N DUP 11
A00404:156:HV37TDSXX:2:2568:22227:31187 chr15 101096450 N chr15 101096597 N DUP 2
A00297:158:HT275DSXX:4:2551:30255:34350 chr15 101096593 N chr15 101096666 N DUP 15
A00404:155:HV27LDSXX:4:1116:29405:29841 chr15 101096019 N chr15 101096501 N DEL 5
A00297:158:HT275DSXX:4:1116:22046:35509 chr15 101096029 N chr15 101096511 N DEL 3
A00404:156:HV37TDSXX:1:2471:16378:16705 chr15 101096333 N chr15 101096556 N DEL 5
A00404:156:HV37TDSXX:2:1667:6126:29293 chr15 101096234 N chr15 101096566 N DUP 15
A00404:155:HV27LDSXX:1:2365:12020:10034 chr15 101096234 N chr15 101096566 N DUP 15
A00404:156:HV37TDSXX:1:1109:11939:29246 chr15 101096234 N chr15 101096566 N DUP 15
A00404:155:HV27LDSXX:4:1339:11369:14011 chr15 101096039 N chr15 101096521 N DEL 5
A00404:155:HV27LDSXX:2:1432:26964:10676 chr15 101096076 N chr15 101096521 N DEL 10
A00297:158:HT275DSXX:1:2524:32181:27884 chr15 101096234 N chr15 101096566 N DUP 15
A00297:158:HT275DSXX:2:2401:20347:24361 chr15 101096307 N chr15 101096419 N DEL 13
A00297:158:HT275DSXX:2:2401:20356:24345 chr15 101096307 N chr15 101096419 N DEL 15
A00404:155:HV27LDSXX:1:1669:31241:13416 chr15 101095938 N chr15 101096307 N DUP 10
A00404:156:HV37TDSXX:1:1365:27887:17785 chr15 101096234 N chr15 101096566 N DUP 15
A00404:156:HV37TDSXX:1:1268:12038:13354 chr15 101096234 N chr15 101096566 N DUP 15
A00404:156:HV37TDSXX:4:1310:27208:31735 chr15 101096084 N chr15 101096529 N DEL 7
A00404:155:HV27LDSXX:3:1103:6388:15530 chr15 101095938 N chr15 101096307 N DUP 8
A00404:156:HV37TDSXX:3:1323:13621:7263 chr15 101096307 N chr15 101096419 N DEL 1
A00404:155:HV27LDSXX:2:2419:4463:2174 chr15 101096234 N chr15 101096603 N DUP 11
A00404:156:HV37TDSXX:1:2124:25147:13385 chr15 101096048 N chr15 101096419 N DEL 4
A00297:158:HT275DSXX:3:2230:29894:1188 chr15 101096234 N chr15 101096603 N DUP 9
A00297:158:HT275DSXX:1:2619:8431:7106 chr15 101096234 N chr15 101096603 N DUP 14
A00297:158:HT275DSXX:3:2366:32262:17315 chr15 101096234 N chr15 101096603 N DUP 15
A00297:158:HT275DSXX:1:1469:23999:12211 chr15 101095975 N chr15 101096344 N DUP 10
A00404:155:HV27LDSXX:2:1678:21187:13510 chr15 101096483 N chr15 101096632 N DEL 15
A00404:156:HV37TDSXX:3:1204:15031:34006 chr15 101096483 N chr15 101096632 N DEL 15
A00404:155:HV27LDSXX:1:2334:16758:16016 chr15 101096483 N chr15 101096632 N DEL 15
A00404:155:HV27LDSXX:1:2334:16893:15906 chr15 101096483 N chr15 101096632 N DEL 15
A00404:155:HV27LDSXX:4:1565:18041:8500 chr15 101096483 N chr15 101096632 N DEL 15
A00404:155:HV27LDSXX:4:2565:16975:16203 chr15 101096483 N chr15 101096632 N DEL 15
A00404:155:HV27LDSXX:4:2449:6189:28119 chr15 101096483 N chr15 101096632 N DEL 15
A00404:155:HV27LDSXX:1:1617:18313:32017 chr15 101096483 N chr15 101096632 N DEL 15
A00297:158:HT275DSXX:4:2445:9634:31798 chr15 101096483 N chr15 101096632 N DEL 15
A00297:158:HT275DSXX:2:2231:1371:24032 chr15 101096483 N chr15 101096632 N DEL 14
A00404:156:HV37TDSXX:2:2678:7563:21042 chr15 101096483 N chr15 101096632 N DEL 13
A00404:156:HV37TDSXX:3:2374:17716:36432 chr15 101096483 N chr15 101096632 N DEL 6
A00404:155:HV27LDSXX:3:2142:27688:16313 chr15 101096483 N chr15 101096632 N DEL 9
A00404:156:HV37TDSXX:2:1342:5113:8187 chr15 101096483 N chr15 101096632 N DEL 8
A00404:155:HV27LDSXX:2:2419:4463:2174 chr15 101095928 N chr15 101096632 N DEL 5
A00404:155:HV27LDSXX:3:1537:22987:1344 chr15 101095928 N chr15 101096632 N DEL 5
A00404:156:HV37TDSXX:1:1264:2428:1125 chr15 101095931 N chr15 101096635 N DEL 5
A00404:156:HV37TDSXX:3:2116:29966:35070 chr15 101095928 N chr15 101096632 N DEL 5
A00404:155:HV27LDSXX:4:2425:20446:21934 chr15 101095935 N chr15 101096639 N DEL 5
A00404:156:HV37TDSXX:3:1138:20076:26772 chr15 101096013 N chr15 101096643 N DEL 4
A00404:155:HV27LDSXX:3:1165:23800:28995 chr8 6104563 N chr8 6104666 N DEL 4
A00297:158:HT275DSXX:1:2231:5294:14262 chr7 2267970 N chr7 2268127 N DEL 5
A00297:158:HT275DSXX:1:1304:24668:21386 chr7 2267914 N chr7 2268069 N DUP 5
A00297:158:HT275DSXX:1:1468:5403:33708 chr7 2268175 N chr7 2268325 N DEL 9
A00404:155:HV27LDSXX:2:2241:24587:21840 chr7 2268185 N chr7 2268285 N DEL 10
A00297:158:HT275DSXX:1:1468:5403:33708 chr7 2268186 N chr7 2268237 N DEL 5
A00297:158:HT275DSXX:1:1468:5575:33755 chr7 2268185 N chr7 2268236 N DEL 5
A00404:155:HV27LDSXX:2:2241:24587:21840 chr7 2268185 N chr7 2268285 N DEL 15
A00404:155:HV27LDSXX:2:1378:28438:20369 chr7 2267929 N chr7 2268086 N DEL 5
A00297:158:HT275DSXX:4:2624:10664:27665 chr7 2268185 N chr7 2268236 N DEL 16
A00404:156:HV37TDSXX:3:1563:10402:12179 chr21 42267578 N chr21 42267953 N DEL 4
A00404:156:HV37TDSXX:3:1622:13386:28369 chr21 42267514 N chr21 42267614 N DEL 7
A00297:158:HT275DSXX:2:2667:25563:24345 chr21 42267674 N chr21 42267917 N DEL 7
A00404:155:HV27LDSXX:4:1208:12129:34616 chr21 42267449 N chr21 42267714 N DEL 1
A00297:158:HT275DSXX:2:1405:26549:24737 chr21 42267814 N chr21 42267969 N DEL 11
A00297:158:HT275DSXX:3:1178:15917:36010 chr21 42267730 N chr21 42267984 N DEL 9
A00404:155:HV27LDSXX:2:1375:18249:19069 chr21 42267699 N chr21 42268008 N DEL 5
A00404:155:HV27LDSXX:1:2340:9896:19038 chr16 88247162 N chr16 88247488 N DEL 3
A00297:158:HT275DSXX:4:1662:26313:21950 chr16 88247168 N chr16 88247482 N DEL 9
A00297:158:HT275DSXX:4:1662:26594:21746 chr16 88247168 N chr16 88247482 N DEL 9
A00404:155:HV27LDSXX:2:1346:14000:35164 chr16 88247176 N chr16 88247678 N DEL 13
A00297:158:HT275DSXX:3:1537:18114:22874 chr16 88247176 N chr16 88247678 N DEL 13
A00297:158:HT275DSXX:1:1521:4661:2957 chr16 88247140 N chr16 88247554 N DEL 50
A00404:156:HV37TDSXX:2:1307:21224:3865 chr16 88247176 N chr16 88247678 N DEL 17
A00404:155:HV27LDSXX:4:2176:19226:20228 chr16 88247176 N chr16 88247678 N DEL 17
A00404:156:HV37TDSXX:2:2647:15239:16454 chr16 88247176 N chr16 88247678 N DEL 17
A00404:155:HV27LDSXX:1:2519:18304:11365 chr16 88247176 N chr16 88247678 N DEL 17
A00297:158:HT275DSXX:2:2343:17481:20588 chr16 88247176 N chr16 88247678 N DEL 17
A00404:156:HV37TDSXX:3:1425:20211:36151 chr16 88247176 N chr16 88247678 N DEL 17
A00297:158:HT275DSXX:2:2413:31132:7341 chr16 88247008 N chr16 88247177 N DEL 13
A00297:158:HT275DSXX:2:1571:31729:15013 chr16 88247201 N chr16 88247641 N DUP 11
A00297:158:HT275DSXX:2:2570:29152:21793 chr16 88247201 N chr16 88247641 N DUP 11
A00404:156:HV37TDSXX:3:1475:17960:11303 chr16 88247201 N chr16 88247641 N DUP 7
A00404:155:HV27LDSXX:4:1243:32045:34444 chr16 88247214 N chr16 88247459 N DUP 7
A00297:158:HT275DSXX:1:2109:27154:27101 chr16 88247218 N chr16 88247851 N DUP 5
A00297:158:HT275DSXX:1:2434:15926:36683 chr16 88247220 N chr16 88247299 N DUP 9
A00404:155:HV27LDSXX:4:2309:16477:7263 chr16 88246947 N chr16 88247367 N DUP 5
A00297:158:HT275DSXX:2:2343:12174:28244 chr16 88246979 N chr16 88247380 N DUP 9
A00297:158:HT275DSXX:2:1470:23448:36464 chr16 88247389 N chr16 88247485 N DEL 12
A00297:158:HT275DSXX:1:2526:3803:2628 chr16 88246969 N chr16 88247457 N DUP 3
A00404:155:HV27LDSXX:1:1313:15365:35055 chr16 88246969 N chr16 88247457 N DUP 8
A00297:158:HT275DSXX:3:1139:5385:3928 chr16 88247366 N chr16 88247483 N DUP 14
A00404:155:HV27LDSXX:4:1143:5394:13745 chr16 88246969 N chr16 88247457 N DUP 12
A00404:156:HV37TDSXX:3:2563:18846:24674 chr16 88246980 N chr16 88247390 N DEL 29
A00404:156:HV37TDSXX:2:1120:1506:8641 chr16 88246980 N chr16 88247390 N DEL 29
A00404:156:HV37TDSXX:2:2263:3314:21574 chr16 88246981 N chr16 88247391 N DEL 14
A00297:158:HT275DSXX:2:2413:31132:7341 chr16 88246969 N chr16 88247457 N DUP 25
A00404:155:HV27LDSXX:1:1652:31864:34695 chr16 88246969 N chr16 88247457 N DUP 26
A00404:155:HV27LDSXX:1:1652:32226:35415 chr16 88246969 N chr16 88247457 N DUP 16
A00404:155:HV27LDSXX:1:2518:25174:29653 chr16 88247048 N chr16 88247530 N DEL 24
A00404:155:HV27LDSXX:4:1111:32371:34006 chr16 88247048 N chr16 88247530 N DEL 24
A00297:158:HT275DSXX:1:2244:5665:13056 chr16 88247048 N chr16 88247530 N DEL 24
A00404:155:HV27LDSXX:1:2519:18304:11365 chr16 88247048 N chr16 88247530 N DEL 23
A00404:156:HV37TDSXX:2:1661:20500:30796 chr16 88247049 N chr16 88247531 N DEL 11
A00404:155:HV27LDSXX:1:1239:30517:8813 chr16 88247048 N chr16 88247530 N DEL 22
A00404:155:HV27LDSXX:3:1403:16911:7326 chr16 88247048 N chr16 88247530 N DEL 22
A00404:156:HV37TDSXX:2:2647:15239:16454 chr16 88247048 N chr16 88247530 N DEL 13
A00297:158:HT275DSXX:2:1432:30011:21809 chr16 88247357 N chr16 88247508 N DEL 2
A00404:155:HV27LDSXX:1:1664:20817:20572 chr16 88247048 N chr16 88247530 N DEL 13
A00404:155:HV27LDSXX:1:2318:6876:25520 chr16 88247008 N chr16 88247530 N DEL 13
A00297:158:HT275DSXX:2:2632:14380:2253 chr16 88247008 N chr16 88247530 N DEL 13
A00404:156:HV37TDSXX:1:2113:32181:9659 chr16 88247008 N chr16 88247530 N DEL 13
A00404:155:HV27LDSXX:3:2472:21956:36761 chr16 88246910 N chr16 88247530 N DEL 13
A00297:158:HT275DSXX:4:1652:31015:30248 chr16 88246910 N chr16 88247530 N DEL 13
A00404:155:HV27LDSXX:2:1320:22037:32236 chr16 88247062 N chr16 88247544 N DEL 1
A00404:155:HV27LDSXX:3:2472:21956:36761 chr16 88247697 N chr16 88247895 N DEL 28
A00297:158:HT275DSXX:3:1147:30255:14873 chr16 88247245 N chr16 88247751 N DEL 9
A00404:155:HV27LDSXX:1:2342:20410:29011 chr16 88247245 N chr16 88247751 N DEL 9
A00404:155:HV27LDSXX:4:2322:13720:24659 chr16 88247245 N chr16 88247751 N DEL 9
A00404:156:HV37TDSXX:3:1633:25572:12054 chr16 88247245 N chr16 88247751 N DEL 9
A00404:156:HV37TDSXX:3:1143:3369:16752 chr16 88247246 N chr16 88247752 N DEL 9
A00297:158:HT275DSXX:1:2577:15374:7075 chr16 88247252 N chr16 88247758 N DEL 8
A00404:156:HV37TDSXX:4:1648:18304:5008 chr16 88247253 N chr16 88247759 N DEL 7
A00297:158:HT275DSXX:2:2632:14380:2253 chr16 88247254 N chr16 88247760 N DEL 6
A00297:158:HT275DSXX:3:2431:10429:32456 chr5 153296468 N chr5 153296644 N DEL 5
A00297:158:HT275DSXX:3:2431:9670:32894 chr5 153296476 N chr5 153296652 N DEL 5
A00404:155:HV27LDSXX:1:1666:15709:22905 chr5 153296643 N chr5 153296819 N DEL 5
A00404:155:HV27LDSXX:1:2232:7129:21919 chr5 153296643 N chr5 153296819 N DEL 5
A00404:156:HV37TDSXX:2:2362:28203:25222 chr5 153296636 N chr5 153296909 N DEL 5
A00404:155:HV27LDSXX:2:1661:19407:4476 chr5 153296663 N chr5 153296837 N DUP 5
A00404:155:HV27LDSXX:4:1301:20446:36245 chr5 153296663 N chr5 153296837 N DUP 5
A00404:155:HV27LDSXX:3:2219:9751:4633 chr5 153296734 N chr5 153296830 N DUP 1
A00404:155:HV27LDSXX:4:1649:4327:36135 chr5 153296933 N chr5 153297104 N DEL 21
A00404:156:HV37TDSXX:3:2624:2103:33004 chr5 153296608 N chr5 153296882 N DEL 21
A00404:155:HV27LDSXX:2:2660:14950:32863 chr5 153296528 N chr5 153296976 N DEL 5
A00404:155:HV27LDSXX:4:1666:6081:31093 chr6 27485638 N chr6 27486205 N DUP 6
A00297:158:HT275DSXX:3:1308:30020:23484 chr6 27485809 N chr6 27485927 N DEL 12
A00297:158:HT275DSXX:3:1234:32307:4961 chr6 27485811 N chr6 27486085 N DEL 19
A00404:156:HV37TDSXX:2:2333:5050:17722 chr6 27485795 N chr6 27486109 N DEL 5
A00404:156:HV37TDSXX:1:2173:21603:29199 chr14 80354774 N chr14 80354872 N DEL 11
A00404:156:HV37TDSXX:2:2340:28682:7232 chr14 80354771 N chr14 80354869 N DEL 14
A00404:155:HV27LDSXX:4:1127:23231:8844 chr12 121993596 N chr12 121993788 N DUP 3
A00297:158:HT275DSXX:2:2443:21893:10974 chr12 117583510 N chr12 117583563 N DEL 13
A00404:156:HV37TDSXX:1:1261:28664:3223 chr12 117583510 N chr12 117583563 N DEL 13
A00404:156:HV37TDSXX:1:2420:19135:18443 chr12 117583513 N chr12 117583566 N DEL 12
A00404:156:HV37TDSXX:2:2651:9751:25332 chr19 48011339 N chr19 48011404 N DEL 4
A00404:156:HV37TDSXX:2:1524:14760:30874 chr19 48011339 N chr19 48011404 N DEL 9
A00404:156:HV37TDSXX:2:1524:14778:31657 chr19 48011339 N chr19 48011404 N DEL 9
A00404:156:HV37TDSXX:4:2123:4237:19820 chr19 48011339 N chr19 48011648 N DEL 11
A00404:156:HV37TDSXX:2:2461:5113:16705 chr19 48011400 N chr19 48011497 N DUP 5
A00404:156:HV37TDSXX:3:2176:18548:15608 chr19 48011380 N chr19 48011596 N DUP 4
A00404:155:HV27LDSXX:1:1524:9453:10911 chr19 48011380 N chr19 48011596 N DUP 6
A00297:158:HT275DSXX:2:2423:19633:8625 chr19 48011282 N chr19 48011604 N DEL 8
A00297:158:HT275DSXX:2:2423:19678:8609 chr19 48011282 N chr19 48011604 N DEL 8
A00297:158:HT275DSXX:1:1452:22833:29982 chr19 48011396 N chr19 48011611 N DEL 1
A00404:155:HV27LDSXX:3:1248:1597:21386 chr19 1063325 N chr19 1063438 N DUP 8
A00404:156:HV37TDSXX:1:2169:16333:25488 chr19 1063294 N chr19 1063446 N DUP 25
A00297:158:HT275DSXX:4:1567:32334:27179 chr19 1063349 N chr19 1063464 N DEL 15
A00404:155:HV27LDSXX:2:1203:25545:7936 chr19 1063349 N chr19 1063464 N DEL 15
A00297:158:HT275DSXX:1:2544:25870:17895 chr19 1063349 N chr19 1063464 N DEL 15
A00404:156:HV37TDSXX:1:1540:1353:32863 chr20 43293284 N chr20 43293395 N DUP 8
A00297:158:HT275DSXX:1:2561:2853:25880 chr19 6730599 N chr19 6730777 N DEL 5
A00404:155:HV27LDSXX:2:2512:18421:20400 chr15 94814138 N chr15 94814295 N DEL 11
A00404:155:HV27LDSXX:2:2206:25870:27445 chr10 92674862 N chr10 92674959 N DUP 5
A00404:155:HV27LDSXX:3:1102:29432:22247 chr10 92674862 N chr10 92674959 N DUP 5
A00297:158:HT275DSXX:3:1206:12491:3114 chr10 92674946 N chr10 92675121 N DEL 9
A00297:158:HT275DSXX:3:2271:2663:27962 chr10 92674969 N chr10 92675270 N DUP 8
A00297:158:HT275DSXX:3:1102:28203:10974 chr10 92675054 N chr10 92675279 N DEL 10
A00404:155:HV27LDSXX:1:2114:26982:19946 chr10 92674948 N chr10 92675123 N DUP 12
A00404:156:HV37TDSXX:4:2357:21070:8015 chr10 92674904 N chr10 92675205 N DUP 5
A00404:155:HV27LDSXX:4:2663:12644:32315 chr10 92674855 N chr10 92675129 N DEL 3
A00404:155:HV27LDSXX:2:2427:2727:5682 chr10 92675152 N chr10 92675278 N DUP 5
A00404:156:HV37TDSXX:1:1435:15655:19210 chr10 92674890 N chr10 92675240 N DUP 5
A00297:158:HT275DSXX:1:1329:29713:36667 chr10 92674890 N chr10 92675240 N DUP 5
A00297:158:HT275DSXX:4:1634:11758:14215 chr10 92674978 N chr10 92675154 N DEL 5
A00404:155:HV27LDSXX:4:2621:4146:30718 chr10 92675012 N chr10 92675188 N DEL 10
A00404:155:HV27LDSXX:1:2159:4191:28134 chr10 92674862 N chr10 92675086 N DUP 4
A00297:158:HT275DSXX:4:2652:13440:9267 chr10 92674841 N chr10 92675242 N DEL 5
A00404:155:HV27LDSXX:4:1104:32434:27289 chr2 63809245 N chr2 63809324 N DUP 1
A00297:158:HT275DSXX:4:2145:27516:5243 chr2 63809264 N chr2 63809345 N DEL 5
A00297:158:HT275DSXX:4:2569:15953:26522 chr2 63809264 N chr2 63809345 N DEL 5
A00297:158:HT275DSXX:2:1253:28863:14372 chr2 63809347 N chr2 63809472 N DUP 1
A00404:155:HV27LDSXX:4:1223:17870:34757 chr2 63809260 N chr2 63809544 N DEL 30
A00297:158:HT275DSXX:2:2329:21630:13808 chr10 112455486 N chr10 112455627 N DEL 5
A00404:156:HV37TDSXX:1:1611:9688:12477 chr6 169067794 N chr6 169067882 N DEL 9
A00404:155:HV27LDSXX:2:2202:12427:34475 chr11 77098679 N chr11 77098805 N DUP 4
A00404:156:HV37TDSXX:4:2576:20980:24580 chr11 77098679 N chr11 77098805 N DUP 5
A00404:155:HV27LDSXX:1:1276:21251:15154 chr11 77098679 N chr11 77098805 N DUP 5
A00404:156:HV37TDSXX:4:2206:4146:3067 chr11 77098698 N chr11 77098824 N DUP 3
A00404:155:HV27LDSXX:3:2437:3794:11256 chr11 77098682 N chr11 77098857 N DUP 2
A00404:155:HV27LDSXX:2:2214:15103:25300 chr19 9701652 N chr19 9701903 N DEL 7
A00404:156:HV37TDSXX:2:2573:9173:26209 chr19 9701657 N chr19 9701808 N DEL 10
A00297:158:HT275DSXX:3:2647:15899:19413 chr19 9701657 N chr19 9701808 N DEL 10
A00404:156:HV37TDSXX:2:2268:26467:30733 chr19 9701658 N chr19 9701835 N DEL 21
A00404:155:HV27LDSXX:3:1408:21649:16971 chr19 9701740 N chr19 9701845 N DEL 7
A00404:155:HV27LDSXX:3:2407:19416:36777 chr19 9701740 N chr19 9701845 N DEL 7
A00297:158:HT275DSXX:4:2555:28004:10629 chr19 9701740 N chr19 9701845 N DEL 14
A00404:155:HV27LDSXX:4:2572:5122:16501 chr19 9701740 N chr19 9701845 N DEL 15
A00297:158:HT275DSXX:4:1167:19922:22498 chr19 9701740 N chr19 9701845 N DEL 24
A00404:155:HV27LDSXX:2:1374:4074:33912 chr19 9701740 N chr19 9701845 N DEL 29
A00404:156:HV37TDSXX:4:1631:16631:16611 chr19 9701740 N chr19 9701845 N DEL 32
A00404:156:HV37TDSXX:4:1631:16731:16877 chr19 9701740 N chr19 9701845 N DEL 32
A00404:156:HV37TDSXX:1:2523:14959:14184 chr19 9701759 N chr19 9701832 N DEL 29
A00297:158:HT275DSXX:2:2264:3640:28808 chr19 9701759 N chr19 9701832 N DEL 35
A00297:158:HT275DSXX:4:2655:25473:22748 chr19 9701759 N chr19 9701832 N DEL 35
A00297:158:HT275DSXX:2:1671:1931:36401 chr19 9701759 N chr19 9701832 N DEL 35
A00404:156:HV37TDSXX:1:2244:17418:23328 chr19 9701759 N chr19 9701832 N DEL 34
A00404:156:HV37TDSXX:2:2159:25726:12696 chr19 9701759 N chr19 9701832 N DEL 33
A00404:156:HV37TDSXX:2:2270:23194:9471 chr19 9701759 N chr19 9701832 N DEL 33
A00404:155:HV27LDSXX:4:1332:17653:30311 chr19 9701666 N chr19 9701875 N DEL 5
A00404:155:HV27LDSXX:2:1228:6985:3850 chr19 9701675 N chr19 9701884 N DEL 6
A00297:158:HT275DSXX:1:1139:10285:3239 chr19 9701678 N chr19 9701887 N DEL 5
A00404:155:HV27LDSXX:4:1407:20094:9643 chr19 9701760 N chr19 9701909 N DEL 12
A00297:158:HT275DSXX:4:1439:18566:29669 chr19 9701826 N chr19 9701929 N DEL 10
A00404:156:HV37TDSXX:3:2578:19551:26678 chr19 9701861 N chr19 9701938 N DEL 1
A00297:158:HT275DSXX:1:1438:26124:14387 chr9 120495996 N chr9 120496929 N DUP 10
A00297:158:HT275DSXX:2:2215:10836:24956 chr9 120496096 N chr9 120496195 N DEL 4
A00297:158:HT275DSXX:3:1652:10185:11522 chr9 120495989 N chr9 120496214 N DUP 5
A00404:156:HV37TDSXX:2:1561:29586:13620 chr9 120496046 N chr9 120496447 N DUP 5
A00404:155:HV27LDSXX:1:2253:3305:8187 chr9 120496046 N chr9 120496271 N DUP 5
A00404:155:HV27LDSXX:3:2603:25364:30107 chr9 120496148 N chr9 120496632 N DEL 6
A00404:155:HV27LDSXX:4:1472:14805:25535 chr9 120496092 N chr9 120496545 N DUP 1
A00297:158:HT275DSXX:2:1571:4246:7654 chr9 120496148 N chr9 120496632 N DEL 25
A00404:155:HV27LDSXX:3:1669:32099:1470 chr9 120496161 N chr9 120496338 N DEL 5
A00404:155:HV27LDSXX:3:2304:19135:31438 chr9 120495991 N chr9 120496120 N DEL 5
A00404:155:HV27LDSXX:4:2442:27145:7326 chr9 120495994 N chr9 120496123 N DEL 5
A00404:155:HV27LDSXX:2:2311:25717:22576 chr9 120496141 N chr9 120496897 N DUP 3
A00404:156:HV37TDSXX:1:1203:18430:28745 chr9 120495963 N chr9 120496141 N DEL 3
A00404:155:HV27LDSXX:3:1364:10041:17754 chr9 120496161 N chr9 120496338 N DEL 5
A00297:158:HT275DSXX:3:2624:26051:29324 chr9 120496271 N chr9 120496902 N DEL 5
A00297:158:HT275DSXX:2:2127:28610:31814 chr9 120496192 N chr9 120496318 N DUP 5
A00297:158:HT275DSXX:2:1674:17481:4679 chr9 120496175 N chr9 120496350 N DUP 2
A00404:156:HV37TDSXX:1:1605:5439:14638 chr9 120496176 N chr9 120496351 N DUP 1
A00297:158:HT275DSXX:1:2666:21847:6292 chr9 120496186 N chr9 120496540 N DUP 6
A00404:156:HV37TDSXX:4:2448:4490:27367 chr9 120496239 N chr9 120496596 N DEL 5
A00297:158:HT275DSXX:2:1473:4029:35023 chr9 120495965 N chr9 120496192 N DEL 5
A00297:158:HT275DSXX:2:2467:14055:7576 chr9 120495965 N chr9 120496192 N DEL 5
A00404:155:HV27LDSXX:1:2635:2663:22701 chr9 120496239 N chr9 120496596 N DEL 5
A00404:155:HV27LDSXX:3:2137:8838:35712 chr9 120496011 N chr9 120496238 N DEL 5
A00404:155:HV27LDSXX:2:1607:18204:13823 chr9 120496313 N chr9 120496670 N DEL 6
A00404:155:HV27LDSXX:2:1313:4969:1673 chr9 120496313 N chr9 120496670 N DEL 6
A00404:155:HV27LDSXX:3:2107:32271:18552 chr9 120496177 N chr9 120496353 N DUP 7
A00404:155:HV27LDSXX:4:2667:30996:13119 chr9 120495951 N chr9 120496353 N DUP 7
A00404:155:HV27LDSXX:4:1565:24939:21073 chr9 120496320 N chr9 120496628 N DEL 5
A00404:155:HV27LDSXX:1:2312:6596:28479 chr9 120496320 N chr9 120496628 N DEL 5
A00404:156:HV37TDSXX:3:1408:10474:27492 chr9 120496035 N chr9 120496262 N DEL 4
A00404:155:HV27LDSXX:4:2465:20455:17534 chr9 120496177 N chr9 120496353 N DUP 7
A00404:155:HV27LDSXX:3:2563:13819:27712 chr9 120496153 N chr9 120496328 N DUP 5
A00404:156:HV37TDSXX:4:2666:4942:23891 chr9 120496153 N chr9 120496328 N DUP 5
A00404:156:HV37TDSXX:4:1336:27109:18223 chr9 120495976 N chr9 120496281 N DEL 1
A00404:155:HV27LDSXX:1:2547:27199:17096 chr9 120496324 N chr9 120496855 N DUP 5
A00404:155:HV27LDSXX:1:2270:13376:19272 chr9 120496338 N chr9 120496513 N DUP 5
A00404:155:HV27LDSXX:1:2515:18530:12101 chr9 120495961 N chr9 120496718 N DUP 5
A00404:155:HV27LDSXX:3:2441:6668:22122 chr9 120496119 N chr9 120496296 N DEL 5
A00404:156:HV37TDSXX:2:1355:11731:15013 chr9 120496219 N chr9 120496298 N DEL 5
A00404:155:HV27LDSXX:1:2130:7581:28776 chr9 120495992 N chr9 120496346 N DEL 5
A00404:156:HV37TDSXX:2:1235:21802:13761 chr9 120495984 N chr9 120496338 N DEL 5
A00297:158:HT275DSXX:3:1434:2627:8703 chr9 120495984 N chr9 120496338 N DEL 5
A00404:156:HV37TDSXX:1:1607:11171:15170 chr9 120496162 N chr9 120496337 N DUP 5
A00404:156:HV37TDSXX:4:1370:29496:8954 chr9 120496162 N chr9 120496337 N DUP 5
A00404:156:HV37TDSXX:1:1609:15013:26115 chr9 120495984 N chr9 120496338 N DEL 5
A00404:156:HV37TDSXX:3:1375:19289:9596 chr9 120495994 N chr9 120496348 N DEL 3
A00297:158:HT275DSXX:4:2278:31738:23390 chr9 120496226 N chr9 120496583 N DEL 4
A00297:158:HT275DSXX:4:1636:13286:15045 chr9 120496214 N chr9 120496571 N DEL 5
A00297:158:HT275DSXX:4:2155:21151:36526 chr9 120496321 N chr9 120496447 N DUP 10
A00404:155:HV27LDSXX:3:2138:12364:12790 chr9 120496214 N chr9 120496571 N DEL 5
A00404:156:HV37TDSXX:3:2538:15817:7247 chr9 120496214 N chr9 120496571 N DEL 5
A00404:155:HV27LDSXX:2:2540:3152:20353 chr9 120495988 N chr9 120496391 N DEL 5
A00297:158:HT275DSXX:4:1321:2320:27868 chr9 120495989 N chr9 120496392 N DEL 5
A00404:155:HV27LDSXX:3:1364:10041:17754 chr9 120496438 N chr9 120497020 N DUP 5
A00297:158:HT275DSXX:2:1233:23167:6574 chr9 120495997 N chr9 120496400 N DEL 5
A00297:158:HT275DSXX:2:1375:21920:19633 chr9 120496222 N chr9 120496579 N DEL 5
A00404:155:HV27LDSXX:2:2410:24080:34303 chr9 120496004 N chr9 120496407 N DEL 5
A00404:155:HV27LDSXX:1:1609:2157:13338 chr9 120496518 N chr9 120496924 N DEL 4
A00404:155:HV27LDSXX:1:2514:25039:9627 chr9 120496490 N chr9 120496669 N DUP 5
A00404:155:HV27LDSXX:4:2371:4743:26741 chr9 120496530 N chr9 120496934 N DEL 6
A00404:156:HV37TDSXX:3:1563:21142:27430 chr9 120495973 N chr9 120496554 N DUP 5
A00404:155:HV27LDSXX:3:2105:3649:12258 chr9 120496710 N chr9 120496934 N DEL 10
A00404:156:HV37TDSXX:3:2575:20528:30812 chr9 120495973 N chr9 120496554 N DUP 5
A00404:156:HV37TDSXX:2:2620:7193:25379 chr9 120495973 N chr9 120496554 N DUP 5
A00404:155:HV27LDSXX:1:1608:15338:18317 chr9 120496459 N chr9 120496863 N DUP 2
A00404:155:HV27LDSXX:4:2667:30996:13119 chr9 120495973 N chr9 120496554 N DUP 5
A00404:156:HV37TDSXX:3:2575:20528:30812 chr9 120495973 N chr9 120496554 N DUP 5
A00297:158:HT275DSXX:3:2233:5701:9392 chr9 120496486 N chr9 120496537 N DUP 2
A00404:155:HV27LDSXX:1:1145:12825:25113 chr9 120496488 N chr9 120496537 N DUP 9
A00404:155:HV27LDSXX:2:1317:24108:25676 chr9 120495973 N chr9 120496554 N DUP 5
A00297:158:HT275DSXX:2:1323:23791:4805 chr9 120496124 N chr9 120496529 N DEL 19
A00297:158:HT275DSXX:4:2329:19370:27305 chr9 120496127 N chr9 120496532 N DEL 18
A00297:158:HT275DSXX:3:1417:14226:32957 chr9 120495965 N chr9 120496546 N DUP 5
A00297:158:HT275DSXX:4:1237:21124:24831 chr9 120495973 N chr9 120496554 N DUP 5
A00404:155:HV27LDSXX:2:1514:32172:13119 chr9 120496616 N chr9 120497020 N DEL 2
A00404:155:HV27LDSXX:1:2326:29568:22263 chr9 120496127 N chr9 120496532 N DEL 15
A00404:155:HV27LDSXX:2:1514:32172:13119 chr9 120496616 N chr9 120497020 N DEL 6
A00404:155:HV27LDSXX:2:1317:24108:25676 chr9 120496554 N chr9 120496731 N DEL 5
A00297:158:HT275DSXX:2:1628:1787:36245 chr9 120496618 N chr9 120496944 N DEL 5
A00297:158:HT275DSXX:3:1142:3450:31360 chr9 120496306 N chr9 120496533 N DEL 6
A00404:156:HV37TDSXX:2:1169:26639:31501 chr9 120496554 N chr9 120496731 N DEL 5
A00404:155:HV27LDSXX:2:2149:32045:36166 chr9 120496319 N chr9 120496548 N DEL 3
A00404:155:HV27LDSXX:3:2104:23285:10441 chr9 120496186 N chr9 120496542 N DEL 5
A00404:155:HV27LDSXX:3:1326:13738:12007 chr9 120496537 N chr9 120496942 N DUP 7
A00404:156:HV37TDSXX:2:2468:5891:3521 chr9 120496183 N chr9 120496535 N DEL 7
A00404:155:HV27LDSXX:3:1420:22037:27915 chr9 120496566 N chr9 120496743 N DEL 10
A00404:155:HV27LDSXX:3:2454:25843:20040 chr9 120496392 N chr9 120496571 N DUP 5
A00297:158:HT275DSXX:4:1608:14651:29183 chr9 120496702 N chr9 120496928 N DEL 3
A00404:155:HV27LDSXX:2:1211:10484:4867 chr9 120496272 N chr9 120496676 N DUP 1
A00404:156:HV37TDSXX:2:1441:31801:13009 chr9 120496698 N chr9 120496924 N DEL 3
A00404:156:HV37TDSXX:4:2420:7853:21574 chr9 120496228 N chr9 120496585 N DEL 1
A00404:155:HV27LDSXX:3:2104:23285:10441 chr9 120496638 N chr9 120497040 N DUP 5
A00404:156:HV37TDSXX:2:2567:8205:15859 chr9 120496526 N chr9 120496658 N DEL 1
A00404:155:HV27LDSXX:3:1317:10013:6778 chr9 120496103 N chr9 120496631 N DEL 7
A00404:156:HV37TDSXX:3:1112:26078:29904 chr9 120496546 N chr9 120496675 N DEL 2
A00297:158:HT275DSXX:1:2537:30653:8015 chr9 120496718 N chr9 120496945 N DEL 12
A00297:158:HT275DSXX:1:2572:28149:36151 chr9 120496186 N chr9 120496670 N DEL 5
A00297:158:HT275DSXX:1:2572:28791:34006 chr9 120496186 N chr9 120496670 N DEL 5
A00404:155:HV27LDSXX:2:1571:7328:34319 chr9 120495970 N chr9 120496727 N DUP 5
A00297:158:HT275DSXX:2:2204:3721:21120 chr9 120496732 N chr9 120496960 N DEL 5
A00297:158:HT275DSXX:3:1373:11053:12555 chr9 120496340 N chr9 120496697 N DEL 5
A00404:155:HV27LDSXX:4:2469:22643:26678 chr9 120495969 N chr9 120496728 N DEL 10
A00297:158:HT275DSXX:3:1405:30237:36417 chr9 120496825 N chr9 120496924 N DEL 9
A00404:155:HV27LDSXX:4:1441:13612:27101 chr9 120496516 N chr9 120496873 N DEL 10
A00404:156:HV37TDSXX:1:1116:29161:15452 chr9 120496333 N chr9 120496898 N DEL 34
A00404:156:HV37TDSXX:4:1635:7139:5963 chr6 37100641 N chr6 37100932 N DEL 5
A00404:156:HV37TDSXX:1:2352:15004:1016 chr6 37100641 N chr6 37100932 N DEL 5
A00404:155:HV27LDSXX:2:2240:22516:34632 chr6 37100641 N chr6 37100932 N DEL 5
A00297:158:HT275DSXX:2:2638:19072:14982 chr19 16349240 N chr19 16349538 N DEL 5
A00404:155:HV27LDSXX:2:2654:28763:18959 chr19 16349240 N chr19 16349538 N DEL 5
A00404:156:HV37TDSXX:1:2362:8034:26428 chr19 16349256 N chr19 16349552 N DUP 5
A00297:158:HT275DSXX:1:1178:1181:23390 chr19 16349256 N chr19 16349552 N DUP 5
A00297:158:HT275DSXX:1:2346:15194:26052 chr19 16349262 N chr19 16349558 N DUP 5
A00404:155:HV27LDSXX:2:1672:5122:9612 chr19 16349262 N chr19 16349558 N DUP 5
A00297:158:HT275DSXX:2:2305:23647:10128 chr19 16349263 N chr19 16349559 N DUP 5
A00297:158:HT275DSXX:1:1203:32723:25661 chr1 187738572 N chr1 187738653 N DUP 1
A00404:156:HV37TDSXX:2:1247:32886:36464 chr3 45890432 N chr3 45890514 N DEL 3
A00404:156:HV37TDSXX:3:1432:28131:13698 chr3 45890431 N chr3 45890513 N DEL 4
A00404:156:HV37TDSXX:4:2133:21007:4679 chr3 45890430 N chr3 45890512 N DEL 5
A00297:158:HT275DSXX:1:1652:1425:19085 chr5 126596225 N chr5 126596521 N DUP 5
A00404:155:HV27LDSXX:2:1517:26214:23970 chr5 126596225 N chr5 126596521 N DUP 5
A00404:155:HV27LDSXX:2:1517:26666:23657 chr5 126596225 N chr5 126596521 N DUP 5
A00404:156:HV37TDSXX:3:2459:3278:10488 chr5 126596186 N chr5 126596482 N DUP 3
A00404:156:HV37TDSXX:3:2457:3712:34225 chr5 126596433 N chr5 126596740 N DUP 5
A00404:156:HV37TDSXX:1:1237:10999:32315 chr5 126596448 N chr5 126596757 N DEL 25
A00404:156:HV37TDSXX:3:2244:7961:23296 chr5 126596452 N chr5 126596761 N DEL 15
A00297:158:HT275DSXX:2:1665:4001:5353 chr11 472061 N chr11 472185 N DEL 5
A00404:155:HV27LDSXX:4:2523:2528:26005 chr11 472084 N chr11 472206 N DUP 5
A00297:158:HT275DSXX:3:2538:9959:29919 chr9 17927484 N chr9 17927573 N DUP 5
A00404:156:HV37TDSXX:4:1166:24948:29042 chr1 28823812 N chr1 28823948 N DEL 5
A00297:158:HT275DSXX:1:2571:31204:11224 chr18 76508713 N chr18 76508904 N DEL 7
A00404:156:HV37TDSXX:1:2556:24071:28119 chr18 76508713 N chr18 76508904 N DEL 7
A00404:155:HV27LDSXX:4:2575:2347:10942 chr18 76508915 N chr18 76509096 N DEL 2
A00404:156:HV37TDSXX:3:2223:29423:8422 chr2 129914492 N chr2 129914743 N DEL 17
A00404:156:HV37TDSXX:3:2223:29423:8422 chr2 129914488 N chr2 129914739 N DEL 35
A00404:156:HV37TDSXX:1:1164:9444:3724 chr2 129914582 N chr2 129914692 N DUP 5
A00404:156:HV37TDSXX:4:1223:24930:9565 chr2 129914549 N chr2 129914660 N DEL 1
A00404:156:HV37TDSXX:4:1310:28122:3255 chr2 129914799 N chr2 129914858 N DEL 5
A00404:156:HV37TDSXX:4:1252:17752:36526 chr2 129914738 N chr2 129914971 N DEL 43
A00404:156:HV37TDSXX:3:1614:19506:27946 chr2 129914798 N chr2 129915058 N DUP 5
A00297:158:HT275DSXX:2:1522:16640:32471 chr2 129914890 N chr2 129915389 N DEL 8
A00404:155:HV27LDSXX:3:1369:11071:4977 chr2 129914554 N chr2 129914835 N DEL 1
A00404:156:HV37TDSXX:2:2659:1958:33880 chr2 129914903 N chr2 129915319 N DEL 30
A00297:158:HT275DSXX:3:1653:13033:6590 chr2 129914478 N chr2 129915017 N DUP 5
A00404:156:HV37TDSXX:3:2449:11659:33395 chr2 129914702 N chr2 129914935 N DEL 5
A00404:156:HV37TDSXX:1:1502:10565:22075 chr2 129915071 N chr2 129915209 N DEL 16
A00297:158:HT275DSXX:3:1165:17969:20243 chr2 129914677 N chr2 129915105 N DEL 41
A00297:158:HT275DSXX:4:2501:23068:22811 chr2 129915134 N chr2 129915218 N DEL 12
A00297:158:HT275DSXX:2:1522:16640:32471 chr2 129915200 N chr2 129915284 N DEL 5
A00404:156:HV37TDSXX:2:1659:4273:27618 chr2 129914508 N chr2 129915294 N DEL 5
A00404:156:HV37TDSXX:2:2448:32434:36996 chr2 129914736 N chr2 129915409 N DEL 14
A00404:156:HV37TDSXX:1:2570:22155:15655 chr6 11936836 N chr6 11936967 N DUP 11
A00404:155:HV27LDSXX:4:1329:26386:5729 chr6 11936836 N chr6 11936967 N DUP 10
A00297:158:HT275DSXX:4:1469:3351:18912 chr6 11936884 N chr6 11936940 N DEL 15
A00404:156:HV37TDSXX:2:1352:22589:19601 chr14 97181459 N chr14 97181537 N DEL 6
A00404:156:HV37TDSXX:2:1130:22733:31438 chr3 14255507 N chr3 14255659 N DUP 1
A00404:155:HV27LDSXX:4:2653:2745:31140 chr3 14255548 N chr3 14255629 N DEL 3
A00404:156:HV37TDSXX:1:1676:9037:6809 chr17 307322 N chr17 307563 N DEL 5
A00297:158:HT275DSXX:3:2408:15185:34021 chr17 307405 N chr17 307470 N DEL 16
A00404:156:HV37TDSXX:2:2670:18891:20964 chr17 307405 N chr17 307470 N DEL 16
A00404:155:HV27LDSXX:2:2406:12717:4382 chr17 307405 N chr17 307470 N DEL 17
A00297:158:HT275DSXX:4:2171:9688:29356 chr17 307405 N chr17 307470 N DEL 20
A00404:155:HV27LDSXX:1:1320:1172:22561 chr17 307405 N chr17 307470 N DEL 20
A00297:158:HT275DSXX:3:1442:12491:18208 chr17 307405 N chr17 307470 N DEL 21
A00297:158:HT275DSXX:3:1177:6144:2487 chr17 307368 N chr17 307433 N DEL 25
A00404:156:HV37TDSXX:3:2335:5068:3662 chr17 307368 N chr17 307433 N DEL 25
A00297:158:HT275DSXX:1:2137:29984:8202 chr17 307368 N chr17 307433 N DEL 23
A00297:158:HT275DSXX:1:1426:17861:31172 chr17 307368 N chr17 307433 N DEL 25
A00404:155:HV27LDSXX:1:1343:23981:2785 chr17 307368 N chr17 307433 N DEL 25
A00404:155:HV27LDSXX:4:2114:9155:3912 chr17 307368 N chr17 307433 N DEL 19
A00404:156:HV37TDSXX:1:2347:4915:18897 chr17 307373 N chr17 307470 N DEL 6
A00404:155:HV27LDSXX:1:2347:29469:4272 chr17 307377 N chr17 307474 N DEL 2
A00404:156:HV37TDSXX:2:2168:25617:32550 chr17 307375 N chr17 307472 N DEL 4
A00404:156:HV37TDSXX:4:1437:10068:35650 chr17 307444 N chr17 307573 N DEL 18
A00404:156:HV37TDSXX:3:2606:29288:27978 chr4 19519947 N chr4 19520532 N DEL 3
A00404:155:HV27LDSXX:2:1650:25301:29653 chr4 19520537 N chr4 19520614 N DEL 17
A00297:158:HT275DSXX:1:2358:14968:6370 chr4 19520537 N chr4 19520614 N DEL 19
A00297:158:HT275DSXX:1:2457:22064:10676 chr4 19520506 N chr4 19520615 N DEL 5
A00404:155:HV27LDSXX:3:1407:1244:25160 chr4 19520506 N chr4 19520615 N DEL 5
A00297:158:HT275DSXX:3:1161:19623:6073 chr9 38628988 N chr9 38629151 N DEL 8
A00404:155:HV27LDSXX:1:1415:20555:17206 chr16 61768465 N chr16 61768554 N DUP 6
A00404:156:HV37TDSXX:3:1315:8133:33833 chr16 61768524 N chr16 61768581 N DUP 6
A00297:158:HT275DSXX:1:1633:23339:9408 chr16 61768476 N chr16 61768559 N DEL 4
A00404:156:HV37TDSXX:4:1465:21043:16016 chr2 239282314 N chr2 239282439 N DEL 4
A00297:158:HT275DSXX:3:2442:30671:11271 chr2 239282410 N chr2 239282493 N DUP 5
A00297:158:HT275DSXX:3:1161:10990:26882 chr4 109597707 N chr4 109598011 N DEL 23
A00297:158:HT275DSXX:2:2566:19831:2801 chr4 109597631 N chr4 109597854 N DUP 5
A00404:156:HV37TDSXX:2:2572:30960:22858 chr4 109597651 N chr4 109597922 N DUP 8
A00404:156:HV37TDSXX:2:2615:28908:31140 chr4 109597635 N chr4 109597761 N DUP 5
A00297:158:HT275DSXX:4:2309:4978:32597 chr4 109597635 N chr4 109597761 N DUP 5
A00404:156:HV37TDSXX:3:2125:8974:16501 chr4 109597630 N chr4 109597855 N DEL 8
A00404:156:HV37TDSXX:2:1211:32777:22247 chr9 136007493 N chr9 136007680 N DUP 4
A00404:156:HV37TDSXX:2:2635:26196:24095 chr9 136007493 N chr9 136007680 N DUP 6
A00404:155:HV27LDSXX:1:1177:23041:33567 chr9 136007493 N chr9 136007680 N DUP 7
A00404:156:HV37TDSXX:4:2306:11315:17487 chr9 136007565 N chr9 136007694 N DUP 7
A00297:158:HT275DSXX:2:2436:20907:9017 chr9 136007644 N chr9 136007715 N DEL 2
A00404:155:HV27LDSXX:4:1124:2546:21966 chr9 136007644 N chr9 136007715 N DEL 2
A00404:155:HV27LDSXX:4:2325:27778:20353 chr9 136007624 N chr9 136007709 N DEL 5
A00404:155:HV27LDSXX:4:1319:27841:26381 chr17 82218337 N chr17 82218614 N DEL 3
A00297:158:HT275DSXX:1:2645:11044:31986 chr17 82218352 N chr17 82218432 N DEL 10
A00404:155:HV27LDSXX:3:1405:5855:21652 chr17 82218371 N chr17 82218531 N DEL 11
A00404:156:HV37TDSXX:1:2173:6126:16861 chr17 82218374 N chr17 82218452 N DUP 1
A00404:155:HV27LDSXX:3:2246:26576:9377 chr17 82218374 N chr17 82218452 N DUP 3
A00404:155:HV27LDSXX:2:1633:14371:7874 chr17 82218374 N chr17 82218452 N DUP 4
A00404:156:HV37TDSXX:4:2202:4969:35556 chr17 82218374 N chr17 82218452 N DUP 5
A00404:155:HV27LDSXX:2:1114:1759:9518 chr17 82218374 N chr17 82218452 N DUP 11
A00404:155:HV27LDSXX:2:1361:17508:4225 chr17 82218522 N chr17 82218639 N DEL 14
A00404:156:HV37TDSXX:3:2542:18050:36824 chr17 82218374 N chr17 82218452 N DUP 11
A00297:158:HT275DSXX:2:2520:25111:17926 chr17 82218453 N chr17 82218531 N DUP 5
A00404:155:HV27LDSXX:1:2426:3794:8187 chr17 82218374 N chr17 82218452 N DUP 11
A00404:155:HV27LDSXX:2:1323:2736:25520 chr17 82218414 N chr17 82218613 N DEL 5
A00297:158:HT275DSXX:3:1272:30219:6699 chr1 52870075 N chr1 52870127 N DEL 38
A00404:155:HV27LDSXX:3:1234:1497:35618 chr16 78422840 N chr16 78422951 N DUP 10
A00404:156:HV37TDSXX:3:1404:12255:21590 chr16 78422840 N chr16 78422951 N DUP 10
A00404:156:HV37TDSXX:3:2250:10818:5572 chr16 78422889 N chr16 78422960 N DEL 9
A00297:158:HT275DSXX:3:1126:30382:30718 chr16 78422890 N chr16 78422961 N DEL 9
A00297:158:HT275DSXX:3:1126:31331:29575 chr16 78422890 N chr16 78422961 N DEL 9
A00404:155:HV27LDSXX:4:2410:29586:24424 chr16 78422845 N chr16 78423008 N DEL 3
A00404:155:HV27LDSXX:4:2346:11767:15608 chr16 78422844 N chr16 78423009 N DEL 4
A00297:158:HT275DSXX:4:1160:31150:11005 chr1 150729439 N chr1 150729711 N DEL 5
A00404:156:HV37TDSXX:2:1320:18168:10692 chr9 76064025 N chr9 76064427 N DEL 2
A00297:158:HT275DSXX:1:2418:20754:29230 chr9 76064071 N chr9 76064471 N DUP 1
A00404:155:HV27LDSXX:1:2347:17255:18630 chr9 76064092 N chr9 76064267 N DUP 5
A00297:158:HT275DSXX:1:2418:20754:29230 chr9 76064025 N chr9 76064425 N DUP 5
A00297:158:HT275DSXX:1:1352:17309:8923 chr9 76064349 N chr9 76064475 N DUP 5
A00297:158:HT275DSXX:4:2157:21893:32769 chr12 124622495 N chr12 124622570 N DEL 5
A00404:156:HV37TDSXX:3:1309:18295:15483 chr12 124622495 N chr12 124622570 N DEL 10
A00404:156:HV37TDSXX:4:2363:26585:34037 chr12 124622495 N chr12 124622570 N DEL 15
A00297:158:HT275DSXX:3:1144:25165:37059 chr10 54421831 N chr10 54422022 N DUP 7
A00297:158:HT275DSXX:2:1620:8151:13949 chr17 45417079 N chr17 45417389 N DEL 25
A00297:158:HT275DSXX:3:1418:18457:26663 chr17 45417902 N chr17 45418189 N DEL 2
A00404:155:HV27LDSXX:1:1204:7075:33661 chr1 9116317 N chr1 9116442 N DEL 2
A00404:155:HV27LDSXX:1:2643:26033:15796 chr1 9116317 N chr1 9116442 N DEL 5
A00404:156:HV37TDSXX:4:1606:20907:2942 chr1 9116282 N chr1 9116382 N DUP 1
A00404:155:HV27LDSXX:4:1208:12581:16391 chr1 9116282 N chr1 9116382 N DUP 1
A00297:158:HT275DSXX:3:1549:11261:28479 chr1 9116314 N chr1 9116470 N DUP 9
A00404:155:HV27LDSXX:4:2103:26485:14481 chr6 27826957 N chr6 27827537 N DEL 5
A00297:158:HT275DSXX:4:2650:16423:21386 chr6 27826957 N chr6 27827537 N DEL 5
A00404:156:HV37TDSXX:1:1201:21169:28479 chr6 27826949 N chr6 27827075 N DUP 4
A00297:158:HT275DSXX:1:2609:5177:18443 chr6 27826957 N chr6 27827360 N DEL 5
A00404:156:HV37TDSXX:1:1156:15609:11710 chr6 27826928 N chr6 27827057 N DEL 3
A00404:156:HV37TDSXX:2:2234:23348:14841 chr6 27827089 N chr6 27827313 N DUP 5
A00297:158:HT275DSXX:1:1230:8061:13103 chr6 27827094 N chr6 27827318 N DUP 5
A00297:158:HT275DSXX:2:2525:15998:29731 chr6 27827133 N chr6 27827360 N DEL 10
A00404:155:HV27LDSXX:1:2201:21233:33786 chr6 27826927 N chr6 27827104 N DEL 1
A00404:156:HV37TDSXX:4:1640:6650:2769 chr6 27826928 N chr6 27827106 N DEL 4
A00404:155:HV27LDSXX:4:1271:10682:31046 chr6 27827237 N chr6 27827415 N DEL 8
A00404:155:HV27LDSXX:4:1248:25789:10050 chr6 27827013 N chr6 27827237 N DUP 5
A00404:155:HV27LDSXX:4:1248:26738:6527 chr6 27827021 N chr6 27827245 N DUP 5
A00404:155:HV27LDSXX:1:1136:3956:14356 chr6 27827029 N chr6 27827609 N DEL 5
A00404:156:HV37TDSXX:2:2424:5981:1611 chr6 27827324 N chr6 27827502 N DEL 1
A00404:156:HV37TDSXX:2:2444:22697:5979 chr6 27826968 N chr6 27827369 N DUP 7
A00404:155:HV27LDSXX:3:2620:21585:22780 chr6 27827035 N chr6 27827360 N DEL 5
A00297:158:HT275DSXX:3:2434:22019:31516 chr6 27827183 N chr6 27827408 N DUP 5
A00297:158:HT275DSXX:1:2609:5177:18443 chr6 27827324 N chr6 27827500 N DUP 5
A00404:155:HV27LDSXX:2:2210:22896:8641 chr6 27826958 N chr6 27827536 N DUP 5
A00297:158:HT275DSXX:1:1650:8865:10770 chr6 27827123 N chr6 27827525 N DUP 5
A00297:158:HT275DSXX:2:2403:14624:32737 chr6 27826958 N chr6 27827536 N DUP 5
A00297:158:HT275DSXX:2:1302:16423:32690 chr6 27827255 N chr6 27827608 N DUP 1
A00404:156:HV37TDSXX:2:2654:18087:18693 chr6 27827136 N chr6 27827361 N DUP 5
A00297:158:HT275DSXX:4:1573:7464:5243 chr6 27826968 N chr6 27827548 N DEL 4
A00404:155:HV27LDSXX:4:1318:25211:9706 chr6 27827029 N chr6 27827609 N DEL 5
A00404:155:HV27LDSXX:4:1318:25346:9502 chr6 27827029 N chr6 27827609 N DEL 5
A00404:155:HV27LDSXX:3:1170:13123:10222 chr6 27827029 N chr6 27827609 N DEL 5
A00404:156:HV37TDSXX:2:2166:30382:29496 chr6 27827029 N chr6 27827609 N DEL 5
A00297:158:HT275DSXX:1:1650:8865:10770 chr6 27827029 N chr6 27827609 N DEL 5
A00404:155:HV27LDSXX:2:2218:21034:23202 chr6 27827029 N chr6 27827609 N DEL 5
A00404:155:HV27LDSXX:2:2218:25744:17049 chr6 27827029 N chr6 27827609 N DEL 5
A00404:156:HV37TDSXX:2:2477:13910:23077 chr6 27827029 N chr6 27827609 N DEL 5
A00297:158:HT275DSXX:2:2643:15944:34084 chr6 27827029 N chr6 27827609 N DEL 5
A00404:156:HV37TDSXX:3:2226:9227:19100 chr6 27827075 N chr6 27827655 N DEL 10
A00297:158:HT275DSXX:2:1223:28944:18333 chr6 27827029 N chr6 27827609 N DEL 5
A00404:155:HV27LDSXX:4:1248:25789:10050 chr6 27827075 N chr6 27827655 N DEL 10
A00404:155:HV27LDSXX:4:1248:26738:6527 chr6 27827075 N chr6 27827655 N DEL 10
A00297:158:HT275DSXX:4:1573:7464:5243 chr6 27826913 N chr6 27827620 N DEL 4
A00404:155:HV27LDSXX:3:1156:24306:31156 chr6 27827276 N chr6 27827680 N DEL 5
A00404:155:HV27LDSXX:2:2456:31548:21621 chr5 28232507 N chr5 28232597 N DUP 1
A00297:158:HT275DSXX:4:2308:30563:8328 chr8 100478568 N chr8 100478637 N DEL 1
A00404:156:HV37TDSXX:2:2342:5538:1094 chr4 156601329 N chr4 156601394 N DEL 1
A00404:156:HV37TDSXX:4:2512:11116:5713 chr4 156601244 N chr4 156601370 N DEL 5
A00404:156:HV37TDSXX:4:1313:21097:33301 chr4 156601247 N chr4 156601373 N DEL 5
A00404:155:HV27LDSXX:4:2665:3848:29731 chr4 156601499 N chr4 156601562 N DEL 10
A00404:155:HV27LDSXX:4:1556:13612:14325 chr11 76934811 N chr11 76934863 N DUP 12
A00404:155:HV27LDSXX:1:2611:3748:7012 chr11 76934811 N chr11 76934863 N DUP 16
A00404:155:HV27LDSXX:3:1135:19569:30091 chr11 76934825 N chr11 76934877 N DUP 1
A00297:158:HT275DSXX:4:1431:8929:15264 chr11 76934824 N chr11 76934876 N DUP 2
A00404:155:HV27LDSXX:2:1160:19117:23359 chr5 38862542 N chr5 38862787 N DEL 15
A00404:155:HV27LDSXX:2:1160:19117:23359 chr5 38862554 N chr5 38862799 N DEL 7
A00404:155:HV27LDSXX:4:1341:21278:1955 chr5 38862521 N chr5 38862842 N DEL 8
A00404:155:HV27LDSXX:1:1237:24786:32017 chr5 38862839 N chr5 38862920 N DEL 3
A00404:155:HV27LDSXX:3:2203:7021:32002 chr2 91443034 N chr2 91443116 N DEL 5
A00404:156:HV37TDSXX:2:1374:2727:30859 chr4 157248727 N chr4 157248844 N DUP 6
A00404:156:HV37TDSXX:3:1659:19325:28823 chrX 15736020 N chrX 15736325 N DEL 14
A00404:155:HV27LDSXX:2:1615:21187:2707 chrX 15736020 N chrX 15736325 N DEL 37
A00404:155:HV27LDSXX:1:1349:26982:9674 chr3 143086414 N chr3 143086543 N DEL 5
A00404:156:HV37TDSXX:3:2639:6940:20995 chr3 143086416 N chr3 143086799 N DEL 2
A00297:158:HT275DSXX:3:2101:27905:23359 chr3 143086398 N chr3 143086448 N DUP 7
A00404:155:HV27LDSXX:1:1245:10746:10770 chr3 143086544 N chr3 143086799 N DEL 10
A00297:158:HT275DSXX:3:2620:13693:3756 chr3 143086544 N chr3 143086799 N DEL 10
A00404:156:HV37TDSXX:2:1223:29695:27023 chr3 143086544 N chr3 143086799 N DEL 10
A00404:155:HV27LDSXX:2:2167:9534:12179 chr3 143086468 N chr3 143086594 N DUP 9
A00404:155:HV27LDSXX:4:2507:9643:22733 chr3 143086566 N chr3 143086821 N DEL 10
A00404:156:HV37TDSXX:1:1419:15962:30639 chr3 143086380 N chr3 143086481 N DEL 2
A00297:158:HT275DSXX:2:1175:22236:11412 chr3 143086381 N chr3 143086482 N DEL 1
A00404:156:HV37TDSXX:2:1665:30174:29074 chr3 143086381 N chr3 143086482 N DEL 1
A00404:155:HV27LDSXX:2:1602:10908:14873 chr3 143086602 N chr3 143086808 N DEL 2
A00404:155:HV27LDSXX:2:1602:11198:14372 chr3 143086602 N chr3 143086808 N DEL 2
A00404:155:HV27LDSXX:4:2222:13756:13698 chr3 143086533 N chr3 143086661 N DEL 4
A00297:158:HT275DSXX:1:1649:25762:17300 chr3 143086533 N chr3 143086661 N DEL 5
A00404:155:HV27LDSXX:1:2219:1931:24001 chr3 143086448 N chr3 143086574 N DUP 10
A00297:158:HT275DSXX:2:1213:21558:20635 chr3 143086468 N chr3 143086594 N DUP 2
A00404:156:HV37TDSXX:2:1647:14959:35227 chr3 143086468 N chr3 143086594 N DUP 10
A00404:155:HV27LDSXX:4:2245:11189:32550 chr3 143086468 N chr3 143086594 N DUP 10
A00404:155:HV27LDSXX:4:1649:8034:32910 chr3 143086641 N chr3 143086769 N DEL 5
A00404:156:HV37TDSXX:3:2269:12626:29496 chr2 177351090 N chr2 177351288 N DEL 3
A00404:156:HV37TDSXX:2:2278:28330:31172 chr2 177351104 N chr2 177351339 N DEL 7
A00404:156:HV37TDSXX:3:1642:29432:34428 chr2 177351200 N chr2 177351464 N DEL 10
A00404:156:HV37TDSXX:4:1471:8784:22247 chr17 81719335 N chr17 81719468 N DUP 1
A00404:156:HV37TDSXX:4:1524:20880:13510 chr17 17317098 N chr17 17317434 N DEL 25
A00404:156:HV37TDSXX:1:1677:15781:6026 chr17 17317098 N chr17 17317434 N DEL 5
A00404:155:HV27LDSXX:2:1570:8712:6183 chr17 17317098 N chr17 17317434 N DEL 5
A00404:156:HV37TDSXX:4:2260:15483:3787 chr17 17317098 N chr17 17317434 N DEL 5
A00297:158:HT275DSXX:4:1603:30608:28541 chr12 108363419 N chr12 108363502 N DUP 2
A00297:158:HT275DSXX:1:2205:30454:3693 chr12 108363479 N chr12 108363684 N DUP 5
A00404:155:HV27LDSXX:2:1357:17372:12665 chrX 147120656 N chrX 147120729 N DUP 15
A00404:156:HV37TDSXX:3:2660:11849:24674 chrX 147120666 N chrX 147120757 N DUP 13
A00404:156:HV37TDSXX:1:1401:11605:18709 chrX 147120677 N chrX 147120746 N DEL 18
A00404:156:HV37TDSXX:1:1401:11921:18255 chrX 147120677 N chrX 147120746 N DEL 18
A00404:155:HV27LDSXX:3:2136:23285:28635 chrX 147120677 N chrX 147120746 N DEL 18
A00404:156:HV37TDSXX:1:2631:8522:16094 chrX 147120677 N chrX 147120746 N DEL 16
A00297:158:HT275DSXX:1:1508:30120:5431 chrX 147120646 N chrX 147120750 N DEL 9
A00297:158:HT275DSXX:4:2315:3007:32002 chrX 147120642 N chrX 147120759 N DEL 2
A00297:158:HT275DSXX:2:2678:18882:1814 chr15 19822540 N chr15 19822722 N DUP 10
A00404:155:HV27LDSXX:2:2447:2636:14011 chr3 196207691 N chr3 196207788 N DUP 2
A00404:156:HV37TDSXX:3:1272:14425:36370 chr3 196207701 N chr3 196207799 N DEL 3
A00404:156:HV37TDSXX:1:2553:1154:32424 chr3 196207691 N chr3 196207788 N DUP 3
A00404:155:HV27LDSXX:4:1204:19135:10207 chr3 196207691 N chr3 196207788 N DUP 7
A00404:156:HV37TDSXX:4:2121:25129:11913 chr3 196207691 N chr3 196207788 N DUP 7
A00297:158:HT275DSXX:2:1506:14787:21371 chr3 196207701 N chr3 196207799 N DEL 7
A00297:158:HT275DSXX:3:1612:6786:24925 chr3 196207691 N chr3 196207788 N DUP 7
A00297:158:HT275DSXX:3:1351:15899:2096 chr3 196207736 N chr3 196207933 N DEL 11
A00404:155:HV27LDSXX:4:2543:22544:36965 chr3 196207736 N chr3 196207933 N DEL 11
A00404:155:HV27LDSXX:4:2543:22742:36996 chr3 196207736 N chr3 196207933 N DEL 11
A00404:155:HV27LDSXX:4:2645:2880:24831 chr3 196207736 N chr3 196207933 N DEL 6
A00404:155:HV27LDSXX:2:2660:17725:7858 chr3 196207744 N chr3 196207941 N DEL 6
A00404:156:HV37TDSXX:1:2527:22923:15702 chr16 28698022 N chr16 28698281 N DEL 5
A00404:156:HV37TDSXX:1:2171:7572:34648 chr16 28698014 N chr16 28698191 N DUP 5
A00404:156:HV37TDSXX:4:2356:18295:6370 chr16 28698044 N chr16 28698303 N DEL 3
A00404:156:HV37TDSXX:1:2141:2230:22764 chr16 28697941 N chr16 28697993 N DEL 8
A00404:156:HV37TDSXX:1:2141:2600:22999 chr16 28697941 N chr16 28697993 N DEL 8
A00404:156:HV37TDSXX:1:1670:13883:13792 chr16 28698090 N chr16 28698220 N DEL 5
A00404:155:HV27LDSXX:3:2226:14299:35994 chr16 28698167 N chr16 28698297 N DEL 5
A00404:155:HV27LDSXX:4:2246:7527:28902 chr16 28697962 N chr16 28698141 N DEL 14
A00297:158:HT275DSXX:4:2614:30933:8594 chr16 28698196 N chr16 28698324 N DUP 5
A00404:155:HV27LDSXX:3:1634:13105:25473 chr16 28698034 N chr16 28698164 N DEL 2
A00404:156:HV37TDSXX:2:2510:4906:8797 chr16 28698151 N chr16 28698280 N DEL 7
A00404:155:HV27LDSXX:2:1567:26078:16689 chr16 28698152 N chr16 28698280 N DEL 9
A00404:155:HV27LDSXX:2:2357:29288:4178 chr16 28697904 N chr16 28698339 N DUP 5
A00297:158:HT275DSXX:1:1509:30436:18850 chr16 28698277 N chr16 28698532 N DUP 3
A00404:155:HV27LDSXX:1:1168:29875:18599 chr16 28698158 N chr16 28698290 N DEL 7
A00404:155:HV27LDSXX:1:1357:3622:34068 chr16 28698262 N chr16 28698440 N DUP 5
A00404:155:HV27LDSXX:3:1419:5358:29058 chr16 28698421 N chr16 28698498 N DUP 5
A00404:156:HV37TDSXX:4:1276:15745:11945 chr7 155366117 N chr7 155366231 N DUP 5
A00297:158:HT275DSXX:4:1355:3540:26099 chr11 79124983 N chr11 79125044 N DEL 12
A00404:156:HV37TDSXX:3:1465:10267:24439 chr11 79124956 N chr11 79125049 N DEL 5
A00404:156:HV37TDSXX:3:1419:2672:25066 chr11 79124959 N chr11 79125052 N DEL 5
A00404:155:HV27LDSXX:4:1318:5782:31767 chr18 52302506 N chr18 52302662 N DUP 4
A00297:158:HT275DSXX:1:2525:28501:2284 chr10 67826769 N chr10 67826928 N DEL 4
A00297:158:HT275DSXX:2:1112:6316:8923 chr10 67826749 N chr10 67826946 N DUP 5
A00404:155:HV27LDSXX:1:1309:1732:25254 chr10 67826869 N chr10 67826946 N DUP 5
A00404:155:HV27LDSXX:1:1309:2121:25739 chr10 67826869 N chr10 67826946 N DUP 5
A00297:158:HT275DSXX:1:2152:26386:8422 chr10 67826742 N chr10 67826976 N DUP 3
A00404:156:HV37TDSXX:2:2612:24026:13667 chr10 67826752 N chr10 67826986 N DUP 3
A00404:156:HV37TDSXX:3:1609:31837:4366 chr10 67826748 N chr10 67826968 N DEL 1
A00297:158:HT275DSXX:3:2533:10321:6934 chr8 48148394 N chr8 48148735 N DUP 8
A00297:158:HT275DSXX:1:1503:4806:9157 chr8 48148539 N chr8 48148654 N DEL 3
A00404:156:HV37TDSXX:2:1133:2672:16924 chr8 48148550 N chr8 48148663 N DUP 5
A00404:155:HV27LDSXX:3:2455:15980:10598 chr8 48148551 N chr8 48148664 N DUP 4
A00404:155:HV27LDSXX:2:2276:24939:27993 chr8 48148387 N chr8 48148728 N DUP 5
A00297:158:HT275DSXX:1:2546:27398:31469 chr8 48148387 N chr8 48148728 N DUP 20
A00404:156:HV37TDSXX:2:2508:30183:27117 chr8 48148387 N chr8 48148728 N DUP 20
A00404:156:HV37TDSXX:2:2508:30192:27038 chr8 48148387 N chr8 48148728 N DUP 20
A00297:158:HT275DSXX:3:2563:29098:35509 chr8 48148387 N chr8 48148728 N DUP 53
A00404:156:HV37TDSXX:3:1426:29785:36667 chr8 48148387 N chr8 48148728 N DUP 54
A00404:156:HV37TDSXX:3:1364:4408:6809 chr10 112806678 N chr10 112806980 N DEL 5
A00404:156:HV37TDSXX:2:1422:3549:10895 chr8 77343888 N chr8 77344001 N DEL 5
A00297:158:HT275DSXX:1:2513:30092:34162 chr8 77343888 N chr8 77344001 N DEL 5
A00404:156:HV37TDSXX:3:1541:24352:7748 chr8 77343909 N chr8 77344024 N DUP 13
A00297:158:HT275DSXX:2:1221:26232:31485 chr8 77343913 N chr8 77344028 N DUP 11
A00404:155:HV27LDSXX:2:2105:17318:23469 chr8 77343917 N chr8 77344032 N DUP 7
A00404:155:HV27LDSXX:4:2451:17580:3004 chr8 77343891 N chr8 77344042 N DUP 9
A00297:158:HT275DSXX:2:2136:4399:12430 chr8 77343910 N chr8 77344003 N DEL 15
A00297:158:HT275DSXX:1:1350:8639:23719 chr8 77343923 N chr8 77344016 N DEL 2
A00404:156:HV37TDSXX:2:2273:30282:12446 chr8 77343815 N chr8 77344013 N DEL 5
A00404:156:HV37TDSXX:1:1374:19515:1626 chr8 77343892 N chr8 77344173 N DUP 10
A00404:155:HV27LDSXX:4:2649:19235:4805 chr8 77343891 N chr8 77344172 N DUP 11
A00404:155:HV27LDSXX:1:1656:13648:3208 chr8 77344003 N chr8 77344172 N DUP 12
A00404:155:HV27LDSXX:4:1160:27199:35603 chr8 77344003 N chr8 77344172 N DUP 13
A00404:155:HV27LDSXX:1:1454:20654:18035 chr8 77344077 N chr8 77344159 N DUP 17
A00404:156:HV37TDSXX:1:1234:27019:6136 chr8 77344077 N chr8 77344159 N DUP 15
A00404:155:HV27LDSXX:2:1176:17463:35900 chr8 77343869 N chr8 77344190 N DUP 12
A00404:156:HV37TDSXX:2:2645:30698:20400 chr8 77344057 N chr8 77344198 N DUP 14
A00404:156:HV37TDSXX:4:2668:32606:4570 chr8 77344057 N chr8 77344198 N DUP 24
A00404:156:HV37TDSXX:3:1342:11623:6339 chr8 77344023 N chr8 77344172 N DUP 23
A00404:155:HV27LDSXX:1:1178:16369:9111 chr8 77344057 N chr8 77344198 N DUP 31
A00404:155:HV27LDSXX:2:2105:17318:23469 chr8 77344023 N chr8 77344172 N DUP 26
A00404:155:HV27LDSXX:4:1572:19117:31720 chr8 77344057 N chr8 77344198 N DUP 32
A00404:156:HV37TDSXX:4:1573:2157:6856 chr8 77344023 N chr8 77344172 N DUP 29
A00404:155:HV27LDSXX:4:2645:15094:30326 chr8 77344033 N chr8 77344196 N DEL 18
A00297:158:HT275DSXX:2:1529:8784:26694 chr8 77344047 N chr8 77344190 N DEL 17
A00404:156:HV37TDSXX:2:1204:6126:35650 chr8 77344047 N chr8 77344190 N DEL 14
A00404:156:HV37TDSXX:3:2607:23583:31313 chr8 77344052 N chr8 77344195 N DEL 11
A00404:155:HV27LDSXX:2:2536:4616:36573 chr8 77344026 N chr8 77344189 N DEL 13
A00297:158:HT275DSXX:2:2272:30852:33661 chr8 77344029 N chr8 77344192 N DEL 12
A00404:155:HV27LDSXX:1:1448:1687:36918 chr8 77344031 N chr8 77344194 N DEL 10
A00404:155:HV27LDSXX:1:2237:11388:29731 chr8 77344034 N chr8 77344197 N DEL 7
A00404:155:HV27LDSXX:3:2257:5213:14528 chr8 77344078 N chr8 77344201 N DEL 3
A00404:156:HV37TDSXX:2:1603:2076:17018 chr8 77344077 N chr8 77344200 N DEL 4
A00404:156:HV37TDSXX:3:2627:20500:34115 chr16 34700156 N chr16 34700304 N DEL 2
A00404:156:HV37TDSXX:2:1669:20907:36354 chr2 1027418 N chr2 1027652 N DUP 5
A00404:156:HV37TDSXX:2:1676:15429:12085 chr3 189440542 N chr3 189440666 N DEL 18
A00404:155:HV27LDSXX:2:2543:24180:20541 chr3 189440588 N chr3 189440649 N DEL 17
A00297:158:HT275DSXX:4:2646:26675:16814 chr3 189440580 N chr3 189440639 N DEL 10
A00404:156:HV37TDSXX:3:2217:27887:18724 chr3 189440580 N chr3 189440639 N DEL 10
A00404:155:HV27LDSXX:3:1505:28411:13557 chr3 189440579 N chr3 189440638 N DEL 20
A00297:158:HT275DSXX:4:1341:30454:24799 chr22 17814894 N chr22 17815023 N DEL 3
A00297:158:HT275DSXX:3:2170:32199:29951 chr22 17814981 N chr22 17815108 N DUP 5
A00297:158:HT275DSXX:1:1335:7265:21997 chr22 17814915 N chr22 17814980 N DEL 5
A00297:158:HT275DSXX:1:1469:22336:5822 chr22 17815084 N chr22 17815147 N DUP 5
A00297:158:HT275DSXX:1:1453:32823:19695 chr22 17814916 N chr22 17815141 N DEL 5
A00404:155:HV27LDSXX:3:1357:8395:12148 chr6 83243648 N chr6 83243823 N DEL 3
A00297:158:HT275DSXX:1:2560:18521:2409 chr6 83243649 N chr6 83243706 N DUP 10
A00404:156:HV37TDSXX:3:2624:19895:15843 chr6 83243649 N chr6 83243706 N DUP 10
A00404:156:HV37TDSXX:4:1520:19190:21386 chr6 83243649 N chr6 83243706 N DUP 10
A00297:158:HT275DSXX:1:2325:13033:1892 chr6 83243649 N chr6 83243706 N DUP 10
A00404:156:HV37TDSXX:4:1668:29604:16564 chr6 83243698 N chr6 83243757 N DEL 10
A00404:156:HV37TDSXX:1:2540:31747:7842 chr6 83243736 N chr6 83243851 N DUP 10
A00404:156:HV37TDSXX:2:2459:17897:23531 chr6 83243698 N chr6 83243757 N DEL 10
A00297:158:HT275DSXX:2:2321:15619:23531 chr6 83243495 N chr6 83243736 N DEL 10
A00404:156:HV37TDSXX:4:2624:6361:8750 chr6 83243661 N chr6 83243749 N DEL 2
A00404:156:HV37TDSXX:4:2624:6488:8750 chr6 83243661 N chr6 83243749 N DEL 2
A00297:158:HT275DSXX:4:2556:22535:26710 chr6 83243765 N chr6 83243851 N DUP 10
A00297:158:HT275DSXX:2:2325:25400:9064 chr6 83243495 N chr6 83243765 N DEL 10
A00297:158:HT275DSXX:2:2223:4246:26569 chr6 83243495 N chr6 83243765 N DEL 10
A00404:156:HV37TDSXX:4:1618:30680:18333 chr6 83243768 N chr6 83243854 N DUP 9
A00297:158:HT275DSXX:3:2354:12274:5431 chr6 83243669 N chr6 83243786 N DEL 10
A00297:158:HT275DSXX:3:2104:11171:16391 chr6 83243659 N chr6 83243776 N DEL 4
A00404:156:HV37TDSXX:2:1323:26521:32831 chr6 83243728 N chr6 83243816 N DEL 3
A00404:155:HV27LDSXX:3:1305:10276:33223 chr6 83243656 N chr6 83243802 N DEL 5
A00404:156:HV37TDSXX:2:1448:16830:26475 chr6 83243659 N chr6 83243805 N DEL 4
A00297:158:HT275DSXX:3:2176:3739:29105 chr6 83243662 N chr6 83243837 N DEL 1
A00404:155:HV27LDSXX:1:1251:20943:3975 chr16 23169260 N chr16 23169348 N DEL 5
A00297:158:HT275DSXX:2:1409:18394:1157 chr3 57002577 N chr3 57002629 N DEL 18
A00297:158:HT275DSXX:2:1244:8006:18208 chr12 499482 N chr12 499827 N DEL 10
A00404:156:HV37TDSXX:4:1348:13874:26083 chr12 499550 N chr12 499743 N DEL 5
A00404:156:HV37TDSXX:2:1126:19732:22138 chr12 499530 N chr12 499763 N DEL 5
A00404:155:HV27LDSXX:1:1318:8992:35540 chr12 499702 N chr12 499855 N DEL 5
A00297:158:HT275DSXX:2:2112:12635:18521 chr11 8978400 N chr11 8978655 N DEL 10
A00297:158:HT275DSXX:2:2112:13286:14074 chr11 8978400 N chr11 8978655 N DEL 10
A00297:158:HT275DSXX:1:2207:23520:24095 chr11 8978506 N chr11 8978859 N DEL 1
A00404:156:HV37TDSXX:3:1224:12897:17033 chr11 8978418 N chr11 8978544 N DUP 1
A00404:155:HV27LDSXX:1:1556:27570:18239 chr11 8978506 N chr11 8978761 N DEL 1
A00297:158:HT275DSXX:4:1402:7726:7106 chr11 8978506 N chr11 8978761 N DEL 2
A00297:158:HT275DSXX:4:1402:8079:8531 chr11 8978506 N chr11 8978761 N DEL 2
A00404:156:HV37TDSXX:4:1428:26992:11851 chr11 8978506 N chr11 8978761 N DEL 2
A00404:155:HV27LDSXX:3:1146:24505:26396 chr11 8978461 N chr11 8978714 N DUP 1
A00404:155:HV27LDSXX:2:1217:9028:14340 chr11 8978517 N chr11 8978819 N DUP 2
A00404:156:HV37TDSXX:1:2462:5204:1955 chr11 8978445 N chr11 8978573 N DEL 1
A00297:158:HT275DSXX:2:2676:32814:25034 chr11 8978578 N chr11 8978704 N DUP 5
A00297:158:HT275DSXX:2:1317:30807:28729 chr11 8978582 N chr11 8978708 N DUP 5
A00297:158:HT275DSXX:2:1331:32090:36620 chr11 8978582 N chr11 8978708 N DUP 5
A00297:158:HT275DSXX:2:1317:30807:28729 chr11 8978588 N chr11 8978714 N DUP 1
A00297:158:HT275DSXX:2:1331:32090:36620 chr11 8978588 N chr11 8978714 N DUP 1
A00404:155:HV27LDSXX:3:1116:5891:27978 chr11 8978678 N chr11 8978952 N DUP 1
A00404:156:HV37TDSXX:4:2239:18421:18490 chr11 8978742 N chr11 8979066 N DEL 6
A00404:156:HV37TDSXX:1:1262:10881:36245 chr11 8978537 N chr11 8978743 N DEL 8
A00404:155:HV27LDSXX:3:2251:7473:2033 chr11 8978435 N chr11 8978768 N DEL 5
A00404:156:HV37TDSXX:2:2633:2338:5134 chr11 8978520 N chr11 8978775 N DEL 1
A00404:156:HV37TDSXX:2:1558:8422:36307 chr11 8978521 N chr11 8978923 N DEL 8
A00404:156:HV37TDSXX:3:2177:23927:30373 chr11 8978521 N chr11 8978923 N DEL 8
A00404:156:HV37TDSXX:3:1513:31295:16485 chr11 8978521 N chr11 8978923 N DEL 7
A00404:155:HV27LDSXX:1:1274:10158:22748 chr11 8978521 N chr11 8978923 N DEL 7
A00404:155:HV27LDSXX:1:2678:11921:21261 chr11 8978521 N chr11 8978923 N DEL 7
A00297:158:HT275DSXX:1:1508:20509:3255 chr11 8978772 N chr11 8979045 N DUP 10
A00297:158:HT275DSXX:1:2337:8341:36072 chr11 8978449 N chr11 8979103 N DUP 4
A00297:158:HT275DSXX:2:2205:24894:6339 chr11 8978555 N chr11 8979084 N DEL 10
A00404:155:HV27LDSXX:4:2351:19208:22795 chr11 8978462 N chr11 8979118 N DEL 1
A00404:155:HV27LDSXX:2:1409:29794:19930 chr5 174169799 N chr5 174169852 N DUP 25
A00297:158:HT275DSXX:2:2539:30816:26209 chr5 174169799 N chr5 174169852 N DUP 37
A00404:155:HV27LDSXX:1:2378:28456:17143 chr5 174169799 N chr5 174169852 N DUP 22
A00404:155:HV27LDSXX:3:1659:7120:16892 chr5 174169843 N chr5 174169920 N DUP 27
A00404:156:HV37TDSXX:1:1311:22236:12070 chr5 174169792 N chr5 174169845 N DUP 4
A00404:156:HV37TDSXX:3:2525:22580:14732 chr5 174169843 N chr5 174169920 N DUP 8
A00404:156:HV37TDSXX:4:2475:3712:1157 chr5 174169843 N chr5 174169920 N DUP 15
A00297:158:HT275DSXX:3:2311:27199:28213 chr5 174169834 N chr5 174169929 N DUP 26
A00404:155:HV27LDSXX:1:2554:8413:22388 chr5 174169834 N chr5 174169929 N DUP 29
A00404:155:HV27LDSXX:2:1220:14109:24674 chr5 174169853 N chr5 174169930 N DUP 21
A00404:155:HV27LDSXX:2:1220:14127:24674 chr5 174169853 N chr5 174169930 N DUP 21
A00297:158:HT275DSXX:3:2235:23511:1157 chr5 174169834 N chr5 174169929 N DUP 22
A00404:155:HV27LDSXX:1:1443:24496:8938 chr5 174169834 N chr5 174169929 N DUP 22
A00404:155:HV27LDSXX:1:1456:28158:4852 chr5 174169834 N chr5 174169929 N DUP 22
A00297:158:HT275DSXX:2:1520:31069:31939 chr5 174169845 N chr5 174169922 N DUP 22
A00404:156:HV37TDSXX:1:1240:23393:28291 chr5 174169797 N chr5 174169888 N DEL 16
A00404:156:HV37TDSXX:3:2216:8341:1783 chr5 174169840 N chr5 174169898 N DEL 5
A00404:156:HV37TDSXX:1:2557:29975:8563 chr1 1056702 N chr1 1056805 N DUP 1
A00404:156:HV37TDSXX:1:1264:24071:28808 chr1 1056702 N chr1 1056805 N DUP 4
A00297:158:HT275DSXX:2:1427:25744:13542 chr1 1056702 N chr1 1056805 N DUP 5
A00297:158:HT275DSXX:1:2273:18457:7968 chr1 1056701 N chr1 1056804 N DUP 5
A00404:155:HV27LDSXX:3:2512:16080:19507 chr1 1056702 N chr1 1056805 N DUP 7
A00404:156:HV37TDSXX:1:1269:6388:25770 chr1 1056702 N chr1 1056805 N DUP 8
A00404:156:HV37TDSXX:4:1545:18331:1141 chr1 1056761 N chr1 1056864 N DEL 14
A00404:155:HV27LDSXX:2:1548:5439:9064 chr1 1056761 N chr1 1056864 N DEL 5
A00404:155:HV27LDSXX:4:1478:31684:36010 chr1 1056761 N chr1 1056864 N DEL 5
A00297:158:HT275DSXX:1:1676:2356:4664 chr1 1056765 N chr1 1056868 N DEL 5
A00404:155:HV27LDSXX:1:1669:2465:11710 chr1 1056761 N chr1 1056864 N DEL 5
A00404:156:HV37TDSXX:4:2432:21468:21292 chr1 1056761 N chr1 1056864 N DEL 5
A00297:158:HT275DSXX:4:1606:29613:2112 chr1 1056761 N chr1 1056864 N DEL 5
A00404:155:HV27LDSXX:2:2425:13892:30718 chr1 1056761 N chr1 1056864 N DEL 5
A00404:155:HV27LDSXX:3:2512:16080:19507 chr1 1056733 N chr1 1056870 N DEL 5
A00404:155:HV27LDSXX:2:1565:10619:5979 chr1 1056735 N chr1 1056872 N DEL 5
A00404:155:HV27LDSXX:1:2135:2184:22748 chr1 1056685 N chr1 1056876 N DEL 3
A00404:155:HV27LDSXX:1:2135:3504:21746 chr1 1056685 N chr1 1056876 N DEL 3
A00297:158:HT275DSXX:1:2646:28022:9972 chr7 65489232 N chr7 65489394 N DUP 1
A00297:158:HT275DSXX:3:2332:19714:9486 chr7 65489229 N chr7 65489495 N DUP 6
A00404:155:HV27LDSXX:4:1674:24957:16250 chr7 65489197 N chr7 65489271 N DUP 7
A00297:158:HT275DSXX:4:1633:23610:25755 chr7 65489253 N chr7 65489311 N DUP 18
A00404:156:HV37TDSXX:4:2413:11957:35258 chr7 65489192 N chr7 65489292 N DUP 18
A00297:158:HT275DSXX:3:2154:18195:19852 chr7 65489192 N chr7 65489458 N DUP 12
A00297:158:HT275DSXX:2:2545:7355:8594 chr7 65489192 N chr7 65489292 N DUP 24
A00404:156:HV37TDSXX:4:2256:24695:29575 chr7 65489192 N chr7 65489292 N DUP 31
A00297:158:HT275DSXX:2:1166:28320:21856 chr7 65489268 N chr7 65489355 N DUP 5
A00297:158:HT275DSXX:2:2165:29107:22748 chr7 65489268 N chr7 65489355 N DUP 5
A00297:158:HT275DSXX:2:2161:32823:3223 chr7 65489269 N chr7 65489356 N DUP 5
A00404:155:HV27LDSXX:1:2433:11632:20823 chr7 65489275 N chr7 65489362 N DUP 3
A00404:156:HV37TDSXX:2:1643:21603:9095 chr7 65489288 N chr7 65489351 N DEL 16
A00404:156:HV37TDSXX:4:2116:7808:19085 chr11 64582052 N chr11 64582290 N DEL 3
A00404:155:HV27LDSXX:1:2557:5683:12900 chr11 64582210 N chr11 64582283 N DEL 8
A00404:156:HV37TDSXX:2:2261:25816:24815 chr11 64582202 N chr11 64582393 N DUP 18
A00404:156:HV37TDSXX:3:2318:3929:4445 chr11 64582286 N chr11 64582434 N DUP 36
A00404:155:HV27LDSXX:1:1350:21576:34851 chr11 64582215 N chr11 64582273 N DEL 1
A00404:155:HV27LDSXX:2:1229:18141:5635 chr11 64582262 N chr11 64582323 N DEL 15
A00404:155:HV27LDSXX:4:1472:1787:30201 chr11 64582286 N chr11 64582434 N DUP 10
A00297:158:HT275DSXX:2:1320:21495:32894 chr11 64582286 N chr11 64582434 N DUP 20
A00297:158:HT275DSXX:2:1320:21829:32784 chr11 64582286 N chr11 64582434 N DUP 20
A00404:155:HV27LDSXX:1:1463:23520:27571 chr11 64582286 N chr11 64582434 N DUP 20
A00404:155:HV27LDSXX:1:1463:23918:27132 chr11 64582286 N chr11 64582434 N DUP 20
A00404:155:HV27LDSXX:2:2430:5086:31657 chr11 64582286 N chr11 64582434 N DUP 20
A00404:155:HV27LDSXX:1:1345:20555:12696 chr11 64582263 N chr11 64582366 N DEL 14
A00297:158:HT275DSXX:3:2356:12861:9768 chr11 64582262 N chr11 64582427 N DEL 3
A00404:156:HV37TDSXX:3:1104:23647:27665 chr3 57119500 N chr3 57119678 N DEL 7
A00404:156:HV37TDSXX:1:2653:20790:15702 chr19 4638025 N chr19 4638203 N DEL 6
A00297:158:HT275DSXX:1:2423:23321:10379 chr20 4610592 N chr20 4610659 N DEL 5
A00404:155:HV27LDSXX:4:1376:5647:10614 chr20 4610555 N chr20 4610661 N DEL 5
A00404:155:HV27LDSXX:3:2413:5132:24721 chr1 230394776 N chr1 230394888 N DUP 5
A00404:155:HV27LDSXX:4:1473:27498:9126 chr1 230395692 N chr1 230395919 N DEL 3
A00404:155:HV27LDSXX:3:1641:2103:8046 chr1 230395813 N chr1 230395923 N DEL 29
A00404:156:HV37TDSXX:4:1254:12084:9392 chr15 40136112 N chr15 40136362 N DEL 4
A00404:155:HV27LDSXX:3:1622:5701:10582 chr15 40136407 N chr15 40136509 N DEL 10
A00297:158:HT275DSXX:1:2463:2329:2550 chr15 40136177 N chr15 40136424 N DUP 4
A00404:155:HV27LDSXX:3:1554:17987:6872 chr15 40136407 N chr15 40136605 N DEL 15
A00404:156:HV37TDSXX:1:1205:14208:14544 chr15 40136424 N chr15 40136526 N DEL 5
A00404:156:HV37TDSXX:1:1573:4354:34021 chr15 40136443 N chr15 40136593 N DEL 5
A00297:158:HT275DSXX:1:2345:26793:10347 chr15 40136142 N chr15 40136734 N DEL 4
A00404:156:HV37TDSXX:3:2522:4607:7122 chr10 6231885 N chr10 6232020 N DEL 2
A00297:158:HT275DSXX:3:2432:11605:22748 chr7 153329487 N chr7 153329622 N DEL 11
A00297:158:HT275DSXX:1:2678:30978:13213 chr7 153329527 N chr7 153329656 N DEL 9
A00297:158:HT275DSXX:2:1351:13376:28667 chr7 153329490 N chr7 153329625 N DEL 12
A00404:156:HV37TDSXX:1:2674:15727:31234 chr7 153329491 N chr7 153329626 N DEL 11
A00404:156:HV37TDSXX:2:2174:12635:5776 chr7 153329487 N chr7 153329626 N DEL 20
A00404:156:HV37TDSXX:1:1163:10474:16282 chr7 153329601 N chr7 153329667 N DEL 7
A00404:156:HV37TDSXX:3:1216:4354:10097 chr7 153329601 N chr7 153329667 N DEL 7
A00404:155:HV27LDSXX:4:2409:10881:1141 chr7 153329601 N chr7 153329667 N DEL 7
A00404:155:HV27LDSXX:4:2409:9679:1219 chr7 153329601 N chr7 153329667 N DEL 7
A00297:158:HT275DSXX:2:2154:26286:14700 chr11 91147292 N chr11 91147349 N DUP 13
A00297:158:HT275DSXX:2:1333:7591:32111 chrX 87234162 N chrX 87234239 N DEL 19
A00404:156:HV37TDSXX:1:1163:29206:24737 chrX 87234162 N chrX 87234239 N DEL 23
A00404:156:HV37TDSXX:1:1352:4634:25801 chrX 87234126 N chrX 87234239 N DEL 24
A00404:156:HV37TDSXX:1:1352:4960:25175 chrX 87234126 N chrX 87234239 N DEL 24
A00404:156:HV37TDSXX:1:1153:29315:16313 chrX 87234080 N chrX 87234332 N DUP 17
A00404:155:HV27LDSXX:3:1628:14443:33927 chrX 87233978 N chrX 87234253 N DEL 1
A00297:158:HT275DSXX:4:1558:16170:27117 chrX 87234093 N chrX 87234490 N DUP 18
A00404:156:HV37TDSXX:1:2555:16414:28416 chr10 133011041 N chr10 133011092 N DEL 54
A00404:155:HV27LDSXX:3:1541:23963:4163 chr10 133011073 N chr10 133011211 N DEL 28
A00404:155:HV27LDSXX:3:1121:9399:29105 chr10 133010969 N chr10 133011137 N DUP 9
A00404:155:HV27LDSXX:4:1472:18032:4225 chr10 133011148 N chr10 133011474 N DEL 11
A00297:158:HT275DSXX:2:1248:4029:32518 chr10 133011085 N chr10 133011341 N DUP 9
A00404:155:HV27LDSXX:4:2177:30427:7592 chr10 133011117 N chr10 133011643 N DUP 11
A00297:158:HT275DSXX:2:1351:1597:31000 chr10 133011074 N chr10 133011516 N DUP 5
A00404:155:HV27LDSXX:1:2219:23619:36104 chr10 133011085 N chr10 133011526 N DUP 11
A00297:158:HT275DSXX:1:2414:17662:6997 chr10 133011645 N chr10 133011782 N DUP 5
A00297:158:HT275DSXX:2:1552:18222:27383 chr10 133011081 N chr10 133011523 N DUP 5
A00404:156:HV37TDSXX:2:2231:18602:21872 chr10 133011081 N chr10 133011523 N DUP 5
A00297:158:HT275DSXX:2:1504:7726:7169 chr10 133011204 N chr10 133011254 N DUP 1
A00297:158:HT275DSXX:3:2561:6180:29606 chr10 133011128 N chr10 133011265 N DUP 18
A00404:156:HV37TDSXX:1:1236:26078:20384 chr10 133011069 N chr10 133011345 N DEL 23
A00404:156:HV37TDSXX:4:1165:24876:8907 chr10 133011228 N chr10 133011367 N DEL 24
A00297:158:HT275DSXX:2:1565:15347:2863 chr10 133011232 N chr10 133011371 N DEL 24
A00404:155:HV27LDSXX:4:1261:1325:33567 chr10 133011066 N chr10 133011342 N DEL 18
A00404:156:HV37TDSXX:3:2342:27434:5353 chr10 133011232 N chr10 133011371 N DEL 24
A00297:158:HT275DSXX:4:2558:12780:4648 chr10 133011128 N chr10 133011265 N DUP 13
A00404:155:HV27LDSXX:3:1541:23963:4163 chr10 133011073 N chr10 133011211 N DEL 14
A00404:155:HV27LDSXX:4:1246:22987:24486 chr10 133011228 N chr10 133011367 N DEL 24
A00404:156:HV37TDSXX:1:2125:23059:33004 chr10 133011263 N chr10 133011672 N DEL 18
A00297:158:HT275DSXX:2:2525:21477:5212 chr10 133011263 N chr10 133011672 N DEL 11
A00404:156:HV37TDSXX:4:2332:25672:34804 chr10 133011090 N chr10 133011331 N DUP 20
A00404:155:HV27LDSXX:1:2615:1127:16470 chr10 133011090 N chr10 133011739 N DUP 30
A00404:155:HV27LDSXX:4:1469:2528:10254 chr10 133011102 N chr10 133011275 N DEL 11
A00297:158:HT275DSXX:2:2360:18801:20744 chr10 133011169 N chr10 133011561 N DEL 17
A00404:156:HV37TDSXX:1:2218:18927:9878 chr10 133011088 N chr10 133011754 N DUP 12
A00297:158:HT275DSXX:3:2418:22733:34632 chr10 133011085 N chr10 133011341 N DUP 7
A00404:155:HV27LDSXX:4:2177:30427:7592 chr10 133011372 N chr10 133011475 N DUP 15
A00297:158:HT275DSXX:2:1306:24388:26443 chr10 133011374 N chr10 133011475 N DUP 22
A00404:155:HV27LDSXX:1:2412:19542:36808 chr10 133011347 N chr10 133011601 N DUP 25
A00404:156:HV37TDSXX:4:2323:22444:11240 chr10 133011077 N chr10 133011351 N DEL 20
A00404:156:HV37TDSXX:2:1157:27624:16172 chr10 133011495 N chr10 133011683 N DEL 12
A00297:158:HT275DSXX:3:1330:6361:8406 chr10 133011378 N chr10 133011598 N DUP 27
A00297:158:HT275DSXX:2:2563:14922:4539 chr10 133011070 N chr10 133011344 N DEL 20
A00404:156:HV37TDSXX:2:2505:25400:19742 chr10 133011042 N chr10 133011877 N DUP 7
A00297:158:HT275DSXX:3:2561:6180:29606 chr10 133011495 N chr10 133011683 N DEL 13
A00404:156:HV37TDSXX:3:2158:25961:8594 chr10 133011438 N chr10 133011505 N DEL 12
A00297:158:HT275DSXX:1:2414:17662:6997 chr10 133011257 N chr10 133011685 N DEL 10
A00404:156:HV37TDSXX:4:2332:25672:34804 chr10 133011495 N chr10 133011683 N DEL 22
A00297:158:HT275DSXX:2:2152:29107:29888 chr10 133011485 N chr10 133011877 N DUP 21
A00404:156:HV37TDSXX:1:1464:19090:6840 chr10 133011682 N chr10 133011853 N DUP 2
A00404:155:HV27LDSXX:2:1311:31584:7623 chr10 133011485 N chr10 133011877 N DUP 22
A00404:156:HV37TDSXX:4:1337:19235:11819 chr10 133011485 N chr10 133011877 N DUP 29
A00404:155:HV27LDSXX:1:1641:6732:33442 chr10 133011143 N chr10 133011552 N DEL 22
A00404:156:HV37TDSXX:4:2262:2700:15248 chr10 133011180 N chr10 133011349 N DEL 41
A00404:155:HV27LDSXX:4:2246:29423:17785 chr10 133011180 N chr10 133011349 N DEL 26
A00404:155:HV27LDSXX:1:1641:6732:33442 chr10 133011180 N chr10 133011349 N DEL 20
A00404:155:HV27LDSXX:3:2374:10321:35086 chr10 133011180 N chr10 133011349 N DEL 20
A00404:155:HV27LDSXX:2:1670:6786:1971 chr10 133011180 N chr10 133011349 N DEL 16
A00297:158:HT275DSXX:2:1331:18457:3834 chr10 133011041 N chr10 133011621 N DEL 5
A00297:158:HT275DSXX:3:1451:16785:20885 chr10 133011476 N chr10 133011698 N DUP 25
A00297:158:HT275DSXX:1:1238:4625:26537 chr10 133011415 N chr10 133011484 N DEL 32
A00404:155:HV27LDSXX:1:1471:17589:28009 chr10 133011152 N chr10 133011476 N DEL 18
A00404:155:HV27LDSXX:3:2148:20030:11099 chr10 133011416 N chr10 133011485 N DEL 25
A00404:155:HV27LDSXX:2:1124:16170:1783 chr10 133011178 N chr10 133011485 N DEL 14
A00404:156:HV37TDSXX:1:1352:11388:33802 chr10 133011471 N chr10 133011521 N DUP 13
A00297:158:HT275DSXX:1:1521:32560:16548 chr10 133011141 N chr10 133011618 N DUP 10
A00404:155:HV27LDSXX:1:1602:8043:10003 chr10 133011090 N chr10 133011601 N DUP 27
A00297:158:HT275DSXX:3:1241:8965:13197 chr10 133011703 N chr10 133011787 N DUP 7
A00297:158:HT275DSXX:4:1363:21567:2801 chr10 133011347 N chr10 133011601 N DUP 36
A00404:155:HV27LDSXX:4:2235:27597:21512 chr10 133011347 N chr10 133011601 N DUP 35
A00297:158:HT275DSXX:1:1602:19316:23923 chr10 133011117 N chr10 133011781 N DUP 17
A00297:158:HT275DSXX:3:2172:20320:36839 chr10 133011117 N chr10 133011643 N DUP 11
A00297:158:HT275DSXX:3:2418:22733:34632 chr10 133011085 N chr10 133011751 N DUP 11
A00404:155:HV27LDSXX:4:1656:10619:19100 chr10 133011110 N chr10 133011776 N DUP 10
A00404:156:HV37TDSXX:2:1315:10158:1360 chr10 133011516 N chr10 133011791 N DEL 8
A00404:156:HV37TDSXX:2:1134:2383:7874 chr10 133011516 N chr10 133011791 N DEL 7
A00297:158:HT275DSXX:3:1316:2618:5055 chr10 133011117 N chr10 133011643 N DUP 11
A00297:158:HT275DSXX:3:1647:27326:15280 chr10 133011085 N chr10 133011528 N DUP 9
A00404:156:HV37TDSXX:3:1272:24099:23187 chr10 133011645 N chr10 133011782 N DUP 5
A00404:155:HV27LDSXX:2:1414:6587:6511 chr10 133011645 N chr10 133011782 N DUP 5
A00297:158:HT275DSXX:2:1310:6795:2018 chr10 133011117 N chr10 133011643 N DUP 11
A00297:158:HT275DSXX:4:2601:21775:2503 chr10 133011135 N chr10 133011797 N DUP 17
A00404:155:HV27LDSXX:4:2354:32723:23093 chr10 133011645 N chr10 133011782 N DUP 5
A00404:155:HV27LDSXX:1:1557:30436:22294 chr10 133011645 N chr10 133011782 N DUP 5
A00404:155:HV27LDSXX:3:2663:9552:5822 chr10 133011117 N chr10 133011643 N DUP 11
A00404:155:HV27LDSXX:2:2157:17716:3865 chr10 133011151 N chr10 133011727 N DUP 9
A00297:158:HT275DSXX:4:1344:22724:35900 chr10 133011092 N chr10 133011707 N DUP 4
A00297:158:HT275DSXX:2:1478:16034:2801 chr10 133011645 N chr10 133011833 N DUP 9
A00297:158:HT275DSXX:4:2211:27814:4319 chr10 133011096 N chr10 133011711 N DUP 7
A00404:155:HV27LDSXX:3:2663:9552:5822 chr10 133011092 N chr10 133011707 N DUP 5
A00404:155:HV27LDSXX:1:1432:20934:7279 chr10 133011645 N chr10 133011782 N DUP 5
A00404:155:HV27LDSXX:1:1471:17589:28009 chr10 133011485 N chr10 133011877 N DUP 32
A00404:156:HV37TDSXX:1:2541:3595:8437 chr10 133011485 N chr10 133011877 N DUP 34
A00297:158:HT275DSXX:4:1450:30427:34209 chr10 133011151 N chr10 133011742 N DUP 14
A00404:156:HV37TDSXX:1:1464:19090:6840 chr10 133011528 N chr10 133011631 N DEL 3
A00404:155:HV27LDSXX:3:2624:2709:19241 chr10 133011416 N chr10 133011485 N DEL 37
A00404:155:HV27LDSXX:4:1210:19886:26882 chr10 133011663 N chr10 133011744 N DUP 13
A00404:155:HV27LDSXX:4:1210:20374:27978 chr10 133011476 N chr10 133011887 N DUP 10
A00404:155:HV27LDSXX:4:2246:29423:17785 chr10 133011663 N chr10 133011744 N DUP 13
A00404:155:HV27LDSXX:4:2235:27597:21512 chr10 133011150 N chr10 133011561 N DEL 25
A00404:155:HV27LDSXX:2:1542:23927:31438 chr10 133011508 N chr10 133011723 N DUP 15
A00404:156:HV37TDSXX:3:2417:7871:12962 chr10 133011663 N chr10 133011744 N DUP 19
A00297:158:HT275DSXX:3:2357:4951:12978 chr10 133011217 N chr10 133011527 N DEL 20
A00404:156:HV37TDSXX:1:2374:28438:35524 chr10 133011476 N chr10 133011887 N DUP 13
A00404:156:HV37TDSXX:3:2412:6488:6684 chr10 133011476 N chr10 133011698 N DUP 21
A00404:155:HV27LDSXX:2:2157:17716:3865 chr10 133011133 N chr10 133011680 N DEL 9
A00404:156:HV37TDSXX:3:2211:22299:21355 chr10 133011158 N chr10 133011705 N DEL 5
A00404:156:HV37TDSXX:2:1266:15185:7122 chr10 133011032 N chr10 133011699 N DEL 6
A00404:156:HV37TDSXX:2:1315:10158:1360 chr10 133011643 N chr10 133011784 N DEL 7
A00297:158:HT275DSXX:3:2469:30915:26506 chr10 133011643 N chr10 133011784 N DEL 7
A00297:158:HT275DSXX:2:2571:26558:2237 chr10 133011643 N chr10 133011784 N DEL 7
A00297:158:HT275DSXX:2:2360:18801:20744 chr10 133011643 N chr10 133011784 N DEL 7
A00297:158:HT275DSXX:4:2355:10673:3975 chr10 133011643 N chr10 133011784 N DEL 7
A00404:156:HV37TDSXX:1:2541:3595:8437 chr10 133011574 N chr10 133011801 N DEL 8
A00404:156:HV37TDSXX:2:2410:21775:7889 chr10 133011524 N chr10 133011757 N DEL 11
A00404:156:HV37TDSXX:4:2262:2700:15248 chr10 133010984 N chr10 133011562 N DEL 11
A00297:158:HT275DSXX:4:2509:32009:8923 chr10 133010874 N chr10 133011945 N DUP 5
A00297:158:HT275DSXX:4:1325:18304:35446 chr10 133010985 N chr10 133011854 N DEL 7
A00404:155:HV27LDSXX:4:2667:14317:21026 chr12 124339377 N chr12 124339558 N DUP 8
A00404:156:HV37TDSXX:3:2552:14561:29872 chr12 124339285 N chr12 124339384 N DEL 5
A00297:158:HT275DSXX:4:1670:11993:36417 chr3 97328048 N chr3 97328105 N DEL 7
A00404:155:HV27LDSXX:2:2416:27633:7513 chr3 97328048 N chr3 97328105 N DEL 31
A00404:155:HV27LDSXX:3:2632:22372:21073 chr3 97328048 N chr3 97328105 N DEL 29
A00404:155:HV27LDSXX:4:2320:25192:5541 chr11 63572243 N chr11 63572328 N DEL 1
A00404:156:HV37TDSXX:1:1261:8332:1955 chr11 44978537 N chr11 44978708 N DEL 10
A00297:158:HT275DSXX:2:1160:14290:36980 chr11 2773261 N chr11 2773406 N DUP 5
A00297:158:HT275DSXX:2:2160:12038:12978 chr11 2773261 N chr11 2773406 N DUP 5
A00404:156:HV37TDSXX:1:1237:32777:8782 chr11 2773342 N chr11 2773476 N DEL 39
A00404:156:HV37TDSXX:1:1504:12590:3662 chr11 2773610 N chr11 2773802 N DUP 1
A00404:156:HV37TDSXX:1:1171:20256:7263 chr2 236707124 N chr2 236707223 N DEL 16
A00404:155:HV27LDSXX:4:1632:20844:23970 chr2 236707331 N chr2 236707424 N DEL 1
A00404:156:HV37TDSXX:3:1305:9697:3067 chr2 236707082 N chr2 236707381 N DEL 38
A00404:156:HV37TDSXX:3:2260:21856:29794 chr9 135927972 N chr9 135928135 N DEL 21
A00404:156:HV37TDSXX:2:2545:9173:36260 chr9 135927848 N chr9 135928157 N DEL 13
A00297:158:HT275DSXX:4:2156:13648:31297 chr9 135928075 N chr9 135928179 N DEL 15
A00404:155:HV27LDSXX:1:1368:11225:34710 chr15 24120137 N chr15 24120200 N DEL 5
A00297:158:HT275DSXX:2:2513:14353:14794 chr15 24120139 N chr15 24120202 N DEL 5
A00297:158:HT275DSXX:2:1633:16595:10316 chr9 404053 N chr9 404144 N DEL 7
A00404:155:HV27LDSXX:2:1525:16306:15358 chr9 404053 N chr9 404144 N DEL 13
A00404:155:HV27LDSXX:3:1331:20799:33098 chr9 404056 N chr9 404151 N DEL 8
A00297:158:HT275DSXX:2:1270:21133:25191 chr9 404053 N chr9 404144 N DEL 18
A00404:155:HV27LDSXX:1:2262:7681:10629 chr9 404057 N chr9 404158 N DEL 1
A00404:155:HV27LDSXX:1:1275:14253:26396 chr4 7657449 N chr4 7657634 N DUP 3
A00404:156:HV37TDSXX:3:1637:20066:16360 chr4 7657495 N chr4 7657640 N DUP 6
A00404:156:HV37TDSXX:4:2539:15456:33144 chr4 7657495 N chr4 7657640 N DUP 7
A00404:156:HV37TDSXX:2:1364:28275:15358 chr4 7657495 N chr4 7657640 N DUP 7
A00404:156:HV37TDSXX:1:1638:15176:5384 chr2 78593354 N chr2 78593495 N DEL 13
A00404:156:HV37TDSXX:1:2638:15076:12633 chr2 78593354 N chr2 78593495 N DEL 13
A00297:158:HT275DSXX:1:1657:17155:2487 chr2 78593359 N chr2 78593500 N DEL 5
A00404:156:HV37TDSXX:4:2575:14904:32878 chr2 78593354 N chr2 78593495 N DEL 7
A00404:155:HV27LDSXX:4:2272:18982:9314 chr2 78593363 N chr2 78593504 N DEL 5
A00297:158:HT275DSXX:3:2509:30779:19507 chr1 3181239 N chr1 3181410 N DUP 25
A00404:155:HV27LDSXX:2:2550:15176:9204 chr1 3181239 N chr1 3181410 N DUP 25
A00404:155:HV27LDSXX:3:1549:5113:11162 chr1 3181241 N chr1 3181412 N DUP 25
A00297:158:HT275DSXX:4:2533:32660:18380 chr1 3181286 N chr1 3181495 N DUP 18
A00404:155:HV27LDSXX:3:1151:11397:10989 chr1 3181286 N chr1 3181495 N DUP 10
A00404:156:HV37TDSXX:2:1110:24044:23876 chr1 3181319 N chr1 3181402 N DUP 19
A00404:155:HV27LDSXX:3:1549:21884:32158 chr1 3181319 N chr1 3181402 N DUP 19
A00404:155:HV27LDSXX:2:1369:11586:13322 chr1 3181319 N chr1 3181390 N DUP 23
A00297:158:HT275DSXX:4:1608:28013:36104 chr1 3181392 N chr1 3181443 N DUP 9
A00297:158:HT275DSXX:1:2519:22128:25128 chr1 3181406 N chr1 3181507 N DUP 25
A00404:155:HV27LDSXX:4:1259:29821:15937 chr1 3181349 N chr1 3181490 N DUP 1
A00297:158:HT275DSXX:2:2339:5240:23813 chr1 3181406 N chr1 3181507 N DUP 21
A00404:155:HV27LDSXX:1:1444:31168:14137 chr1 3181368 N chr1 3181495 N DUP 11
A00404:156:HV37TDSXX:2:1172:23430:24878 chr1 3181367 N chr1 3181482 N DUP 1
A00404:155:HV27LDSXX:2:1506:32344:1642 chr2 60056669 N chr2 60056820 N DEL 5
A00297:158:HT275DSXX:1:2667:2410:17597 chr8 141658335 N chr8 141658495 N DEL 1
A00404:155:HV27LDSXX:4:1549:2003:33426 chr8 141658352 N chr8 141658506 N DEL 24
A00404:155:HV27LDSXX:4:1549:2013:33411 chr8 141658352 N chr8 141658506 N DEL 24
A00404:155:HV27LDSXX:4:1111:28556:17816 chr8 141658352 N chr8 141658506 N DEL 26
A00297:158:HT275DSXX:1:2605:30581:2096 chr8 141658400 N chr8 141658485 N DEL 16
A00404:155:HV27LDSXX:1:2242:25129:7373 chr8 141658400 N chr8 141658485 N DEL 19
A00404:155:HV27LDSXX:2:2242:11731:23375 chr8 141658365 N chr8 141658564 N DEL 7
A00297:158:HT275DSXX:2:2550:26124:13166 chr16 2802216 N chr16 2802374 N DEL 5
A00297:158:HT275DSXX:2:1252:3341:13949 chr16 2802207 N chr16 2802597 N DEL 7
A00297:158:HT275DSXX:4:1518:22643:4570 chr16 2802122 N chr16 2802173 N DEL 15
A00404:155:HV27LDSXX:3:1208:26087:33176 chr16 2802263 N chr16 2802535 N DUP 5
A00404:156:HV37TDSXX:1:2206:20518:35086 chr11 124166316 N chr11 124166369 N DEL 26
A00404:156:HV37TDSXX:1:2613:13991:16830 chr11 124166321 N chr11 124166374 N DEL 25
A00404:155:HV27LDSXX:2:1113:29595:20932 chr11 124166316 N chr11 124166369 N DEL 25
A00297:158:HT275DSXX:3:2123:25464:30029 chr11 124166316 N chr11 124166369 N DEL 18
A00297:158:HT275DSXX:3:2564:21097:11631 chr11 124166320 N chr11 124166373 N DEL 11
A00404:156:HV37TDSXX:1:2373:19126:35055 chr9 103014827 N chr9 103014933 N DEL 5
A00404:156:HV37TDSXX:3:1265:27254:28307 chr9 103014827 N chr9 103014933 N DEL 5
A00404:156:HV37TDSXX:4:1671:21875:23093 chr9 103014827 N chr9 103014933 N DEL 21
A00404:155:HV27LDSXX:1:1530:14353:5995 chr9 103014827 N chr9 103014933 N DEL 16
A00404:155:HV27LDSXX:3:2510:9507:13448 chr9 103014703 N chr9 103014934 N DEL 5
A00404:156:HV37TDSXX:2:1231:12961:11381 chr9 103014703 N chr9 103014934 N DEL 5
A00297:158:HT275DSXX:3:2629:25554:3411 chr9 103014706 N chr9 103014937 N DEL 5
A00297:158:HT275DSXX:4:2152:19506:12602 chr9 103014706 N chr9 103014937 N DEL 5
A00297:158:HT275DSXX:3:2446:4218:19194 chr9 103014709 N chr9 103014940 N DEL 5
A00404:155:HV27LDSXX:1:1125:32615:29543 chr9 103014709 N chr9 103014940 N DEL 5
A00404:155:HV27LDSXX:1:1126:30427:1016 chr9 103014709 N chr9 103014940 N DEL 5
A00404:155:HV27LDSXX:3:2510:9507:13448 chr9 103015227 N chr9 103015303 N DEL 3
A00297:158:HT275DSXX:1:2365:10185:25488 chr9 103015227 N chr9 103015303 N DEL 4
A00404:155:HV27LDSXX:3:1257:21504:28463 chr9 103015227 N chr9 103015303 N DEL 4
A00404:155:HV27LDSXX:4:2250:10122:15139 chr6 67407645 N chr6 67407708 N DEL 12
A00404:155:HV27LDSXX:1:1348:21386:8061 chr10 68182406 N chr10 68182513 N DUP 7
A00404:155:HV27LDSXX:1:1359:29604:25895 chr10 68182397 N chr10 68182456 N DEL 7
A00404:155:HV27LDSXX:1:1647:21043:36119 chr10 68182397 N chr10 68182456 N DEL 7
A00404:156:HV37TDSXX:4:2147:16667:35650 chr10 68182397 N chr10 68182456 N DEL 7
A00404:155:HV27LDSXX:1:1318:28194:31876 chr10 68182409 N chr10 68182468 N DEL 3
A00297:158:HT275DSXX:1:2344:14217:26490 chr10 68182376 N chr10 68182603 N DUP 7
A00297:158:HT275DSXX:2:2507:2067:34757 chr10 68182364 N chr10 68182567 N DUP 2
A00404:156:HV37TDSXX:4:1549:26015:18145 chr10 68182364 N chr10 68182567 N DUP 2
A00404:155:HV27LDSXX:1:1134:12183:13385 chr10 68182376 N chr10 68182603 N DUP 6
A00404:156:HV37TDSXX:1:2276:5665:36385 chr5 169290049 N chr5 169290122 N DEL 5
A00404:156:HV37TDSXX:2:1454:23900:23437 chr5 169290049 N chr5 169290122 N DEL 5
A00404:156:HV37TDSXX:4:2166:11695:17957 chr5 169290306 N chr5 169290379 N DEL 52
A00404:156:HV37TDSXX:2:2261:25220:2018 chr5 169290357 N chr5 169290465 N DUP 7
A00404:156:HV37TDSXX:4:2266:14271:22169 chr5 169290465 N chr5 169290932 N DEL 7
A00404:156:HV37TDSXX:1:2320:27516:35462 chr5 169290465 N chr5 169290932 N DEL 7
A00404:156:HV37TDSXX:1:1260:12789:13651 chr5 169290465 N chr5 169290932 N DEL 7
A00297:158:HT275DSXX:2:2523:2121:17127 chr5 169290520 N chr5 169290605 N DEL 2
A00404:156:HV37TDSXX:3:1446:31186:27258 chr5 169290150 N chr5 169290523 N DEL 51
A00404:156:HV37TDSXX:2:1204:26693:32628 chr5 169290126 N chr5 169290547 N DEL 25
A00404:155:HV27LDSXX:1:1256:1099:22780 chr5 169290605 N chr5 169290736 N DUP 5
A00404:155:HV27LDSXX:4:2220:26142:26443 chr5 169290302 N chr5 169290780 N DUP 4
A00297:158:HT275DSXX:1:2524:5086:14278 chr5 169290391 N chr5 169291051 N DEL 5
A00404:155:HV27LDSXX:4:2232:11424:35023 chr7 70845747 N chr7 70845806 N DEL 13
A00404:155:HV27LDSXX:3:1123:28528:15671 chr3 13682219 N chr3 13682282 N DUP 7
A00404:156:HV37TDSXX:2:2539:30906:24455 chr3 13682228 N chr3 13682297 N DUP 12
A00404:155:HV27LDSXX:1:2652:7717:27915 chr3 13682228 N chr3 13682297 N DUP 12
A00404:156:HV37TDSXX:1:2359:13593:18427 chr1 6107137 N chr1 6108038 N DUP 1
A00297:158:HT275DSXX:3:2277:17481:14262 chr1 6107376 N chr1 6107678 N DEL 5
A00404:155:HV27LDSXX:3:2435:11080:24659 chr1 6107951 N chr1 6108049 N DUP 5
A00404:155:HV27LDSXX:2:2469:19642:15937 chr1 6107432 N chr1 6108331 N DEL 5
A00297:158:HT275DSXX:3:1263:28221:20838 chr1 6108055 N chr1 6108355 N DEL 3
A00297:158:HT275DSXX:3:1407:12915:19006 chr1 6107199 N chr1 6108357 N DEL 6
A00404:155:HV27LDSXX:4:1110:7979:23923 chr11 67984167 N chr11 67984316 N DEL 15
A00404:156:HV37TDSXX:1:1277:14009:25786 chrX 6532894 N chrX 6532966 N DEL 19
A00404:156:HV37TDSXX:4:2332:10068:24001 chrX 6532913 N chrX 6532977 N DEL 13
A00297:158:HT275DSXX:3:1656:20916:11600 chrX 6532941 N chrX 6532995 N DUP 6
A00297:158:HT275DSXX:2:1319:18466:1752 chrX 6533023 N chrX 6533298 N DEL 16
A00297:158:HT275DSXX:4:2570:6705:2988 chrX 6533057 N chrX 6533115 N DUP 4
A00404:156:HV37TDSXX:4:1558:17210:27414 chrX 6533081 N chrX 6533517 N DEL 9
A00297:158:HT275DSXX:3:2111:14751:9752 chrX 6532870 N chrX 6533431 N DUP 28
A00404:156:HV37TDSXX:2:1542:18954:27117 chrX 6533089 N chrX 6533500 N DEL 17
A00297:158:HT275DSXX:2:1473:15004:3897 chrX 6532983 N chrX 6533637 N DEL 5
A00404:155:HV27LDSXX:4:1354:32597:25003 chr16 34713844 N chr16 34714143 N DUP 5
A00297:158:HT275DSXX:3:1155:13440:8171 chr16 34713998 N chr16 34714170 N DUP 4
A00297:158:HT275DSXX:3:1155:13810:7874 chr16 34713998 N chr16 34714170 N DUP 4
A00297:158:HT275DSXX:3:2157:12400:11725 chr16 34713998 N chr16 34714170 N DUP 4
A00297:158:HT275DSXX:3:2229:15402:21559 chr16 34713998 N chr16 34714170 N DUP 4
A00297:158:HT275DSXX:3:1622:24379:6417 chr16 34713953 N chr16 34714125 N DUP 5
A00404:156:HV37TDSXX:1:1309:5258:28855 chr16 34713953 N chr16 34714125 N DUP 5
A00404:156:HV37TDSXX:1:1611:31910:29199 chr16 34713953 N chr16 34714125 N DUP 5
A00404:155:HV27LDSXX:4:2508:28718:24893 chr16 34713953 N chr16 34714125 N DUP 5
A00404:156:HV37TDSXX:3:2168:21504:36198 chr16 34713953 N chr16 34714125 N DUP 5
A00404:155:HV27LDSXX:4:1273:23439:3912 chr16 34714054 N chr16 34714125 N DUP 5
A00404:155:HV27LDSXX:4:2204:6081:30499 chr16 34714054 N chr16 34714125 N DUP 5
A00297:158:HT275DSXX:1:1428:21350:28479 chr16 34714054 N chr16 34714125 N DUP 5
A00404:156:HV37TDSXX:2:1146:12771:23077 chr16 34714054 N chr16 34714125 N DUP 5
A00404:155:HV27LDSXX:1:2578:12011:23610 chr16 34714054 N chr16 34714125 N DUP 5
A00404:156:HV37TDSXX:2:2221:31412:10394 chr16 34714054 N chr16 34714125 N DUP 5
A00404:156:HV37TDSXX:2:1241:1389:22185 chr16 34714054 N chr16 34714125 N DUP 5
A00404:156:HV37TDSXX:3:2507:31720:35070 chr16 34714054 N chr16 34714125 N DUP 5
A00297:158:HT275DSXX:4:1435:26069:31203 chr16 34714054 N chr16 34714125 N DUP 5
A00297:158:HT275DSXX:4:1134:10221:26240 chr16 34714054 N chr16 34714125 N DUP 8
A00404:156:HV37TDSXX:3:1541:25852:31297 chr16 34714054 N chr16 34714125 N DUP 8
A00404:156:HV37TDSXX:2:2350:27263:27132 chr16 34714054 N chr16 34714125 N DUP 10
A00404:156:HV37TDSXX:3:2126:31394:17284 chr16 34714054 N chr16 34714125 N DUP 10
A00297:158:HT275DSXX:2:1329:3947:6010 chr16 34714054 N chr16 34714125 N DUP 10
A00297:158:HT275DSXX:3:2661:26865:30796 chr16 11598988 N chr16 11599288 N DEL 5
A00404:155:HV27LDSXX:1:2125:7591:13103 chr16 11599013 N chr16 11599311 N DUP 3
A00404:155:HV27LDSXX:1:2125:7600:13119 chr16 11599013 N chr16 11599311 N DUP 3
A00404:156:HV37TDSXX:3:1521:24243:14732 chr16 11599068 N chr16 11599368 N DEL 21
A00404:156:HV37TDSXX:2:1416:10619:35697 chr16 11599034 N chr16 11599334 N DEL 20
A00297:158:HT275DSXX:2:2572:10809:34898 chr16 11599044 N chr16 11599344 N DEL 3
A00404:156:HV37TDSXX:2:1416:9905:36871 chr16 11599161 N chr16 11599460 N DEL 5
A00404:156:HV37TDSXX:4:2404:18810:17347 chr7 158456242 N chr7 158456577 N DUP 5
A00297:158:HT275DSXX:2:1114:24117:11412 chr7 158456158 N chr7 158456289 N DUP 5
A00297:158:HT275DSXX:1:2307:10330:22357 chr7 158456158 N chr7 158456289 N DUP 5
A00297:158:HT275DSXX:1:1348:1588:18176 chr7 158456158 N chr7 158456289 N DUP 5
A00404:155:HV27LDSXX:1:2665:2130:6903 chr7 158456158 N chr7 158456289 N DUP 5
A00297:158:HT275DSXX:4:1352:29677:37012 chr7 158456364 N chr7 158456671 N DEL 10
A00297:158:HT275DSXX:2:1228:7636:23202 chr7 158456366 N chr7 158456571 N DEL 2
A00297:158:HT275DSXX:3:1442:28474:21778 chr7 158456304 N chr7 158456507 N DUP 5
A00297:158:HT275DSXX:4:1352:29677:37012 chr7 158456364 N chr7 158456671 N DEL 15
A00404:156:HV37TDSXX:1:2174:2392:1282 chr7 158456385 N chr7 158456692 N DEL 5
A00297:158:HT275DSXX:1:2126:11822:10817 chr7 158456417 N chr7 158456622 N DEL 15
A00404:155:HV27LDSXX:2:1221:13693:11021 chr7 158456484 N chr7 158456740 N DEL 2
A00297:158:HT275DSXX:1:2119:31015:25708 chr7 158456361 N chr7 158456564 N DUP 5
A00404:155:HV27LDSXX:3:1123:30987:9784 chr7 158456315 N chr7 158456469 N DEL 9
A00404:155:HV27LDSXX:1:2332:27941:20572 chr7 158456177 N chr7 158456514 N DEL 10
A00404:156:HV37TDSXX:3:1138:25292:20870 chr7 158456551 N chr7 158456601 N DUP 5
A00404:155:HV27LDSXX:3:1266:28330:18302 chr7 158456558 N chr7 158456661 N DEL 18
A00404:155:HV27LDSXX:1:1311:27335:32957 chr7 158456493 N chr7 158456545 N DEL 10
A00404:156:HV37TDSXX:4:1549:7889:20603 chr7 158456202 N chr7 158456692 N DEL 5
A00297:158:HT275DSXX:3:2128:30183:30530 chr7 158456653 N chr7 158456705 N DEL 2
A00404:156:HV37TDSXX:4:2453:6189:8954 chr9 133382624 N chr9 133383100 N DEL 3
A00404:156:HV37TDSXX:3:1257:17418:24017 chr9 133383009 N chr9 133383142 N DEL 5
A00297:158:HT275DSXX:3:2367:5330:5838 chr9 133383049 N chr9 133383180 N DUP 5
A00404:155:HV27LDSXX:1:2421:16631:13041 chr9 133383120 N chr9 133383430 N DUP 3
A00404:155:HV27LDSXX:2:2668:20057:9518 chr9 133383319 N chr9 133383432 N DUP 7
A00297:158:HT275DSXX:3:1419:8675:10160 chr9 133383407 N chr9 133383603 N DEL 10
A00404:155:HV27LDSXX:2:2361:29008:32315 chr9 133383443 N chr9 133383606 N DUP 28
A00404:156:HV37TDSXX:1:2416:19524:4899 chr9 133383443 N chr9 133383606 N DUP 25
A00404:156:HV37TDSXX:1:1533:28944:20494 chr9 133383443 N chr9 133383606 N DUP 17
A00404:156:HV37TDSXX:3:1419:23927:10770 chr9 133382708 N chr9 133383445 N DEL 10
A00404:156:HV37TDSXX:2:2547:5005:20556 chr9 133383451 N chr9 133383614 N DUP 7
A00404:156:HV37TDSXX:2:2310:12192:11992 chr9 133383445 N chr9 133383608 N DUP 13
A00404:156:HV37TDSXX:3:2463:8983:28604 chr9 133383453 N chr9 133383616 N DUP 5
A00404:155:HV27LDSXX:3:1123:21151:13855 chr9 133383587 N chr9 133383736 N DEL 5
A00404:155:HV27LDSXX:3:1123:22788:14622 chr9 133383587 N chr9 133383736 N DEL 5
A00297:158:HT275DSXX:1:2433:6180:29982 chr9 133383587 N chr9 133383736 N DEL 9
A00404:155:HV27LDSXX:2:1256:21531:35524 chr9 133383587 N chr9 133383736 N DEL 9
A00297:158:HT275DSXX:4:2210:1570:36808 chr9 133383587 N chr9 133383736 N DEL 10
A00297:158:HT275DSXX:2:2507:14940:26303 chr9 133383587 N chr9 133383736 N DEL 13
A00404:156:HV37TDSXX:3:2666:2627:21699 chr9 133383587 N chr9 133383736 N DEL 25
A00297:158:HT275DSXX:2:1277:25816:28948 chr9 133383587 N chr9 133383736 N DEL 33
A00297:158:HT275DSXX:2:2164:19877:13933 chr9 133383587 N chr9 133383736 N DEL 33
A00297:158:HT275DSXX:2:2164:19985:13714 chr9 133383587 N chr9 133383736 N DEL 33
A00404:156:HV37TDSXX:3:1209:17481:10817 chr9 133383587 N chr9 133383736 N DEL 37
A00297:158:HT275DSXX:1:2430:6894:36104 chr9 133382912 N chr9 133383685 N DUP 21
A00297:158:HT275DSXX:3:1524:4291:4820 chr9 133383198 N chr9 133383728 N DUP 6
A00404:156:HV37TDSXX:3:1574:12400:26412 chr9 133383198 N chr9 133383728 N DUP 7
A00404:155:HV27LDSXX:1:1676:26539:17049 chr9 133383537 N chr9 133383657 N DEL 32
A00297:158:HT275DSXX:1:2443:12454:9533 chr9 133383443 N chr9 133383754 N DUP 22
A00404:155:HV27LDSXX:2:1223:17381:30091 chr9 133382939 N chr9 133383660 N DEL 9
A00404:155:HV27LDSXX:4:1132:23701:33426 chr9 133382911 N chr9 133383662 N DEL 7
A00404:155:HV27LDSXX:2:1252:9634:23625 chr9 133382912 N chr9 133383663 N DEL 6
A00404:155:HV27LDSXX:1:1209:30707:30655 chr9 133382925 N chr9 133383780 N DUP 16
A00297:158:HT275DSXX:3:1253:2953:24706 chr9 133382896 N chr9 133383781 N DUP 22
A00404:155:HV27LDSXX:1:2242:14416:31939 chr9 133383443 N chr9 133383754 N DUP 30
A00297:158:HT275DSXX:3:2475:11605:32424 chr9 133383443 N chr9 133383754 N DUP 32
A00404:155:HV27LDSXX:4:1416:6686:4053 chr9 133383587 N chr9 133383736 N DEL 16
A00297:158:HT275DSXX:2:1147:17689:4758 chr9 133383587 N chr9 133383736 N DEL 10
A00404:155:HV27LDSXX:1:1535:3296:35196 chr9 133383587 N chr9 133383736 N DEL 5
A00404:156:HV37TDSXX:3:2530:6903:15515 chr9 133383587 N chr9 133383736 N DEL 5
A00297:158:HT275DSXX:1:2344:18295:27070 chr9 133383589 N chr9 133383738 N DEL 5
A00297:158:HT275DSXX:1:2344:18511:18458 chr9 133383589 N chr9 133383738 N DEL 5
A00404:155:HV27LDSXX:2:2527:20021:22482 chr9 133383590 N chr9 133383739 N DEL 5
A00404:156:HV37TDSXX:3:1128:26503:7247 chr9 133383590 N chr9 133383739 N DEL 5
A00297:158:HT275DSXX:1:2560:13792:6965 chr9 133383212 N chr9 133383744 N DEL 5
A00404:156:HV37TDSXX:2:2122:21359:32064 chr9 133383261 N chr9 133383746 N DEL 3
A00404:155:HV27LDSXX:1:1563:11288:6793 chr12 124333989 N chr12 124334124 N DEL 3
A00297:158:HT275DSXX:1:2345:17707:17253 chr12 124333989 N chr12 124334124 N DEL 4
A00297:158:HT275DSXX:4:1230:15980:7467 chr12 124334014 N chr12 124334117 N DEL 10
A00297:158:HT275DSXX:2:2236:13431:30358 chr12 124333990 N chr12 124334155 N DUP 31
A00404:156:HV37TDSXX:1:2145:1597:7169 chr12 124334033 N chr12 124334154 N DUP 32
A00297:158:HT275DSXX:3:1476:13792:13667 chr12 124334033 N chr12 124334154 N DUP 29
A00404:155:HV27LDSXX:1:2376:10963:16219 chr12 124334033 N chr12 124334154 N DUP 27
A00404:156:HV37TDSXX:4:1313:32244:19382 chr12 124334033 N chr12 124334154 N DUP 25
A00297:158:HT275DSXX:4:2208:12554:32033 chr12 124334033 N chr12 124334154 N DUP 25
A00297:158:HT275DSXX:3:2418:13566:3662 chr12 124333990 N chr12 124334155 N DUP 13
A00404:155:HV27LDSXX:3:1159:24270:12430 chr12 124334019 N chr12 124334154 N DUP 2
A00297:158:HT275DSXX:3:1416:25003:2487 chr12 124334006 N chr12 124334141 N DUP 3
A00404:155:HV27LDSXX:4:1446:15329:30953 chr12 124334036 N chr12 124334125 N DUP 14
A00404:156:HV37TDSXX:3:2502:31340:35352 chr12 124334049 N chr12 124334170 N DUP 8
A00297:158:HT275DSXX:1:2112:8693:17863 chr12 124333989 N chr12 124334124 N DEL 10
A00404:155:HV27LDSXX:3:1234:19795:4366 chr5 135754153 N chr5 135754292 N DEL 5
A00297:158:HT275DSXX:3:1474:19072:19492 chr8 94591333 N chr8 94591511 N DEL 5
A00404:155:HV27LDSXX:3:2604:18141:19758 chr8 94591314 N chr8 94591391 N DUP 5
A00297:158:HT275DSXX:3:1157:17888:5008 chr8 94591334 N chr8 94591510 N DUP 5
A00297:158:HT275DSXX:2:2462:25491:9126 chr8 94591461 N chr8 94591762 N DUP 4
A00404:155:HV27LDSXX:1:1115:22200:10379 chr8 94591279 N chr8 94591455 N DUP 5
A00404:155:HV27LDSXX:1:2342:2799:27978 chr8 94591426 N chr8 94591477 N DEL 1
A00297:158:HT275DSXX:3:1474:19072:19492 chr8 94591608 N chr8 94591785 N DEL 5
A00404:155:HV27LDSXX:3:1355:4083:28917 chr8 94591608 N chr8 94591785 N DEL 5
A00297:158:HT275DSXX:4:1566:3857:34100 chr8 94591608 N chr8 94591785 N DEL 5
A00404:156:HV37TDSXX:1:2641:6479:21887 chr8 94591408 N chr8 94591586 N DEL 5
A00404:155:HV27LDSXX:4:1332:8721:13307 chr8 94591288 N chr8 94591669 N DUP 1
A00297:158:HT275DSXX:1:1374:29423:15280 chr8 94591366 N chr8 94591718 N DUP 14
A00297:158:HT275DSXX:3:1409:16360:11976 chr8 94591428 N chr8 94591731 N DEL 14
A00404:155:HV27LDSXX:2:1618:12373:23296 chr8 94591428 N chr8 94591731 N DEL 14
A00404:156:HV37TDSXX:4:1558:17517:27414 chr8 94591428 N chr8 94591731 N DEL 14
A00404:155:HV27LDSXX:4:1232:6171:13401 chr8 94591455 N chr8 94591758 N DEL 8
A00404:155:HV27LDSXX:2:1375:17011:28479 chr8 94591756 N chr8 94591886 N DUP 10
A00404:155:HV27LDSXX:1:2117:29487:3176 chr5 57518786 N chr5 57518903 N DEL 26
A00404:156:HV37TDSXX:1:1675:17327:5415 chr3 127155936 N chr3 127156005 N DEL 4
A00297:158:HT275DSXX:4:2672:9995:25880 chr3 127155917 N chr3 127156182 N DUP 5
A00297:158:HT275DSXX:3:1167:31575:30592 chr3 127155917 N chr3 127156182 N DUP 5
A00404:156:HV37TDSXX:3:1364:17815:10081 chr3 127155917 N chr3 127156182 N DUP 5
A00404:156:HV37TDSXX:4:2445:7591:34178 chr3 127155940 N chr3 127156177 N DEL 5
A00404:155:HV27LDSXX:1:2656:26006:22983 chr21 44504203 N chr21 44504373 N DEL 5
A00404:156:HV37TDSXX:1:2222:27019:27712 chr21 44504114 N chr21 44504377 N DEL 14
A00404:155:HV27LDSXX:4:2421:14452:27085 chr1 75906598 N chr1 75906660 N DUP 19
A00297:158:HT275DSXX:2:1121:32922:32049 chr1 75906598 N chr1 75906660 N DUP 26
A00297:158:HT275DSXX:2:1220:2437:7467 chr1 75906598 N chr1 75906660 N DUP 26
A00297:158:HT275DSXX:2:1618:31024:36558 chr1 75906594 N chr1 75906692 N DUP 11
A00297:158:HT275DSXX:2:1619:29686:22874 chr1 75906594 N chr1 75906692 N DUP 11
A00404:155:HV27LDSXX:4:1361:19587:34100 chr1 75906621 N chr1 75906715 N DUP 5
A00297:158:HT275DSXX:4:2328:12762:9690 chr22 47069799 N chr22 47069942 N DEL 4
A00404:155:HV27LDSXX:3:2350:27670:20948 chr22 47069799 N chr22 47069942 N DEL 7
A00297:158:HT275DSXX:4:2601:15555:31344 chr22 47069799 N chr22 47069942 N DEL 11
A00297:158:HT275DSXX:3:1401:32841:29027 chr22 47069799 N chr22 47069942 N DEL 17
A00297:158:HT275DSXX:2:2237:25220:13197 chr22 47069799 N chr22 47069942 N DEL 17
A00404:156:HV37TDSXX:1:1432:14498:17331 chr22 47069799 N chr22 47069942 N DEL 17
A00404:155:HV27LDSXX:4:1346:18900:17534 chr22 47069799 N chr22 47069942 N DEL 17
A00404:156:HV37TDSXX:2:2243:13404:31125 chr22 47069875 N chr22 47070163 N DEL 5
A00297:158:HT275DSXX:4:1165:30228:32957 chr22 47069711 N chr22 47069875 N DUP 6
A00404:156:HV37TDSXX:2:1627:25590:9330 chr22 47069711 N chr22 47069875 N DUP 9
A00297:158:HT275DSXX:2:2127:6967:3662 chr22 47069856 N chr22 47069951 N DEL 18
A00404:156:HV37TDSXX:1:2268:25608:17691 chr22 47069962 N chr22 47070057 N DUP 24
A00404:156:HV37TDSXX:2:2611:20808:5932 chr22 47069856 N chr22 47069951 N DEL 22
A00297:158:HT275DSXX:2:1335:14651:19038 chr22 47069856 N chr22 47069951 N DEL 22
A00404:156:HV37TDSXX:2:1442:7419:13338 chr22 47069820 N chr22 47070057 N DUP 18
A00404:156:HV37TDSXX:2:1303:1832:25394 chr22 47069820 N chr22 47070057 N DUP 21
A00297:158:HT275DSXX:1:2475:4218:22952 chr22 47069749 N chr22 47069962 N DEL 9
A00297:158:HT275DSXX:1:2475:5385:24283 chr22 47069749 N chr22 47069962 N DEL 9
A00404:155:HV27LDSXX:2:2104:15501:21480 chr22 47069749 N chr22 47069962 N DEL 9
A00404:156:HV37TDSXX:2:2346:11017:22921 chr22 47069820 N chr22 47070057 N DUP 21
A00404:155:HV27LDSXX:2:1115:19352:18724 chr22 47069866 N chr22 47070010 N DEL 11
A00404:156:HV37TDSXX:4:1473:3586:17628 chr22 47069763 N chr22 47069976 N DEL 1
A00404:155:HV27LDSXX:1:1668:13648:28541 chr22 47069866 N chr22 47070010 N DEL 11
A00297:158:HT275DSXX:4:2429:26431:36151 chr22 47069866 N chr22 47070010 N DEL 11
A00404:156:HV37TDSXX:3:2248:30481:5744 chr22 47069866 N chr22 47070010 N DEL 11
A00297:158:HT275DSXX:3:2406:3703:21465 chr22 47069866 N chr22 47070010 N DEL 11
A00297:158:HT275DSXX:2:1417:15167:35336 chr22 47069866 N chr22 47070010 N DEL 11
A00404:156:HV37TDSXX:3:1267:5593:30780 chr22 47069866 N chr22 47070010 N DEL 11
A00404:155:HV27LDSXX:1:1274:2654:34460 chr22 47069866 N chr22 47070010 N DEL 11
A00404:155:HV27LDSXX:1:2174:31295:28416 chr22 47069866 N chr22 47070010 N DEL 11
A00404:156:HV37TDSXX:4:2233:6289:21621 chr22 47069866 N chr22 47070010 N DEL 11
A00404:155:HV27LDSXX:3:1333:11162:5666 chr22 47069866 N chr22 47070010 N DEL 11
A00404:156:HV37TDSXX:1:1113:18918:20322 chr22 47069866 N chr22 47070010 N DEL 11
A00297:158:HT275DSXX:4:2548:7491:14967 chr22 47069870 N chr22 47070014 N DEL 11
A00297:158:HT275DSXX:2:1645:2636:35524 chr22 47069876 N chr22 47070020 N DEL 5
A00404:156:HV37TDSXX:2:1555:17219:28588 chr1 125082639 N chr1 125082854 N DUP 5
A00404:156:HV37TDSXX:1:2217:26205:1783 chr1 125082639 N chr1 125082854 N DUP 5
A00297:158:HT275DSXX:2:2271:12210:10864 chr1 125082745 N chr1 125082816 N DUP 1
A00297:158:HT275DSXX:4:2219:15402:14262 chr1 125082696 N chr1 125082914 N DUP 2
A00404:156:HV37TDSXX:1:1205:19099:15562 chr1 125082844 N chr1 125082918 N DUP 1
A00404:156:HV37TDSXX:3:2253:24135:21746 chr1 125082893 N chr1 125082964 N DUP 5
A00404:155:HV27LDSXX:3:1630:17662:7310 chr5 56835433 N chr5 56835500 N DEL 3
A00404:155:HV27LDSXX:2:2556:28031:4914 chr5 56835433 N chr5 56835500 N DEL 7
A00404:155:HV27LDSXX:2:1470:28284:3004 chr5 56835445 N chr5 56835512 N DEL 3
A00404:155:HV27LDSXX:3:1348:24813:29309 chr5 56835437 N chr5 56835504 N DEL 11
A00404:156:HV37TDSXX:2:2622:23267:12164 chr5 56835437 N chr5 56835504 N DEL 11
A00297:158:HT275DSXX:3:2528:23764:2253 chr5 56835445 N chr5 56835512 N DEL 3
A00297:158:HT275DSXX:2:1315:17327:35790 chr5 56835442 N chr5 56835509 N DEL 5
A00404:155:HV27LDSXX:3:2352:17436:16031 chr21 7915792 N chr21 7915902 N DEL 5
A00297:158:HT275DSXX:3:2543:13657:2440 chr21 7915791 N chr21 7915959 N DEL 5
A00404:156:HV37TDSXX:4:2275:13160:35869 chr21 7915791 N chr21 7915975 N DEL 5
A00404:155:HV27LDSXX:4:1530:1407:32925 chr21 7915803 N chr21 7916036 N DEL 5
A00404:156:HV37TDSXX:1:1578:5846:2973 chr1 32720524 N chr1 32720599 N DEL 5
A00404:156:HV37TDSXX:2:2501:6985:24017 chr5 149729701 N chr5 149729820 N DEL 1
A00404:156:HV37TDSXX:2:2226:25201:30076 chr5 149729700 N chr5 149729821 N DEL 5
A00404:155:HV27LDSXX:3:2524:7581:10300 chr12 131635072 N chr12 131635263 N DUP 5
A00404:156:HV37TDSXX:2:1211:1561:18192 chr2 11380617 N chr2 11380696 N DUP 24
A00404:156:HV37TDSXX:4:1114:15049:9424 chr2 11380617 N chr2 11380696 N DUP 24
A00404:155:HV27LDSXX:2:1441:13720:28040 chr2 11380617 N chr2 11380714 N DUP 18
A00404:156:HV37TDSXX:2:1211:1090:20259 chr2 11380617 N chr2 11380696 N DUP 24
A00297:158:HT275DSXX:2:2628:30978:14716 chr2 11380596 N chr2 11380739 N DUP 14
A00404:156:HV37TDSXX:1:1247:8214:29465 chr1 125181621 N chr1 125181694 N DEL 3
A00404:156:HV37TDSXX:4:2444:23439:6292 chr1 125181621 N chr1 125181694 N DEL 5
A00404:155:HV27LDSXX:2:2117:13467:10786 chr1 125181621 N chr1 125181694 N DEL 5
A00297:158:HT275DSXX:1:1533:28221:33802 chr1 125181621 N chr1 125181694 N DEL 3
A00404:155:HV27LDSXX:3:1339:26078:2879 chr1 125181534 N chr1 125181627 N DUP 6
A00404:155:HV27LDSXX:1:2109:4390:3834 chr1 125181621 N chr1 125181694 N DEL 5
A00297:158:HT275DSXX:1:2363:25518:12305 chr1 125181621 N chr1 125181694 N DEL 2
A00404:156:HV37TDSXX:2:2370:17083:33332 chr1 125181621 N chr1 125181694 N DEL 5
A00404:156:HV37TDSXX:1:1533:8757:12493 chr1 125181549 N chr1 125181619 N DUP 8
A00404:156:HV37TDSXX:4:1404:11776:10019 chr1 125181621 N chr1 125181694 N DEL 2
A00404:156:HV37TDSXX:2:2470:1624:20462 chr1 125181473 N chr1 125181573 N DUP 8
A00404:155:HV27LDSXX:2:2128:3034:25942 chr1 125181621 N chr1 125181694 N DEL 5
A00404:155:HV27LDSXX:2:2668:11288:26177 chr1 125181383 N chr1 125181626 N DUP 3
A00404:156:HV37TDSXX:1:2429:18087:7858 chr1 125181621 N chr1 125181694 N DEL 5
A00297:158:HT275DSXX:2:1524:15899:12273 chr1 125181621 N chr1 125181694 N DEL 3
A00404:156:HV37TDSXX:2:2674:17083:25097 chr1 125181621 N chr1 125181694 N DEL 4
A00404:156:HV37TDSXX:3:2678:6325:27508 chr1 125181528 N chr1 125181693 N DUP 5
A00404:156:HV37TDSXX:1:1236:12002:25911 chr1 125181621 N chr1 125181694 N DEL 5
A00404:156:HV37TDSXX:3:2278:14678:9627 chr1 125181549 N chr1 125181619 N DUP 10
A00404:155:HV27LDSXX:3:2236:10574:18991 chr1 125181473 N chr1 125181573 N DUP 9
A00404:155:HV27LDSXX:3:2558:2230:18286 chr1 125181621 N chr1 125181694 N DEL 5
A00297:158:HT275DSXX:3:2523:2031:14716 chr1 125181530 N chr1 125181623 N DUP 5
A00404:156:HV37TDSXX:3:2240:22525:30577 chr1 125181621 N chr1 125181694 N DEL 5
A00297:158:HT275DSXX:2:1617:27489:1251 chr1 125181621 N chr1 125181694 N DEL 5
A00404:155:HV27LDSXX:4:1407:6189:4664 chr1 125181621 N chr1 125181694 N DEL 5
A00404:155:HV27LDSXX:2:1432:6180:13698 chr1 125181621 N chr1 125181694 N DEL 3
A00297:158:HT275DSXX:1:1426:13964:22075 chr1 125181621 N chr1 125181694 N DEL 5
A00404:156:HV37TDSXX:1:2136:13395:25379 chr1 125181449 N chr1 125181574 N DEL 5
A00297:158:HT275DSXX:1:1247:3459:23516 chr1 125181452 N chr1 125181577 N DEL 5
A00297:158:HT275DSXX:3:1112:10366:32158 chr8 37785292 N chr8 37785594 N DEL 1
A00297:158:HT275DSXX:3:1122:14362:5384 chr1 37579633 N chr1 37579983 N DEL 22
A00404:155:HV27LDSXX:2:1108:18349:5274 chr7 58036480 N chr7 58036580 N DUP 8
A00404:155:HV27LDSXX:2:2108:17888:13557 chr7 58036480 N chr7 58036580 N DUP 8
A00404:155:HV27LDSXX:2:2328:13241:5008 chr7 58036456 N chr7 58036605 N DUP 8
A00404:155:HV27LDSXX:3:1537:16541:33865 chr7 58036454 N chr7 58036580 N DUP 38
A00297:158:HT275DSXX:3:2644:13060:14278 chr3 195710380 N chr3 195710516 N DEL 5
A00404:156:HV37TDSXX:4:1430:15103:18818 chr3 195710430 N chr3 195710926 N DEL 5
A00404:156:HV37TDSXX:4:2469:30653:7138 chr3 195710457 N chr3 195711133 N DEL 10
A00297:158:HT275DSXX:4:1646:25717:31532 chr3 195710447 N chr3 195710673 N DEL 10
A00404:156:HV37TDSXX:4:1411:27416:15687 chr3 195710447 N chr3 195710673 N DEL 15
A00404:156:HV37TDSXX:4:2423:3577:28385 chr3 195710507 N chr3 195711529 N DEL 1
A00404:155:HV27LDSXX:4:1562:8079:32080 chr3 195710447 N chr3 195710673 N DEL 3
A00404:155:HV27LDSXX:1:1614:11053:26240 chr3 195710549 N chr3 195711571 N DEL 5
A00404:155:HV27LDSXX:1:2573:10854:19570 chr3 195710549 N chr3 195711571 N DEL 5
A00404:155:HV27LDSXX:1:1357:4291:32816 chr3 195710549 N chr3 195711571 N DEL 5
A00404:156:HV37TDSXX:2:1644:7428:31673 chr3 195710549 N chr3 195711571 N DEL 5
A00404:156:HV37TDSXX:1:2139:18430:9079 chr3 195710507 N chr3 195711529 N DEL 5
A00404:156:HV37TDSXX:3:1214:6126:33927 chr3 195710465 N chr3 195710599 N DUP 3
A00404:156:HV37TDSXX:2:1440:6515:20478 chr3 195710562 N chr3 195711148 N DEL 14
A00404:155:HV27LDSXX:1:2512:9950:33943 chr3 195710599 N chr3 195711095 N DEL 15
A00404:155:HV27LDSXX:3:2669:11948:10285 chr3 195710618 N chr3 195710979 N DEL 5
A00297:158:HT275DSXX:2:2233:13141:3145 chr3 195710644 N chr3 195711005 N DEL 4
A00404:155:HV27LDSXX:4:1342:30192:19930 chr3 195710618 N chr3 195710979 N DEL 5
A00297:158:HT275DSXX:4:1633:3893:23171 chr3 195710644 N chr3 195711005 N DEL 5
A00297:158:HT275DSXX:4:1565:31521:36886 chr3 195710428 N chr3 195710652 N DUP 5
A00297:158:HT275DSXX:3:2478:1072:8265 chr3 195710428 N chr3 195710652 N DUP 5
A00404:156:HV37TDSXX:2:2127:1624:36683 chr3 195710428 N chr3 195710652 N DUP 5
A00297:158:HT275DSXX:4:2273:10655:24831 chr3 195710428 N chr3 195710652 N DUP 5
A00404:156:HV37TDSXX:3:2536:4255:20040 chr3 195710428 N chr3 195710652 N DUP 5
A00297:158:HT275DSXX:1:2477:11397:16063 chr3 195710655 N chr3 195710926 N DEL 5
A00404:155:HV27LDSXX:4:1221:1316:36057 chr3 195710637 N chr3 195711043 N DEL 10
A00404:155:HV27LDSXX:3:2371:26639:30937 chr3 195710454 N chr3 195710590 N DEL 5
A00404:155:HV27LDSXX:1:1327:14452:4789 chr3 195710455 N chr3 195710591 N DEL 5
A00297:158:HT275DSXX:3:1532:18087:12900 chr3 195710542 N chr3 195710633 N DEL 15
A00404:155:HV27LDSXX:3:2107:6072:1611 chr3 195710687 N chr3 195710913 N DEL 5
A00404:155:HV27LDSXX:4:2424:9516:16250 chr3 195710700 N chr3 195710836 N DEL 15
A00404:155:HV27LDSXX:4:2424:9805:16157 chr3 195710700 N chr3 195710836 N DEL 15
A00297:158:HT275DSXX:2:1603:19434:8688 chr3 195710528 N chr3 195710619 N DEL 5
A00297:158:HT275DSXX:1:1464:17011:36025 chr3 195710700 N chr3 195710836 N DEL 15
A00404:155:HV27LDSXX:4:1221:1208:35336 chr3 195710687 N chr3 195710913 N DEL 5
A00404:155:HV27LDSXX:2:1308:3179:7435 chr3 195710655 N chr3 195710926 N DEL 20
A00297:158:HT275DSXX:3:2128:25816:11068 chr3 195710722 N chr3 195711308 N DEL 20
A00404:155:HV27LDSXX:2:2254:32027:22169 chr3 195710644 N chr3 195711095 N DEL 8
A00297:158:HT275DSXX:4:2369:13015:3928 chr3 195710700 N chr3 195710836 N DEL 20
A00404:155:HV27LDSXX:3:1537:6289:21778 chr3 195710700 N chr3 195711286 N DEL 21
A00297:158:HT275DSXX:4:2359:17155:14763 chr3 195710431 N chr3 195710700 N DUP 3
A00404:156:HV37TDSXX:2:1434:27299:32518 chr3 195710700 N chr3 195711286 N DEL 22
A00404:156:HV37TDSXX:1:1260:3622:34788 chr3 195710673 N chr3 195711032 N DUP 5
A00404:156:HV37TDSXX:3:1472:32741:27007 chr3 195710663 N chr3 195710889 N DEL 4
A00404:156:HV37TDSXX:4:2104:24270:28995 chr3 195710673 N chr3 195711032 N DUP 5
A00404:155:HV27LDSXX:2:2164:10366:31031 chr3 195710480 N chr3 195710706 N DEL 3
A00404:155:HV27LDSXX:1:1209:1759:36573 chr3 195710767 N chr3 195711083 N DEL 10
A00404:155:HV27LDSXX:4:2113:9833:5807 chr3 195710428 N chr3 195711012 N DUP 1
A00404:155:HV27LDSXX:1:2573:10854:19570 chr3 195710475 N chr3 195711151 N DEL 4
A00404:155:HV27LDSXX:4:2220:8513:34554 chr3 195710745 N chr3 195711286 N DEL 10
A00297:158:HT275DSXX:2:2620:12707:21120 chr3 195710590 N chr3 195711219 N DUP 30
A00404:155:HV27LDSXX:3:2501:9082:8359 chr3 195710777 N chr3 195711093 N DEL 10
A00404:156:HV37TDSXX:3:1472:32741:27007 chr3 195710931 N chr3 195711112 N DEL 7
A00404:155:HV27LDSXX:4:1571:27317:31454 chr3 195711087 N chr3 195711268 N DEL 5
A00297:158:HT275DSXX:2:1609:14516:18897 chr3 195710833 N chr3 195711192 N DUP 16
A00404:156:HV37TDSXX:1:1326:21242:35211 chr3 195710682 N chr3 195711401 N DUP 12
A00404:155:HV27LDSXX:4:2113:14371:2143 chr3 195710666 N chr3 195710802 N DEL 2
A00404:155:HV27LDSXX:4:1571:27317:31454 chr3 195710666 N chr3 195710802 N DEL 2
A00404:156:HV37TDSXX:3:2530:3007:26209 chr3 195710742 N chr3 195710833 N DEL 15
A00297:158:HT275DSXX:4:1116:32280:19288 chr3 195710653 N chr3 195710877 N DUP 5
A00404:155:HV27LDSXX:4:1108:31467:8171 chr3 195710745 N chr3 195710836 N DEL 17
A00297:158:HT275DSXX:4:1545:11089:20666 chr3 195710745 N chr3 195710836 N DEL 15
A00404:155:HV27LDSXX:3:2533:18982:31172 chr3 195710907 N chr3 195710996 N DUP 14
A00404:156:HV37TDSXX:1:1645:21296:18803 chr3 195710836 N chr3 195710925 N DUP 22
A00404:155:HV27LDSXX:4:1537:7798:19664 chr3 195710475 N chr3 195711196 N DEL 8
A00297:158:HT275DSXX:3:2638:18457:5306 chr3 195711058 N chr3 195711372 N DUP 10
A00404:156:HV37TDSXX:1:1648:28962:16517 chr3 195710643 N chr3 195711002 N DUP 14
A00404:156:HV37TDSXX:2:2268:31467:2378 chr3 195710878 N chr3 195711012 N DUP 13
A00404:155:HV27LDSXX:1:1646:7500:28510 chr3 195710873 N chr3 195711142 N DUP 10
A00404:156:HV37TDSXX:4:2108:32154:19977 chr3 195710732 N chr3 195710868 N DEL 10
A00404:155:HV27LDSXX:4:1310:2266:30749 chr3 195710633 N chr3 195711217 N DUP 15
A00404:155:HV27LDSXX:4:1342:30192:19930 chr3 195710788 N chr3 195710879 N DEL 15
A00297:158:HT275DSXX:2:1169:12328:1799 chr3 195710547 N chr3 195710863 N DEL 10
A00404:156:HV37TDSXX:2:2330:4074:2096 chr3 195710547 N chr3 195710863 N DEL 10
A00404:155:HV27LDSXX:4:1564:12165:30389 chr3 195710878 N chr3 195711372 N DUP 10
A00297:158:HT275DSXX:1:2452:3694:5447 chr3 195710542 N chr3 195710633 N DEL 16
A00404:155:HV27LDSXX:1:2625:5321:2785 chr3 195710683 N chr3 195711357 N DUP 6
A00404:155:HV27LDSXX:1:2609:11342:22420 chr3 195710537 N chr3 195710898 N DEL 14
A00404:156:HV37TDSXX:1:1245:11017:14340 chr3 195710925 N chr3 195711151 N DEL 14
A00404:156:HV37TDSXX:2:1424:9435:26757 chr3 195710661 N chr3 195711200 N DUP 16
A00404:155:HV27LDSXX:4:1564:12165:30389 chr3 195710876 N chr3 195711010 N DUP 2
A00404:155:HV27LDSXX:2:2652:29577:33739 chr3 195710537 N chr3 195710898 N DEL 8
A00404:155:HV27LDSXX:4:1516:25654:32550 chr3 195710882 N chr3 195711016 N DUP 5
A00404:155:HV27LDSXX:1:2609:11342:22420 chr3 195710658 N chr3 195710884 N DEL 5
A00404:155:HV27LDSXX:4:2238:4010:11819 chr3 195711182 N chr3 195711273 N DEL 10
A00404:156:HV37TDSXX:1:1245:11017:14340 chr3 195710541 N chr3 195710902 N DEL 5
A00404:156:HV37TDSXX:1:1277:13774:5995 chr3 195710664 N chr3 195710890 N DEL 3
A00404:155:HV27LDSXX:3:1477:1334:4147 chr3 195711103 N chr3 195711372 N DUP 15
A00297:158:HT275DSXX:1:2101:25500:5008 chr3 195710667 N chr3 195710801 N DUP 2
A00297:158:HT275DSXX:2:1360:14190:29888 chr3 195710700 N chr3 195711286 N DEL 16
A00404:155:HV27LDSXX:2:1409:28483:3286 chr3 195710700 N chr3 195711286 N DEL 16
A00297:158:HT275DSXX:2:2646:16369:28401 chr3 195710700 N chr3 195711286 N DEL 15
A00404:155:HV27LDSXX:2:1564:11758:35164 chr3 195710700 N chr3 195711286 N DEL 15
A00404:155:HV27LDSXX:2:1564:12906:34992 chr3 195710700 N chr3 195711286 N DEL 15
A00297:158:HT275DSXX:2:2444:25581:4679 chr3 195710449 N chr3 195710900 N DEL 5
A00404:156:HV37TDSXX:2:2344:13476:2127 chr3 195710656 N chr3 195710925 N DUP 20
A00404:155:HV27LDSXX:3:2412:1380:7169 chr3 195710428 N chr3 195711012 N DUP 1
A00404:156:HV37TDSXX:1:1469:1570:36871 chr3 195710643 N chr3 195711002 N DUP 6
A00404:155:HV27LDSXX:1:2539:13566:33630 chr3 195710970 N chr3 195711331 N DEL 5
A00404:155:HV27LDSXX:3:2260:29613:26381 chr3 195710428 N chr3 195711012 N DUP 5
A00297:158:HT275DSXX:2:1609:14516:18897 chr3 195711012 N chr3 195711148 N DEL 8
A00404:155:HV27LDSXX:1:2539:13566:33630 chr3 195710878 N chr3 195711012 N DUP 21
A00404:155:HV27LDSXX:2:2351:9435:15358 chr3 195711012 N chr3 195711148 N DEL 15
A00404:155:HV27LDSXX:4:2134:14769:29481 chr3 195710789 N chr3 195711013 N DUP 10
A00297:158:HT275DSXX:2:2618:13783:10614 chr3 195710789 N chr3 195711013 N DUP 15
A00404:155:HV27LDSXX:4:1511:17192:1204 chr3 195710789 N chr3 195711013 N DUP 15
A00297:158:HT275DSXX:1:1569:8061:9095 chr3 195711148 N chr3 195711372 N DUP 10
A00297:158:HT275DSXX:3:2372:4083:18458 chr3 195710542 N chr3 195710633 N DEL 16
A00404:155:HV27LDSXX:3:1220:21838:13855 chr3 195710516 N chr3 195711057 N DEL 3
A00404:156:HV37TDSXX:1:1307:30915:31172 chr3 195710475 N chr3 195711061 N DEL 7
A00297:158:HT275DSXX:1:2276:28293:8813 chr3 195711108 N chr3 195711377 N DUP 10
A00404:155:HV27LDSXX:4:2206:1334:36025 chr3 195710701 N chr3 195711375 N DUP 13
A00404:156:HV37TDSXX:4:1232:31467:26584 chr3 195710732 N chr3 195711093 N DEL 11
A00404:155:HV27LDSXX:1:2515:30770:8187 chr3 195711033 N chr3 195711347 N DUP 5
A00404:156:HV37TDSXX:1:1307:30915:31172 chr3 195711124 N chr3 195711348 N DUP 10
A00404:155:HV27LDSXX:2:1251:14516:25473 chr3 195711148 N chr3 195711372 N DUP 7
A00404:156:HV37TDSXX:4:1433:32226:19163 chr3 195710798 N chr3 195711069 N DEL 5
A00404:156:HV37TDSXX:1:2174:12093:7310 chr3 195710745 N chr3 195710836 N DEL 25
A00404:155:HV27LDSXX:1:1208:31259:11631 chr3 195710665 N chr3 195711071 N DEL 2
A00404:155:HV27LDSXX:1:2208:32018:16141 chr3 195710665 N chr3 195711071 N DEL 2
A00404:155:HV27LDSXX:3:2340:17508:25895 chr3 195711103 N chr3 195711372 N DUP 15
A00404:156:HV37TDSXX:4:1232:31467:26584 chr3 195710711 N chr3 195711072 N DEL 4
A00404:155:HV27LDSXX:2:2509:5023:35650 chr3 195711103 N chr3 195711372 N DUP 15
A00404:155:HV27LDSXX:1:1451:32127:23563 chr3 195710898 N chr3 195711124 N DEL 10
A00404:156:HV37TDSXX:1:2635:27480:17738 chr3 195710672 N chr3 195711078 N DEL 5
A00404:155:HV27LDSXX:1:1305:19940:33583 chr3 195710732 N chr3 195711093 N DEL 5
A00404:156:HV37TDSXX:3:2217:6686:25880 chr3 195710672 N chr3 195711033 N DEL 5
A00404:155:HV27LDSXX:4:2430:27534:28322 chr3 195710913 N chr3 195711362 N DUP 7
A00404:155:HV27LDSXX:2:2535:6180:8500 chr3 195711147 N chr3 195711371 N DUP 5
A00404:156:HV37TDSXX:2:1168:11550:34679 chr3 195710547 N chr3 195711088 N DEL 5
A00404:155:HV27LDSXX:1:1121:28384:32612 chr3 195711148 N chr3 195711372 N DUP 10
A00404:156:HV37TDSXX:1:1102:22968:36511 chr3 195710502 N chr3 195711401 N DUP 15
A00404:155:HV27LDSXX:3:1404:15953:26960 chr3 195710574 N chr3 195710888 N DUP 20
A00297:158:HT275DSXX:4:2108:13819:15092 chr3 195711088 N chr3 195711357 N DUP 10
A00404:155:HV27LDSXX:4:2430:27534:28322 chr3 195711123 N chr3 195711347 N DUP 5
A00404:155:HV27LDSXX:3:2617:9878:21574 chr3 195710507 N chr3 195711093 N DEL 5
A00404:156:HV37TDSXX:1:1245:10773:13416 chr3 195711091 N chr3 195711360 N DUP 7
A00297:158:HT275DSXX:2:2620:12707:21120 chr3 195710427 N chr3 195711371 N DUP 10
A00404:155:HV27LDSXX:2:1302:23592:27132 chr3 195710643 N chr3 195710957 N DUP 16
A00404:156:HV37TDSXX:4:1430:15103:18818 chr3 195710428 N chr3 195711372 N DUP 8
A00297:158:HT275DSXX:2:2602:13829:13416 chr3 195710746 N chr3 195711330 N DUP 8
A00404:155:HV27LDSXX:2:2652:29577:33739 chr3 195710878 N chr3 195711012 N DUP 20
A00404:155:HV27LDSXX:4:1433:28537:13526 chr3 195710789 N chr3 195711148 N DUP 15
A00404:155:HV27LDSXX:1:1314:23348:12430 chr3 195710921 N chr3 195711147 N DEL 5
A00404:156:HV37TDSXX:3:1415:27697:3364 chr3 195710468 N chr3 195711189 N DEL 5
A00297:158:HT275DSXX:2:2618:13783:10614 chr3 195710897 N chr3 195711123 N DEL 5
A00404:156:HV37TDSXX:4:1617:23900:23469 chr3 195710746 N chr3 195711330 N DUP 12
A00404:156:HV37TDSXX:4:1617:23900:23657 chr3 195710746 N chr3 195711330 N DUP 12
A00404:155:HV27LDSXX:1:1208:31259:11631 chr3 195710654 N chr3 195711105 N DEL 8
A00404:156:HV37TDSXX:3:1349:21052:5134 chr3 195710798 N chr3 195711202 N DUP 11
A00297:158:HT275DSXX:2:1449:20383:20635 chr3 195710735 N chr3 195710871 N DEL 7
A00404:155:HV27LDSXX:4:1140:2528:36871 chr3 195710429 N chr3 195711193 N DUP 3
A00404:155:HV27LDSXX:2:1302:23592:27132 chr3 195710628 N chr3 195710897 N DUP 9
A00404:156:HV37TDSXX:1:2340:23511:28964 chr3 195711047 N chr3 195711361 N DUP 10
A00404:156:HV37TDSXX:4:2167:1533:26631 chr3 195710925 N chr3 195711061 N DEL 5
A00297:158:HT275DSXX:2:1169:12328:1799 chr3 195710722 N chr3 195711128 N DEL 5
A00404:156:HV37TDSXX:2:2344:13476:2127 chr3 195711148 N chr3 195711372 N DUP 10
A00297:158:HT275DSXX:3:1441:25129:33833 chr3 195710668 N chr3 195711074 N DEL 5
A00297:158:HT275DSXX:4:2273:10655:24831 chr3 195710482 N chr3 195711113 N DEL 5
A00297:158:HT275DSXX:1:2178:3441:10614 chr3 195710878 N chr3 195711012 N DUP 22
A00404:156:HV37TDSXX:4:2167:1533:26631 chr3 195710897 N chr3 195711123 N DEL 5
A00404:155:HV27LDSXX:2:2351:9435:15358 chr3 195711097 N chr3 195711186 N DUP 5
A00297:158:HT275DSXX:3:2676:21965:17769 chr3 195710633 N chr3 195711217 N DUP 15
A00404:155:HV27LDSXX:3:2302:8703:10363 chr3 195710672 N chr3 195711123 N DEL 5
A00404:155:HV27LDSXX:4:2174:6126:6872 chr3 195710475 N chr3 195711151 N DEL 10
A00297:158:HT275DSXX:3:2513:17698:25316 chr3 195710878 N chr3 195711012 N DUP 15
A00404:156:HV37TDSXX:2:2663:20681:32800 chr3 195710732 N chr3 195711138 N DEL 10
A00297:158:HT275DSXX:4:1474:8585:15577 chr3 195711223 N chr3 195711357 N DUP 7
A00404:155:HV27LDSXX:2:1416:2419:10629 chr3 195710507 N chr3 195711273 N DEL 7
A00404:156:HV37TDSXX:1:2215:26196:4460 chr3 195710781 N chr3 195711277 N DEL 7
A00297:158:HT275DSXX:2:2518:7527:35697 chr3 195710458 N chr3 195711044 N DEL 5
A00297:158:HT275DSXX:1:2361:18502:3693 chr3 195711058 N chr3 195711372 N DUP 10
A00297:158:HT275DSXX:1:2162:26187:19382 chr3 195711193 N chr3 195711284 N DEL 5
A00404:155:HV27LDSXX:1:1209:1759:36573 chr3 195710656 N chr3 195710745 N DUP 10
A00404:155:HV27LDSXX:2:1308:3179:7435 chr3 195711148 N chr3 195711372 N DUP 10
A00404:156:HV37TDSXX:4:1118:23538:3991 chr3 195710878 N chr3 195711012 N DUP 15
A00404:155:HV27LDSXX:4:1511:17192:1204 chr3 195711058 N chr3 195711372 N DUP 9
A00404:156:HV37TDSXX:2:1168:11550:34679 chr3 195710701 N chr3 195711195 N DUP 16
A00404:156:HV37TDSXX:4:1433:32226:19163 chr3 195711193 N chr3 195711284 N DEL 5
A00404:155:HV27LDSXX:3:1134:23475:34820 chr3 195710475 N chr3 195711151 N DEL 10
A00297:158:HT275DSXX:3:2303:29586:8641 chr3 195711187 N chr3 195711278 N DEL 5
A00297:158:HT275DSXX:4:2369:13015:3928 chr3 195710470 N chr3 195711191 N DEL 5
A00404:156:HV37TDSXX:2:2268:31467:2378 chr3 195710970 N chr3 195711061 N DEL 15
A00404:155:HV27LDSXX:3:2533:18982:31172 chr3 195710475 N chr3 195711151 N DEL 5
A00404:155:HV27LDSXX:2:1162:31575:35352 chr3 195710898 N chr3 195711032 N DUP 10
A00297:158:HT275DSXX:1:1635:29053:25661 chr3 195710513 N chr3 195711144 N DEL 4
A00404:156:HV37TDSXX:3:1349:21052:5134 chr3 195710427 N chr3 195710921 N DUP 15
A00297:158:HT275DSXX:4:2118:31367:12195 chr3 195710594 N chr3 195710773 N DUP 10
A00297:158:HT275DSXX:3:2465:31195:4445 chr3 195710808 N chr3 195711169 N DEL 5
A00404:155:HV27LDSXX:3:1477:1334:4147 chr3 195710628 N chr3 195710897 N DUP 15
A00297:158:HT275DSXX:1:1153:15049:2503 chr3 195710628 N chr3 195710897 N DUP 15
A00297:158:HT275DSXX:1:2670:18403:26569 chr3 195710725 N chr3 195711477 N DEL 21
A00404:155:HV27LDSXX:4:2325:27697:12352 chr3 195710711 N chr3 195711162 N DEL 4
A00297:158:HT275DSXX:1:1249:16947:36699 chr3 195710713 N chr3 195711164 N DEL 2
A00404:156:HV37TDSXX:1:2215:26196:4460 chr3 195710789 N chr3 195711238 N DUP 15
A00404:156:HV37TDSXX:2:2663:20690:32377 chr3 195710503 N chr3 195711267 N DUP 5
A00297:158:HT275DSXX:3:2468:17761:29183 chr3 195710647 N chr3 195710961 N DUP 20
A00297:158:HT275DSXX:4:1474:8585:15577 chr3 195710925 N chr3 195711061 N DEL 10
A00404:156:HV37TDSXX:4:1641:5538:28651 chr3 195710872 N chr3 195711186 N DUP 4
A00404:156:HV37TDSXX:4:2654:20274:23954 chr3 195710837 N chr3 195710926 N DUP 25
A00297:158:HT275DSXX:4:2108:13819:15092 chr3 195710777 N chr3 195710958 N DEL 10
A00404:155:HV27LDSXX:2:2550:9435:6997 chr3 195710837 N chr3 195711241 N DUP 10
A00404:155:HV27LDSXX:2:1251:14516:25473 chr3 195710426 N chr3 195711280 N DUP 5
A00404:155:HV27LDSXX:4:1140:2528:36871 chr3 195710547 N chr3 195710863 N DEL 15
A00297:158:HT275DSXX:4:1327:19262:30185 chr3 195710594 N chr3 195711223 N DUP 5
A00404:156:HV37TDSXX:4:1613:9091:15922 chr3 195710510 N chr3 195711096 N DEL 5
A00297:158:HT275DSXX:1:1442:3568:32002 chr3 195710475 N chr3 195710836 N DEL 10
A00404:156:HV37TDSXX:4:1538:19361:3396 chr3 195710516 N chr3 195711057 N DEL 3
A00404:156:HV37TDSXX:2:2138:12237:12571 chr3 195710823 N chr3 195711229 N DEL 12
A00404:155:HV27LDSXX:1:2208:32018:16141 chr3 195710654 N chr3 195711195 N DEL 5
A00404:155:HV27LDSXX:2:2371:20491:21010 chr3 195710661 N chr3 195711202 N DEL 5
A00404:156:HV37TDSXX:2:2374:14045:23156 chr3 195710837 N chr3 195711151 N DUP 5
A00404:155:HV27LDSXX:3:2464:7961:29340 chr3 195710547 N chr3 195711223 N DEL 5
A00297:158:HT275DSXX:4:2658:28646:22921 chr3 195710745 N chr3 195710836 N DEL 20
A00404:156:HV37TDSXX:2:1455:19587:5353 chr3 195711048 N chr3 195711362 N DUP 7
A00404:156:HV37TDSXX:3:1401:22019:10692 chr3 195710823 N chr3 195711362 N DUP 5
A00404:156:HV37TDSXX:4:2358:21034:17816 chr3 195710507 N chr3 195711273 N DEL 20
A00297:158:HT275DSXX:2:1174:18059:28823 chr3 195711258 N chr3 195711347 N DUP 5
A00297:158:HT275DSXX:4:2371:11062:11130 chr3 195711012 N chr3 195711283 N DEL 10
A00404:155:HV27LDSXX:4:2134:14769:29481 chr3 195711179 N chr3 195711270 N DEL 10
A00404:156:HV37TDSXX:1:2139:18430:9079 chr3 195710507 N chr3 195711228 N DEL 5
A00297:158:HT275DSXX:1:2162:26187:19382 chr3 195710657 N chr3 195711241 N DUP 5
A00297:158:HT275DSXX:4:2658:28646:22921 chr3 195710657 N chr3 195711331 N DUP 5
A00297:158:HT275DSXX:2:1561:1768:8249 chr3 195710511 N chr3 195711232 N DEL 5
A00404:155:HV27LDSXX:3:2371:26639:30937 chr3 195710788 N chr3 195710879 N DEL 10
A00404:156:HV37TDSXX:4:1370:27733:11882 chr3 195710657 N chr3 195711331 N DUP 5
A00404:156:HV37TDSXX:1:2565:12924:1767 chr3 195711011 N chr3 195711237 N DEL 1
A00404:155:HV27LDSXX:2:2362:17644:27821 chr3 195710830 N chr3 195710966 N DEL 7
A00404:156:HV37TDSXX:3:2504:26160:2895 chr3 195710878 N chr3 195711012 N DUP 23
A00404:155:HV27LDSXX:1:2642:20826:29042 chr3 195711089 N chr3 195711270 N DEL 5
A00404:156:HV37TDSXX:1:1245:10773:13416 chr3 195710537 N chr3 195710898 N DEL 5
A00404:155:HV27LDSXX:1:1646:7500:28510 chr3 195710898 N chr3 195711032 N DUP 10
A00297:158:HT275DSXX:3:1538:1832:5697 chr3 195711099 N chr3 195711280 N DEL 5
A00404:155:HV27LDSXX:3:1144:24008:1329 chr3 195710700 N chr3 195711286 N DEL 16
A00404:156:HV37TDSXX:4:2504:20537:3270 chr3 195710700 N chr3 195711286 N DEL 15
A00297:158:HT275DSXX:1:2347:18828:25770 chr3 195710777 N chr3 195710958 N DEL 10
A00404:155:HV27LDSXX:2:2254:32027:22169 chr3 195710700 N chr3 195711286 N DEL 15
A00297:158:HT275DSXX:4:1545:11089:20666 chr3 195710833 N chr3 195711192 N DUP 6
A00404:155:HV27LDSXX:4:2532:30590:5776 chr3 195710700 N chr3 195711286 N DEL 15
A00297:158:HT275DSXX:2:1174:18059:28823 chr3 195710788 N chr3 195711284 N DEL 5
A00404:155:HV27LDSXX:3:1420:1434:34350 chr3 195710700 N chr3 195711286 N DEL 15
A00404:155:HV27LDSXX:1:1320:29812:26788 chr3 195710788 N chr3 195711284 N DEL 5
A00404:155:HV27LDSXX:1:2321:28022:15421 chr3 195710788 N chr3 195711284 N DEL 5
A00297:158:HT275DSXX:1:1569:8061:9095 chr3 195710428 N chr3 195711372 N DUP 2
A00297:158:HT275DSXX:2:1144:24975:11146 chr3 195710878 N chr3 195711372 N DUP 15
A00297:158:HT275DSXX:3:1478:1307:31688 chr3 195710518 N chr3 195711284 N DEL 5
A00404:155:HV27LDSXX:3:2204:25807:15530 chr3 195710836 N chr3 195710925 N DUP 20
A00404:156:HV37TDSXX:3:1165:17933:19899 chr3 195710970 N chr3 195711331 N DEL 5
A00404:156:HV37TDSXX:4:1144:27887:25488 chr3 195711148 N chr3 195711372 N DUP 10
A00404:155:HV27LDSXX:1:1121:28384:32612 chr3 195710789 N chr3 195711373 N DUP 10
A00404:156:HV37TDSXX:2:2374:14045:23156 chr3 195710836 N chr3 195710925 N DUP 25
A00404:155:HV27LDSXX:3:2462:8712:7529 chr3 195710475 N chr3 195711331 N DEL 5
A00404:155:HV27LDSXX:4:2206:1334:36025 chr3 195710833 N chr3 195710922 N DUP 20
A00297:158:HT275DSXX:1:2310:18909:15389 chr3 195710789 N chr3 195711013 N DUP 15
A00404:155:HV27LDSXX:1:2131:28483:10113 chr3 195710475 N chr3 195711331 N DEL 5
A00297:158:HT275DSXX:1:2657:20564:23265 chr3 195710476 N chr3 195711332 N DEL 5
A00297:158:HT275DSXX:3:2314:15338:17534 chr3 195711452 N chr3 195711619 N DEL 7
A00404:155:HV27LDSXX:1:1458:30798:21480 chr3 195711407 N chr3 195711574 N DEL 16
A00297:158:HT275DSXX:1:2452:3694:5447 chr3 195711183 N chr3 195711409 N DEL 20
A00404:156:HV37TDSXX:2:1627:29387:32471 chr3 195710897 N chr3 195711393 N DEL 15
A00404:156:HV37TDSXX:2:2511:16206:30718 chr3 195710595 N chr3 195711406 N DEL 11
A00404:155:HV27LDSXX:3:1144:24008:1329 chr3 195710595 N chr3 195711406 N DEL 10
A00404:156:HV37TDSXX:4:1511:26521:36276 chr3 195710595 N chr3 195711406 N DEL 10
A00297:158:HT275DSXX:3:1116:18521:25958 chr3 195710595 N chr3 195711406 N DEL 10
A00404:155:HV27LDSXX:3:1676:7853:5040 chr3 195710459 N chr3 195711405 N DEL 19
A00297:158:HT275DSXX:3:1432:23764:20008 chr3 195710643 N chr3 195711409 N DEL 7
A00404:155:HV27LDSXX:3:2361:10547:23797 chr3 195710461 N chr3 195711407 N DEL 13
A00404:155:HV27LDSXX:4:1338:32018:12446 chr3 195710516 N chr3 195711417 N DEL 3
A00404:155:HV27LDSXX:4:2174:6126:6872 chr3 195710509 N chr3 195711410 N DEL 10
A00404:156:HV37TDSXX:1:2522:9390:31219 chr3 195711182 N chr3 195711453 N DEL 5
A00404:156:HV37TDSXX:1:2522:9941:32111 chr3 195711182 N chr3 195711453 N DEL 5
A00404:155:HV27LDSXX:1:2211:11867:7764 chr3 195711182 N chr3 195711453 N DEL 5
A00297:158:HT275DSXX:2:1559:31548:13103 chr3 195710642 N chr3 195711453 N DEL 20
A00297:158:HT275DSXX:2:2541:16658:29778 chr3 195711182 N chr3 195711453 N DEL 5
A00404:155:HV27LDSXX:4:1206:11216:20008 chr3 195711196 N chr3 195711467 N DEL 5
A00404:155:HV27LDSXX:3:1420:1434:34350 chr3 195710732 N chr3 195711453 N DEL 5
A00404:156:HV37TDSXX:3:2626:14850:3317 chr3 195711088 N chr3 195711523 N DUP 4
A00404:155:HV27LDSXX:3:1131:6777:22811 chr3 195710732 N chr3 195711453 N DEL 5
A00404:155:HV27LDSXX:2:2437:4679:35556 chr3 195710507 N chr3 195711453 N DEL 5
A00297:158:HT275DSXX:4:1604:1597:29277 chr3 195711088 N chr3 195711523 N DUP 5
A00404:156:HV37TDSXX:4:2119:32768:16626 chr3 195710520 N chr3 195711466 N DEL 5
A00404:155:HV27LDSXX:2:2535:6180:8500 chr3 195710507 N chr3 195711453 N DEL 5
A00297:158:HT275DSXX:2:1168:5412:34820 chr3 195710516 N chr3 195711462 N DEL 5
A00404:156:HV37TDSXX:4:2173:32081:22044 chr3 195711135 N chr3 195711572 N DEL 14
A00297:158:HT275DSXX:3:2268:9588:3975 chr3 195711132 N chr3 195711614 N DEL 8
A00404:156:HV37TDSXX:3:2601:3152:10488 chr3 195711132 N chr3 195711614 N DEL 6
A00297:158:HT275DSXX:4:2211:28646:1658 chr3 195711051 N chr3 195711578 N DEL 11
A00404:155:HV27LDSXX:3:2542:16947:20823 chr3 195711047 N chr3 195711574 N DEL 28
A00297:158:HT275DSXX:1:2625:28664:29434 chr3 195711047 N chr3 195711574 N DEL 23
A00297:158:HT275DSXX:2:2319:5132:15327 chr3 195711047 N chr3 195711574 N DEL 23
A00404:155:HV27LDSXX:4:2623:1416:35822 chr3 195711047 N chr3 195711574 N DEL 23
A00404:155:HV27LDSXX:3:2233:19334:28119 chr3 195710826 N chr3 195711623 N DEL 13
A00404:155:HV27LDSXX:2:1533:4453:36323 chr3 195710547 N chr3 195711614 N DEL 8
A00404:155:HV27LDSXX:4:1108:31467:8171 chr3 195711051 N chr3 195711578 N DEL 11
A00404:156:HV37TDSXX:2:2326:6822:18568 chr3 195710745 N chr3 195711587 N DEL 9
A00404:156:HV37TDSXX:2:1511:14579:32534 chr3 195710547 N chr3 195711614 N DEL 5
A00404:155:HV27LDSXX:3:2405:23755:35180 chr3 195710547 N chr3 195711614 N DEL 5
A00404:156:HV37TDSXX:3:1415:27697:3364 chr3 195710547 N chr3 195711614 N DEL 5
A00297:158:HT275DSXX:3:2216:16360:5368 chr3 195710547 N chr3 195711614 N DEL 5
A00297:158:HT275DSXX:3:2216:16378:5368 chr3 195710547 N chr3 195711614 N DEL 5
A00297:158:HT275DSXX:1:1233:18973:26209 chr3 195710547 N chr3 195711614 N DEL 5
A00404:156:HV37TDSXX:2:2511:16206:30718 chr3 195710547 N chr3 195711614 N DEL 5
A00404:155:HV27LDSXX:2:2119:31684:25081 chr3 195710547 N chr3 195711614 N DEL 5
A00297:158:HT275DSXX:3:2373:7491:23891 chr3 195710547 N chr3 195711614 N DEL 5
A00404:156:HV37TDSXX:4:2458:25807:20071 chr3 195710547 N chr3 195711614 N DEL 5
A00404:155:HV27LDSXX:3:2116:25608:25050 chr3 195710999 N chr3 195711616 N DEL 5
A00404:155:HV27LDSXX:3:2635:6171:16783 chr2 10200604 N chr2 10200853 N DEL 9
A00404:155:HV27LDSXX:3:2369:27742:11835 chr2 10200604 N chr2 10200853 N DEL 10
A00404:155:HV27LDSXX:4:2278:26937:11976 chr2 10200564 N chr2 10200625 N DUP 5
A00404:155:HV27LDSXX:2:1441:6234:13949 chr2 10200564 N chr2 10200625 N DUP 5
A00404:155:HV27LDSXX:2:1441:8187:16297 chr2 10200564 N chr2 10200625 N DUP 5
A00404:156:HV37TDSXX:2:2604:12364:9377 chr2 10200539 N chr2 10200631 N DUP 15
A00297:158:HT275DSXX:1:2245:17716:35775 chr2 10200607 N chr2 10200794 N DEL 31
A00404:155:HV27LDSXX:1:2203:14751:26850 chr2 10200554 N chr2 10200679 N DUP 14
A00404:156:HV37TDSXX:1:2433:30933:34961 chr2 10200554 N chr2 10200679 N DUP 19
A00404:155:HV27LDSXX:1:1161:32398:13041 chr2 10200658 N chr2 10200721 N DEL 5
A00297:158:HT275DSXX:3:1159:5267:2722 chr2 10200665 N chr2 10200728 N DEL 3
A00404:155:HV27LDSXX:4:2239:28411:32972 chr2 10200560 N chr2 10200747 N DEL 5
A00404:155:HV27LDSXX:2:2253:30409:31266 chr2 10200607 N chr2 10200794 N DEL 7
A00404:156:HV37TDSXX:2:1132:15745:28134 chr2 10200676 N chr2 10200799 N DEL 14
A00297:158:HT275DSXX:1:1416:29894:22764 chr2 10200710 N chr2 10200866 N DEL 10
A00297:158:HT275DSXX:2:1575:26856:1971 chr2 10200576 N chr2 10200794 N DEL 5
A00404:155:HV27LDSXX:3:1353:11650:1877 chr2 10200712 N chr2 10200868 N DEL 5
A00297:158:HT275DSXX:2:2621:19090:7279 chr2 10200712 N chr2 10200868 N DEL 5
A00404:155:HV27LDSXX:1:2149:3332:15875 chr2 10200712 N chr2 10200868 N DEL 5
A00404:155:HV27LDSXX:1:2149:5249:24455 chr2 10200712 N chr2 10200868 N DEL 5
A00404:155:HV27LDSXX:2:2362:16224:20791 chr2 10200588 N chr2 10200868 N DEL 5
A00404:156:HV37TDSXX:4:2577:10339:25254 chr2 10200586 N chr2 10200866 N DEL 7
A00404:155:HV27LDSXX:1:1428:12780:30733 chr3 8439721 N chr3 8439962 N DEL 2
A00404:156:HV37TDSXX:1:2377:16333:2816 chr3 8439775 N chr3 8439974 N DUP 3
A00404:156:HV37TDSXX:3:2145:27651:26209 chr3 8439618 N chr3 8440055 N DEL 2
A00297:158:HT275DSXX:1:1317:9498:29778 chr3 8439822 N chr3 8440142 N DEL 20
A00404:155:HV27LDSXX:1:1225:1967:28573 chr7 56151451 N chr7 56151626 N DUP 10
A00404:155:HV27LDSXX:2:2336:25654:34741 chr7 56151497 N chr7 56151623 N DUP 5
A00404:155:HV27LDSXX:2:2337:27498:4241 chr7 56151497 N chr7 56151623 N DUP 5
A00297:158:HT275DSXX:3:2340:2031:34882 chr7 56151504 N chr7 56151630 N DUP 5
A00404:155:HV27LDSXX:1:1440:31439:15546 chr7 56151568 N chr7 56151969 N DUP 5
A00404:155:HV27LDSXX:1:2669:25355:6104 chr7 56151412 N chr7 56151635 N DUP 4
A00404:155:HV27LDSXX:2:1122:16622:22701 chr7 56151616 N chr7 56151841 N DUP 2
A00297:158:HT275DSXX:3:2340:2031:34882 chr7 56151665 N chr7 56151842 N DUP 2
A00404:155:HV27LDSXX:2:1435:8648:25739 chr7 56151673 N chr7 56151899 N DUP 5
A00404:155:HV27LDSXX:3:1410:11785:16266 chr7 56151556 N chr7 56151732 N DEL 5
A00404:155:HV27LDSXX:3:2606:11966:22279 chr7 56151528 N chr7 56151704 N DEL 5
A00297:158:HT275DSXX:3:2607:29451:36025 chr7 56151528 N chr7 56151704 N DEL 5
A00404:155:HV27LDSXX:2:2336:25654:34741 chr7 56151528 N chr7 56151704 N DEL 5
A00297:158:HT275DSXX:4:2252:27932:9940 chr7 56151714 N chr7 56151940 N DUP 5
A00404:155:HV27LDSXX:4:2413:31033:9925 chr7 56151717 N chr7 56151943 N DUP 2
A00404:155:HV27LDSXX:2:2313:25229:26616 chr7 56151638 N chr7 56151863 N DUP 16
A00404:155:HV27LDSXX:2:2313:28971:31407 chr7 56151638 N chr7 56151863 N DUP 16
A00404:155:HV27LDSXX:4:2244:21703:4570 chr7 56151569 N chr7 56151892 N DUP 26
A00297:158:HT275DSXX:3:2456:10294:19852 chr7 56151477 N chr7 56151830 N DEL 15
A00404:155:HV27LDSXX:4:2659:3043:7639 chr7 56151474 N chr7 56151827 N DEL 7
A00404:156:HV37TDSXX:3:2338:5403:2394 chr7 56151602 N chr7 56151830 N DEL 10
A00404:155:HV27LDSXX:3:2167:10926:34194 chr7 56151838 N chr7 56152063 N DUP 5
A00297:158:HT275DSXX:3:2173:4797:16031 chr7 56151497 N chr7 56151851 N DEL 6
A00297:158:HT275DSXX:3:2173:9118:9486 chr7 56151497 N chr7 56151851 N DEL 6
A00297:158:HT275DSXX:4:1426:10556:6903 chr7 56151433 N chr7 56151836 N DEL 8
A00297:158:HT275DSXX:2:2657:21377:24017 chr7 56151497 N chr7 56151851 N DEL 5
A00404:155:HV27LDSXX:4:1524:14253:13150 chr7 56151828 N chr7 56152053 N DUP 3
A00404:155:HV27LDSXX:4:1524:15320:18223 chr7 56151828 N chr7 56152053 N DUP 3
A00297:158:HT275DSXX:3:2139:25934:34976 chr16 46385137 N chr16 46385252 N DEL 5
A00297:158:HT275DSXX:1:2232:31964:4304 chr16 46385045 N chr16 46385276 N DUP 2
A00404:156:HV37TDSXX:1:2154:26196:6026 chr16 46385175 N chr16 46385241 N DEL 5
A00404:156:HV37TDSXX:2:2406:11351:3270 chr16 46385135 N chr16 46385320 N DUP 1
A00404:156:HV37TDSXX:3:2464:22480:34538 chr16 46385074 N chr16 46385217 N DUP 5
A00404:155:HV27LDSXX:4:2261:3965:25394 chr16 46385248 N chr16 46385368 N DUP 5
A00404:155:HV27LDSXX:3:2170:19316:10457 chr16 46385309 N chr16 46385380 N DUP 5
A00404:156:HV37TDSXX:2:1654:29478:10113 chr16 46385067 N chr16 46385373 N DUP 5
A00404:156:HV37TDSXX:4:2559:29243:15154 chr16 46385099 N chr16 46385237 N DEL 3
A00297:158:HT275DSXX:3:2663:20292:6198 chr16 46385248 N chr16 46385368 N DUP 1
A00404:156:HV37TDSXX:3:1304:20085:1955 chr11 110890877 N chr11 110890948 N DEL 5
A00297:158:HT275DSXX:4:2139:31819:12602 chr11 110890877 N chr11 110890948 N DEL 5
A00297:158:HT275DSXX:4:1450:11252:21699 chr11 110890892 N chr11 110890947 N DEL 5
A00404:155:HV27LDSXX:4:1609:22878:1188 chr11 110890892 N chr11 110890947 N DEL 5
A00297:158:HT275DSXX:1:1302:4924:7670 chr11 110890892 N chr11 110890947 N DEL 11
A00404:156:HV37TDSXX:3:1558:13738:33677 chr11 110890892 N chr11 110890947 N DEL 15
A00404:156:HV37TDSXX:1:1536:4598:23202 chr11 110890743 N chr11 110890930 N DUP 15
A00404:155:HV27LDSXX:4:2257:18096:17049 chr11 110890701 N chr11 110890952 N DEL 11
A00404:155:HV27LDSXX:3:1158:15474:29575 chr11 110890702 N chr11 110890953 N DEL 10
A00297:158:HT275DSXX:4:1642:3378:25942 chr11 110890723 N chr11 110890956 N DEL 7
A00404:155:HV27LDSXX:1:1361:14525:26021 chr1 1944317 N chr1 1944394 N DEL 5
A00297:158:HT275DSXX:2:2363:12861:9267 chr11 62213191 N chr11 62213244 N DEL 12
A00404:156:HV37TDSXX:1:2274:18050:6261 chr13 27051988 N chr13 27052070 N DEL 7
A00404:156:HV37TDSXX:1:1133:10945:11772 chr13 27051972 N chr13 27052077 N DEL 7
A00404:155:HV27LDSXX:1:2430:22733:14497 chr13 27051973 N chr13 27052078 N DEL 7
A00297:158:HT275DSXX:3:1349:25843:35039 chr13 27051973 N chr13 27052078 N DEL 7
A00404:155:HV27LDSXX:2:1419:15682:15593 chr13 27051974 N chr13 27052079 N DEL 6
A00404:155:HV27LDSXX:3:2601:15772:28651 chr13 27051975 N chr13 27052080 N DEL 5
A00404:156:HV37TDSXX:3:2424:17056:33129 chr13 27052028 N chr13 27052093 N DEL 1
A00297:158:HT275DSXX:4:2268:26440:5384 chr1 232725423 N chr1 232725587 N DEL 7
A00404:156:HV37TDSXX:1:1554:11849:20760 chr1 232725423 N chr1 232725592 N DEL 7
A00404:156:HV37TDSXX:2:1557:22634:1799 chr12 132392041 N chr12 132392097 N DEL 4
A00297:158:HT275DSXX:4:1121:11035:12305 chr12 132392123 N chr12 132392210 N DEL 24
A00297:158:HT275DSXX:1:2564:28049:35164 chr12 132392171 N chr12 132392258 N DEL 14
A00297:158:HT275DSXX:4:1119:16984:34945 chr12 132392151 N chr12 132392637 N DEL 5
A00404:155:HV27LDSXX:4:1657:13602:26553 chr12 132392230 N chr12 132392714 N DUP 5
A00404:156:HV37TDSXX:4:2623:9598:26631 chr12 132392231 N chr12 132392715 N DUP 5
A00404:155:HV27LDSXX:1:2227:26973:35117 chr12 132392352 N chr12 132392410 N DEL 5
A00404:156:HV37TDSXX:4:2504:9860:35634 chr12 132392358 N chr12 132392728 N DUP 5
A00297:158:HT275DSXX:3:2172:25355:1251 chr12 132392074 N chr12 132392531 N DEL 5
A00297:158:HT275DSXX:3:2143:5611:16282 chr12 132392268 N chr12 132392668 N DEL 4
A00404:155:HV27LDSXX:1:2417:3938:23093 chr12 132392357 N chr12 132392756 N DEL 27
A00404:156:HV37TDSXX:1:2563:9191:17628 chrX 102738499 N chrX 102738713 N DEL 25
A00404:155:HV27LDSXX:3:1414:10194:32518 chr7 56371799 N chr7 56371946 N DEL 5
A00404:156:HV37TDSXX:3:2124:31087:5478 chr7 56371860 N chr7 56372041 N DEL 11
A00297:158:HT275DSXX:4:2573:27317:34178 chr7 56371809 N chr7 56371956 N DEL 5
A00297:158:HT275DSXX:2:1411:2239:9095 chr7 56371825 N chr7 56372005 N DEL 26
A00404:155:HV27LDSXX:4:1420:15899:23516 chr7 56371844 N chr7 56371940 N DUP 1
A00404:155:HV27LDSXX:2:2607:21603:27320 chr7 56371850 N chr7 56371947 N DUP 8
A00404:155:HV27LDSXX:1:1534:1958:5979 chr7 56371921 N chr7 56372053 N DEL 24
A00404:155:HV27LDSXX:1:1252:20211:8124 chr7 56371800 N chr7 56371896 N DUP 5
A00404:156:HV37TDSXX:4:1627:5367:9909 chr7 56371825 N chr7 56372005 N DEL 24
A00404:156:HV37TDSXX:4:1224:7256:33098 chr7 56371799 N chr7 56371946 N DEL 5
A00404:155:HV27LDSXX:3:2560:31873:35149 chr7 56371829 N chr7 56371927 N DEL 18
A00404:156:HV37TDSXX:2:1337:19723:7341 chr7 56371808 N chr7 56371906 N DEL 6
A00297:158:HT275DSXX:3:2305:8693:18270 chr7 56371799 N chr7 56371946 N DEL 5
A00404:156:HV37TDSXX:3:2619:18566:8844 chr7 56371871 N chr7 56372052 N DEL 8
A00404:155:HV27LDSXX:3:2116:23411:20462 chr7 56371839 N chr7 56371937 N DEL 5
A00404:156:HV37TDSXX:4:1241:25373:2566 chr7 56371830 N chr7 56371926 N DUP 2
A00404:156:HV37TDSXX:2:1109:11939:34914 chr7 56371823 N chr7 56371970 N DEL 5
A00404:156:HV37TDSXX:1:2127:17390:31203 chr7 56371834 N chr7 56371932 N DEL 5
A00404:156:HV37TDSXX:1:1540:16188:35540 chr7 56371848 N chr7 56371995 N DEL 5
A00404:156:HV37TDSXX:2:2212:13910:24111 chr7 56371799 N chr7 56371946 N DEL 18
A00404:156:HV37TDSXX:2:2103:18340:22608 chr7 56371810 N chr7 56371957 N DEL 4
A00404:156:HV37TDSXX:4:2316:6271:13730 chr7 56371823 N chr7 56371970 N DEL 35
A00404:156:HV37TDSXX:3:2447:25870:23625 chr7 56371799 N chr7 56371946 N DEL 38
A00404:155:HV27LDSXX:4:2646:19488:10191 chr7 56371832 N chr7 56371979 N DEL 5
A00404:156:HV37TDSXX:2:2372:22064:17691 chr7 56371793 N chr7 56372070 N DEL 5
A00404:156:HV37TDSXX:2:1359:18819:23625 chr7 56371805 N chr7 56371952 N DEL 9
A00404:156:HV37TDSXX:1:2424:28854:17550 chr7 56371824 N chr7 56371969 N DUP 5
A00404:155:HV27LDSXX:2:2565:10267:11537 chr7 56371836 N chr7 56371983 N DEL 5
A00404:156:HV37TDSXX:3:2117:23538:35681 chr1 22578850 N chr1 22579145 N DUP 5
A00297:158:HT275DSXX:3:2451:31467:29246 chr17 7077470 N chr17 7077683 N DEL 20
A00297:158:HT275DSXX:3:1476:25093:22122 chr17 7077470 N chr17 7077683 N DEL 20
A00404:155:HV27LDSXX:4:2110:10230:21778 chr17 7077444 N chr17 7077693 N DEL 20
A00404:155:HV27LDSXX:1:1341:31367:7216 chr17 7077470 N chr17 7077683 N DEL 20
A00404:155:HV27LDSXX:1:2340:32181:27539 chr17 7077470 N chr17 7077683 N DEL 20
A00297:158:HT275DSXX:1:1545:2157:16376 chr17 7077471 N chr17 7077684 N DEL 14
A00297:158:HT275DSXX:1:1622:11315:27352 chr8 63865366 N chr8 63865439 N DUP 36
A00404:155:HV27LDSXX:3:2551:13548:25081 chr8 63865366 N chr8 63865439 N DUP 40
A00404:156:HV37TDSXX:4:1166:25256:29888 chr8 63865366 N chr8 63865439 N DUP 45
A00404:155:HV27LDSXX:2:2107:25102:31313 chr8 63865366 N chr8 63865439 N DUP 48
A00404:155:HV27LDSXX:4:2338:32850:24846 chr8 63865366 N chr8 63865439 N DUP 38
A00297:158:HT275DSXX:1:2659:9552:30217 chr8 63865366 N chr8 63865439 N DUP 51
A00297:158:HT275DSXX:4:1224:21739:10645 chr8 63865363 N chr8 63865458 N DEL 7
A00404:156:HV37TDSXX:2:2635:1913:24189 chr17 17779923 N chr17 17780223 N DUP 12
A00404:155:HV27LDSXX:1:2454:11577:22514 chr17 17779942 N chr17 17780232 N DEL 15
A00404:155:HV27LDSXX:1:2248:31521:23171 chr7 142890263 N chr7 142890479 N DEL 30
A00404:155:HV27LDSXX:3:1574:26015:5838 chr7 142890263 N chr7 142890479 N DEL 41
A00404:156:HV37TDSXX:4:1234:3983:17127 chr7 142890274 N chr7 142890356 N DUP 9
A00404:156:HV37TDSXX:4:1475:24397:20948 chr7 142890274 N chr7 142890356 N DUP 9
A00297:158:HT275DSXX:3:1140:18728:1204 chr7 142890266 N chr7 142890706 N DEL 31
A00404:155:HV27LDSXX:2:2557:11541:33160 chr7 142890264 N chr7 142890394 N DUP 9
A00404:155:HV27LDSXX:2:2206:14841:2738 chr7 142890264 N chr7 142890394 N DUP 9
A00297:158:HT275DSXX:3:1369:5430:27023 chr7 142890264 N chr7 142890394 N DUP 9
A00404:155:HV27LDSXX:2:1256:28782:16767 chr7 142890264 N chr7 142890394 N DUP 9
A00297:158:HT275DSXX:3:1345:27679:13416 chr7 142890300 N chr7 142890416 N DUP 18
A00297:158:HT275DSXX:3:1462:27868:2190 chr7 142890278 N chr7 142890426 N DEL 2
A00297:158:HT275DSXX:1:1259:30346:3317 chr7 142890279 N chr7 142890427 N DEL 1
A00404:155:HV27LDSXX:3:2246:13051:4304 chr7 142890294 N chr7 142890424 N DEL 4
A00404:155:HV27LDSXX:3:2140:32850:22592 chr7 142890266 N chr7 142890552 N DUP 7
A00404:155:HV27LDSXX:4:1127:5602:28447 chr7 142890266 N chr7 142890552 N DUP 7
A00404:156:HV37TDSXX:1:2568:6198:6934 chr7 142890266 N chr7 142890552 N DUP 7
A00404:156:HV37TDSXX:1:2568:6262:7044 chr7 142890266 N chr7 142890552 N DUP 7
A00404:156:HV37TDSXX:2:1216:8513:11788 chr7 142890266 N chr7 142890552 N DUP 7
A00404:155:HV27LDSXX:4:1103:6108:15953 chr7 142890350 N chr7 142890484 N DEL 4
A00404:156:HV37TDSXX:4:2613:20952:29011 chr7 142890266 N chr7 142890552 N DUP 8
A00404:155:HV27LDSXX:4:2563:1814:25113 chr7 142890268 N chr7 142890616 N DUP 1
A00404:155:HV27LDSXX:4:2448:8278:25066 chr7 142890424 N chr7 142890555 N DEL 7
A00297:158:HT275DSXX:2:1278:13874:30624 chr7 142890310 N chr7 142890590 N DEL 18
A00297:158:HT275DSXX:2:2343:9426:27962 chr7 142890314 N chr7 142890594 N DEL 11
A00404:155:HV27LDSXX:1:1542:25708:33865 chr7 142890289 N chr7 142890639 N DEL 5
A00404:156:HV37TDSXX:3:2523:4607:28040 chr7 142890289 N chr7 142890639 N DEL 5
A00404:155:HV27LDSXX:1:1407:21576:6073 chr7 142890509 N chr7 142890764 N DUP 7
A00297:158:HT275DSXX:2:2170:12933:10927 chr7 142890509 N chr7 142890764 N DUP 7
A00404:155:HV27LDSXX:4:1618:32380:12915 chr7 142890509 N chr7 142890764 N DUP 7
A00404:155:HV27LDSXX:1:2554:24578:34663 chr7 142890509 N chr7 142890764 N DUP 7
A00404:156:HV37TDSXX:1:1243:8883:26209 chr7 142890397 N chr7 142890764 N DUP 12
A00404:156:HV37TDSXX:3:2523:4607:28040 chr7 142890354 N chr7 142890776 N DEL 6
A00404:156:HV37TDSXX:3:2653:14109:12962 chr7 142890346 N chr7 142890818 N DEL 16
A00404:155:HV27LDSXX:2:2308:29975:35994 chr7 142890293 N chr7 142890829 N DEL 4
A00404:155:HV27LDSXX:3:2543:29866:21026 chr7 142890356 N chr7 142890828 N DEL 5
A00404:156:HV37TDSXX:2:1304:16306:23563 chr7 142890498 N chr7 142890837 N DEL 6
A00404:156:HV37TDSXX:1:1642:26096:29465 chr7 142890279 N chr7 142890969 N DEL 6
A00404:156:HV37TDSXX:3:1565:29704:36495 chr7 142890279 N chr7 142890969 N DEL 6
A00297:158:HT275DSXX:3:1637:25943:21339 chr7 142890324 N chr7 142890968 N DEL 7
A00404:156:HV37TDSXX:2:2363:3287:26725 chr7 142890290 N chr7 142890980 N DEL 1
A00404:155:HV27LDSXX:3:2622:13277:24048 chr2 96461941 N chr2 96462241 N DUP 5
A00404:156:HV37TDSXX:4:2571:9616:7936 chr2 96461942 N chr2 96462242 N DUP 5
A00404:156:HV37TDSXX:2:2617:20528:14403 chr2 96462139 N chr2 96462265 N DUP 5
A00404:156:HV37TDSXX:2:2219:17815:25927 chr2 96462317 N chr2 96462416 N DEL 1
A00404:155:HV27LDSXX:1:1209:3784:33536 chr2 96461941 N chr2 96462339 N DUP 5
A00404:156:HV37TDSXX:2:1650:5764:26099 chr2 96462219 N chr2 96462316 N DUP 5
A00404:156:HV37TDSXX:3:2420:25744:27352 chr2 96462316 N chr2 96462544 N DEL 10
A00297:158:HT275DSXX:3:2508:26756:33802 chr2 96462219 N chr2 96462316 N DUP 5
A00404:155:HV27LDSXX:2:2354:10203:11397 chr2 96462219 N chr2 96462316 N DUP 5
A00404:156:HV37TDSXX:4:2130:4336:19899 chr2 96461961 N chr2 96462263 N DEL 5
A00404:156:HV37TDSXX:2:2650:14425:4805 chr2 96462219 N chr2 96462316 N DUP 5
A00297:158:HT275DSXX:4:2630:17861:28823 chr2 96462316 N chr2 96462544 N DEL 10
A00404:155:HV27LDSXX:1:1138:22679:26647 chr2 96462316 N chr2 96462544 N DEL 10
A00297:158:HT275DSXX:3:1234:20048:24251 chr2 96462465 N chr2 96462544 N DEL 18
A00297:158:HT275DSXX:2:1664:16803:4601 chr2 96462305 N chr2 96462404 N DEL 5
A00404:156:HV37TDSXX:3:2104:25581:36683 chr2 96461956 N chr2 96462355 N DEL 7
A00404:155:HV27LDSXX:3:2520:32696:25207 chr2 96462229 N chr2 96462377 N DEL 4
A00404:155:HV27LDSXX:4:1363:2148:33677 chr2 96462264 N chr2 96462413 N DEL 10
A00297:158:HT275DSXX:1:1514:17463:4993 chr2 96462256 N chr2 96462404 N DEL 5
A00404:156:HV37TDSXX:4:1311:22896:10050 chr2 96461961 N chr2 96462459 N DUP 5
A00404:156:HV37TDSXX:3:2427:11984:8187 chr2 96462096 N chr2 96462544 N DUP 2
A00404:155:HV27LDSXX:1:1147:11586:14982 chr2 96462302 N chr2 96462449 N DEL 7
A00404:156:HV37TDSXX:3:1572:7283:7592 chr2 96461963 N chr2 96462463 N DEL 7
A00404:156:HV37TDSXX:3:2427:11984:8187 chr2 96461957 N chr2 96462454 N DEL 7
A00297:158:HT275DSXX:1:2263:8386:6120 chr2 96462010 N chr2 96462510 N DEL 1
A00404:155:HV27LDSXX:1:2638:1913:21684 chr2 96462366 N chr2 96462543 N DUP 5
A00404:155:HV27LDSXX:4:1219:18132:5087 chr2 96462366 N chr2 96462543 N DUP 5
A00404:155:HV27LDSXX:1:1333:16116:24079 chr2 96462256 N chr2 96462582 N DEL 5
A00404:155:HV27LDSXX:4:1219:18132:5087 chr2 96462256 N chr2 96462582 N DEL 5
A00297:158:HT275DSXX:1:1510:2437:12602 chr2 96462218 N chr2 96462366 N DEL 5
A00404:156:HV37TDSXX:4:1671:30996:2942 chr2 96462257 N chr2 96462582 N DEL 12
A00297:158:HT275DSXX:3:2407:31593:33536 chr2 96462257 N chr2 96462582 N DEL 12
A00404:155:HV27LDSXX:2:2338:6325:31861 chr2 96462113 N chr2 96462563 N DEL 5
A00404:156:HV37TDSXX:2:1176:27462:6151 chr2 96462448 N chr2 96462624 N DUP 6
A00404:156:HV37TDSXX:3:2144:2465:2660 chr2 96461914 N chr2 96462641 N DEL 1
A00404:155:HV27LDSXX:3:2331:21224:18834 chr2 96462620 N chr2 96462672 N DEL 7
A00404:156:HV37TDSXX:1:1353:27398:36511 chr4 38162007 N chr4 38162145 N DEL 4
A00404:156:HV37TDSXX:2:2510:22833:28354 chr20 25220612 N chr20 25220672 N DEL 55
A00404:156:HV37TDSXX:1:1522:27850:9204 chr22 10572398 N chr22 10572543 N DUP 12
A00404:156:HV37TDSXX:1:1522:28709:8907 chr22 10572398 N chr22 10572543 N DUP 12
A00297:158:HT275DSXX:4:1417:13548:35697 chr13 33685181 N chr13 33685363 N DEL 5
A00297:158:HT275DSXX:2:1566:3459:22482 chr13 33685181 N chr13 33685363 N DEL 5
A00404:156:HV37TDSXX:3:1518:21305:30467 chr13 33685181 N chr13 33685363 N DEL 5
A00297:158:HT275DSXX:2:2249:21567:26036 chr2 69902780 N chr2 69902869 N DUP 1
A00404:155:HV27LDSXX:3:2211:31286:30405 chr2 69902780 N chr2 69902869 N DUP 1
A00297:158:HT275DSXX:4:1548:18204:27790 chr1 231011289 N chr1 231011368 N DUP 6
A00297:158:HT275DSXX:2:1335:7844:5368 chr1 231011289 N chr1 231011368 N DUP 8
A00297:158:HT275DSXX:4:2334:16396:17394 chr1 231011378 N chr1 231011497 N DUP 1
A00404:155:HV27LDSXX:1:1621:26639:2315 chr1 231011346 N chr1 231011509 N DUP 2
A00297:158:HT275DSXX:2:2504:13928:1877 chr22 39596329 N chr22 39596453 N DEL 5
A00404:156:HV37TDSXX:2:2414:6732:22670 chr22 39596320 N chr22 39596508 N DUP 23
A00404:156:HV37TDSXX:2:2414:7934:21183 chr22 39596320 N chr22 39596508 N DUP 18
A00404:156:HV37TDSXX:4:2462:25825:6668 chr22 39596320 N chr22 39596508 N DUP 20
A00404:156:HV37TDSXX:2:2235:29622:21887 chr22 39596431 N chr22 39596500 N DEL 16
A00404:155:HV27LDSXX:4:1463:1850:22983 chr22 39596423 N chr22 39596492 N DEL 19
A00404:155:HV27LDSXX:1:2628:14977:13745 chr22 39596423 N chr22 39596492 N DEL 28
A00404:155:HV27LDSXX:4:1278:2419:11443 chr22 39596464 N chr22 39596602 N DEL 31
A00404:156:HV37TDSXX:2:1530:4291:29622 chr22 39596423 N chr22 39596492 N DEL 19
A00404:155:HV27LDSXX:2:1230:13584:24706 chr22 39596289 N chr22 39596619 N DEL 1
A00404:155:HV27LDSXX:1:1465:28248:25582 chr22 39596615 N chr22 39596707 N DEL 39
A00297:158:HT275DSXX:2:1523:20030:30890 chr22 39596347 N chr22 39596676 N DEL 3
A00297:158:HT275DSXX:2:1611:22525:5368 chr6 160789269 N chr6 160789643 N DEL 5
A00404:156:HV37TDSXX:1:2564:23448:23657 chr6 160789269 N chr6 160789643 N DEL 5
A00297:158:HT275DSXX:4:1576:4978:25332 chr6 160789290 N chr6 160790110 N DEL 1
A00404:156:HV37TDSXX:1:2405:27498:28197 chr6 160789232 N chr6 160789357 N DUP 1
A00404:156:HV37TDSXX:4:2508:6063:11584 chr6 160789488 N chr6 160789843 N DEL 3
A00404:155:HV27LDSXX:3:1655:5846:24298 chr6 160789301 N chr6 160789390 N DEL 1
A00297:158:HT275DSXX:1:2104:23520:15859 chr6 160789580 N chr6 160790107 N DEL 5
A00404:156:HV37TDSXX:3:2325:16360:22216 chr6 160789580 N chr6 160790107 N DEL 5
A00404:155:HV27LDSXX:1:1602:23231:3239 chr6 160789580 N chr6 160790107 N DEL 5
A00404:156:HV37TDSXX:1:1150:16504:11537 chr6 160789580 N chr6 160790107 N DEL 5
A00404:155:HV27LDSXX:1:1102:19714:22733 chr6 160789580 N chr6 160790107 N DEL 5
A00297:158:HT275DSXX:2:1611:22525:5368 chr6 160789596 N chr6 160790121 N DUP 5
A00297:158:HT275DSXX:4:2218:1796:2816 chr6 160789305 N chr6 160789599 N DEL 4
A00404:156:HV37TDSXX:1:1168:17300:19805 chr6 160789314 N chr6 160789608 N DEL 2
A00404:155:HV27LDSXX:2:2644:31566:13917 chr6 160789736 N chr6 160789934 N DEL 5
A00404:156:HV37TDSXX:3:2166:20094:17942 chr6 160789370 N chr6 160789735 N DUP 5
A00297:158:HT275DSXX:3:1521:31991:1532 chr6 160789900 N chr6 160790029 N DEL 4
A00404:156:HV37TDSXX:2:1426:21576:20666 chr6 160789900 N chr6 160790029 N DEL 5
A00404:156:HV37TDSXX:1:2314:25654:15890 chr6 160789900 N chr6 160790029 N DEL 5
A00297:158:HT275DSXX:1:2569:28293:18114 chr6 160789900 N chr6 160790029 N DEL 5
A00404:156:HV37TDSXX:2:1637:29107:31140 chr6 160789924 N chr6 160790051 N DUP 5
A00404:155:HV27LDSXX:2:1115:20265:15421 chr6 160789312 N chr6 160789924 N DEL 5
A00404:155:HV27LDSXX:2:2536:21477:26193 chr6 160790034 N chr6 160790154 N DUP 13
A00404:156:HV37TDSXX:3:1530:5132:11412 chr6 160789990 N chr6 160790155 N DUP 12
A00297:158:HT275DSXX:1:1672:30915:10160 chr6 160789990 N chr6 160790155 N DUP 12
A00404:155:HV27LDSXX:1:1132:16504:4867 chr6 160789990 N chr6 160790155 N DUP 12
A00404:155:HV27LDSXX:1:1132:18132:4586 chr6 160789990 N chr6 160790155 N DUP 12
A00297:158:HT275DSXX:2:1625:25672:14011 chr6 160789990 N chr6 160790155 N DUP 12
A00404:155:HV27LDSXX:4:1228:26431:31234 chr6 160789990 N chr6 160790155 N DUP 12
A00297:158:HT275DSXX:1:1569:9887:1705 chr6 160789251 N chr6 160790150 N DEL 7
A00404:155:HV27LDSXX:3:1336:25699:11397 chr6 160790047 N chr6 160790213 N DEL 5
A00297:158:HT275DSXX:2:2556:16613:29074 chr6 160789309 N chr6 160790214 N DEL 5
A00297:158:HT275DSXX:1:2547:24740:13557 chr6 160789309 N chr6 160790214 N DEL 5
A00404:155:HV27LDSXX:4:2519:24288:36417 chr6 160789311 N chr6 160790216 N DEL 5
A00404:156:HV37TDSXX:3:1155:28293:33176 chr6 160789241 N chr6 160790226 N DEL 2
A00404:156:HV37TDSXX:2:1536:27398:21355 chr9 137355584 N chr9 137355763 N DEL 5
A00297:158:HT275DSXX:3:1415:10529:33223 chr9 137355584 N chr9 137355763 N DEL 10
A00404:155:HV27LDSXX:1:1404:17698:26788 chr9 137355611 N chr9 137355790 N DEL 6
A00297:158:HT275DSXX:1:2438:8721:25676 chr9 137355627 N chr9 137355828 N DEL 11
A00297:158:HT275DSXX:3:2358:20717:12352 chr9 137355627 N chr9 137355828 N DEL 14
A00297:158:HT275DSXX:1:1254:29478:12148 chr9 137355623 N chr9 137355723 N DEL 12
A00404:156:HV37TDSXX:2:1677:8368:11350 chr9 137355620 N chr9 137355720 N DEL 17
A00404:156:HV37TDSXX:2:1677:9191:11929 chr9 137355620 N chr9 137355720 N DEL 17
A00404:156:HV37TDSXX:4:1153:31033:21198 chr9 137355620 N chr9 137355720 N DEL 17
A00297:158:HT275DSXX:2:2630:8359:14528 chr9 137355620 N chr9 137355720 N DEL 17
A00297:158:HT275DSXX:3:2532:2013:18818 chr9 137355627 N chr9 137355828 N DEL 21
A00404:155:HV27LDSXX:1:1655:15609:2754 chr9 137355564 N chr9 137355613 N DUP 9
A00404:155:HV27LDSXX:2:1570:15546:36432 chr9 137355584 N chr9 137355763 N DEL 13
A00297:158:HT275DSXX:2:1103:27398:10802 chr9 137355584 N chr9 137355763 N DEL 13
A00297:158:HT275DSXX:2:1103:27606:10786 chr9 137355584 N chr9 137355763 N DEL 13
A00404:155:HV27LDSXX:4:1619:25717:8797 chr9 137355620 N chr9 137355720 N DEL 20
A00404:156:HV37TDSXX:3:1532:10194:2581 chr9 137355620 N chr9 137355720 N DEL 10
A00404:155:HV27LDSXX:1:2176:12735:15749 chr9 137355620 N chr9 137355720 N DEL 10
A00297:158:HT275DSXX:4:2569:14118:27070 chr9 137355600 N chr9 137355812 N DUP 22
A00297:158:HT275DSXX:4:2453:2022:21684 chr9 137355618 N chr9 137355687 N DUP 4
A00404:155:HV27LDSXX:1:2251:19289:2613 chr9 137355578 N chr9 137355655 N DUP 1
A00404:155:HV27LDSXX:4:2318:8178:23829 chr9 137355578 N chr9 137355655 N DUP 1
A00404:155:HV27LDSXX:3:2170:30065:2769 chr9 137355602 N chr9 137355651 N DUP 17
A00404:155:HV27LDSXX:4:1139:22390:30436 chr9 137355755 N chr9 137355883 N DUP 21
A00404:156:HV37TDSXX:2:2156:23366:27680 chr9 137355745 N chr9 137355866 N DUP 45
A00404:155:HV27LDSXX:2:2345:25120:28933 chr9 137355633 N chr9 137355695 N DUP 16
A00404:155:HV27LDSXX:2:2366:20311:22827 chr9 137355568 N chr9 137355680 N DUP 11
A00404:155:HV27LDSXX:2:2363:8160:8766 chr9 137355600 N chr9 137355741 N DUP 17
A00404:155:HV27LDSXX:4:2128:7672:7451 chr9 137355617 N chr9 137355837 N DUP 18
A00297:158:HT275DSXX:2:2214:15691:21527 chr9 137355821 N chr9 137355877 N DUP 23
A00297:158:HT275DSXX:3:1450:12653:26381 chr9 137355711 N chr9 137355835 N DEL 13
A00404:155:HV27LDSXX:1:2264:20482:14043 chr9 137355612 N chr9 137355854 N DUP 18
A00297:158:HT275DSXX:4:1438:6668:16172 chr9 137355628 N chr9 137355705 N DUP 30
A00404:156:HV37TDSXX:1:2648:15573:21950 chr9 137355564 N chr9 137355613 N DUP 16
A00297:158:HT275DSXX:2:2153:12192:14998 chr9 137355600 N chr9 137355820 N DUP 20
A00404:155:HV27LDSXX:4:2454:12979:10942 chr9 137355612 N chr9 137355796 N DUP 13
A00404:156:HV37TDSXX:4:1628:1497:19053 chr9 137355600 N chr9 137355834 N DUP 23
A00297:158:HT275DSXX:2:1266:25382:12947 chr9 137355600 N chr9 137355870 N DUP 16
A00404:156:HV37TDSXX:4:1157:24460:6558 chr9 137355619 N chr9 137355688 N DUP 24
A00404:155:HV27LDSXX:1:2264:20482:14043 chr9 137355821 N chr9 137355877 N DUP 30
A00404:155:HV27LDSXX:2:2161:15275:9408 chr9 137355697 N chr9 137355778 N DEL 14
A00297:158:HT275DSXX:4:2320:9236:8844 chr9 137355601 N chr9 137355742 N DUP 7
A00297:158:HT275DSXX:1:1439:9462:33285 chr9 137355687 N chr9 137355823 N DUP 15
A00404:156:HV37TDSXX:2:2623:22652:22122 chr9 137355631 N chr9 137355837 N DUP 15
A00404:155:HV27LDSXX:4:2219:28926:5995 chr9 137355601 N chr9 137355742 N DUP 8
A00404:155:HV27LDSXX:4:1358:13503:7780 chr9 137355674 N chr9 137355754 N DEL 15
A00297:158:HT275DSXX:2:1657:23619:5697 chr9 137355564 N chr9 137355662 N DUP 16
A00404:155:HV27LDSXX:2:2220:5855:23500 chr9 137355621 N chr9 137355741 N DUP 12
A00404:155:HV27LDSXX:2:2220:6253:21245 chr9 137355621 N chr9 137355741 N DUP 12
A00297:158:HT275DSXX:2:1504:18132:29481 chr9 137355614 N chr9 137355820 N DUP 17
A00297:158:HT275DSXX:2:1505:17960:34287 chr9 137355614 N chr9 137355820 N DUP 17
A00297:158:HT275DSXX:2:1505:17978:34256 chr9 137355614 N chr9 137355820 N DUP 17
A00404:155:HV27LDSXX:4:1336:20021:5885 chr9 137355614 N chr9 137355712 N DUP 13
A00297:158:HT275DSXX:1:2332:5041:11099 chr9 137355733 N chr9 137355828 N DEL 21
A00404:155:HV27LDSXX:4:1358:13503:7780 chr9 137355677 N chr9 137355762 N DUP 15
A00404:156:HV37TDSXX:2:2543:6632:3959 chr9 137355733 N chr9 137355828 N DEL 21
A00404:155:HV27LDSXX:1:2639:16378:32487 chr9 137355745 N chr9 137355866 N DUP 45
A00297:158:HT275DSXX:2:2307:12029:4445 chr9 137355711 N chr9 137355828 N DEL 15
A00404:155:HV27LDSXX:3:2254:14705:22138 chr9 137355593 N chr9 137355726 N DUP 21
A00404:155:HV27LDSXX:1:1678:7129:20322 chr9 137355747 N chr9 137355882 N DUP 29
A00404:155:HV27LDSXX:3:2459:32108:27352 chr9 137355716 N chr9 137355782 N DEL 17
A00404:155:HV27LDSXX:1:2361:4056:23735 chr9 137355698 N chr9 137355785 N DEL 37
A00404:155:HV27LDSXX:2:2345:22498:22858 chr9 137355600 N chr9 137355820 N DUP 11
A00404:155:HV27LDSXX:1:2659:27308:26929 chr9 137355733 N chr9 137355828 N DEL 15
A00297:158:HT275DSXX:4:2321:10999:15436 chr9 137355677 N chr9 137355762 N DUP 22
A00297:158:HT275DSXX:4:1675:3965:16783 chr9 137355677 N chr9 137355849 N DUP 12
A00404:156:HV37TDSXX:4:2227:4869:10551 chr9 137355704 N chr9 137355828 N DEL 26
A00297:158:HT275DSXX:3:2250:27624:5869 chr9 137355715 N chr9 137355853 N DEL 22
A00404:155:HV27LDSXX:2:1145:29758:5776 chr9 137355662 N chr9 137355828 N DEL 16
A00297:158:HT275DSXX:2:1658:4336:36464 chr9 137355670 N chr9 137355836 N DEL 16
A00297:158:HT275DSXX:2:2660:1479:1172 chr9 137355670 N chr9 137355836 N DEL 16
A00297:158:HT275DSXX:1:2502:3848:15389 chr9 137355740 N chr9 137355806 N DEL 5
A00404:156:HV37TDSXX:1:2439:9109:32894 chr9 137355733 N chr9 137355871 N DEL 18
A00404:156:HV37TDSXX:2:1426:9155:34194 chr9 137355634 N chr9 137355828 N DEL 21
A00404:156:HV37TDSXX:2:1426:9805:33692 chr9 137355634 N chr9 137355828 N DEL 21
A00404:155:HV27LDSXX:3:2167:17463:4492 chr9 137355634 N chr9 137355828 N DEL 21
A00404:156:HV37TDSXX:2:2454:17354:20212 chr9 137355634 N chr9 137355828 N DEL 20
A00297:158:HT275DSXX:2:1339:24325:20697 chr9 137355634 N chr9 137355828 N DEL 18
A00297:158:HT275DSXX:1:2634:26784:23516 chr9 137355634 N chr9 137355828 N DEL 16
A00404:155:HV27LDSXX:2:1536:21350:18051 chr9 137355634 N chr9 137355828 N DEL 16
A00404:156:HV37TDSXX:2:1408:9815:15452 chr9 137355634 N chr9 137355828 N DEL 15
A00297:158:HT275DSXX:1:2502:3848:15389 chr9 137355655 N chr9 137355843 N DEL 11
A00297:158:HT275DSXX:1:1263:5258:36839 chr9 137355676 N chr9 137355857 N DEL 19
A00404:155:HV27LDSXX:3:1261:15004:34585 chr6 31068210 N chr6 31068287 N DEL 5
A00404:156:HV37TDSXX:3:2421:22010:34006 chr6 31068343 N chr6 31068407 N DEL 14
A00404:155:HV27LDSXX:3:1221:17933:17550 chr6 31068343 N chr6 31068407 N DEL 14
A00404:155:HV27LDSXX:4:1163:29225:31250 chr6 31068344 N chr6 31068408 N DEL 14
A00404:156:HV37TDSXX:1:1157:25093:2550 chr11 71090237 N chr11 71090507 N DEL 9
A00404:155:HV27LDSXX:3:1174:13838:23547 chr11 71090237 N chr11 71090600 N DEL 13
A00297:158:HT275DSXX:2:2143:24876:29512 chr11 71090320 N chr11 71090499 N DEL 3
A00404:155:HV27LDSXX:4:1310:13865:24032 chr11 71090320 N chr11 71090499 N DEL 3
A00404:156:HV37TDSXX:1:2111:20591:33896 chr11 71090320 N chr11 71090499 N DEL 3
A00404:156:HV37TDSXX:4:2602:2926:4679 chr11 71090246 N chr11 71090334 N DEL 6
A00404:156:HV37TDSXX:1:2342:27715:29074 chr11 71090412 N chr11 71090591 N DUP 15
A00404:156:HV37TDSXX:1:2342:28537:30217 chr11 71090412 N chr11 71090591 N DUP 15
A00404:156:HV37TDSXX:1:1268:31403:16517 chr11 71090412 N chr11 71090591 N DUP 12
A00404:155:HV27LDSXX:3:1174:13838:23547 chr11 71090240 N chr11 71090413 N DEL 25
A00404:156:HV37TDSXX:4:2301:12391:3630 chr11 71090417 N chr11 71090592 N DEL 9
A00297:158:HT275DSXX:1:1228:26458:35258 chr11 71090248 N chr11 71090441 N DUP 13
A00404:155:HV27LDSXX:3:1577:17897:24878 chr11 71090341 N chr11 71090690 N DEL 31
A00404:156:HV37TDSXX:1:1157:25093:2550 chr11 71090421 N chr11 71090600 N DUP 15
A00297:158:HT275DSXX:2:2139:10836:10019 chr11 71090412 N chr11 71090591 N DUP 20
A00404:155:HV27LDSXX:4:1461:21621:32737 chr11 71090341 N chr11 71090690 N DEL 31
A00404:155:HV27LDSXX:3:1135:3179:12508 chr11 71090502 N chr11 71090592 N DEL 27
A00404:156:HV37TDSXX:1:2664:9778:24502 chr11 71090341 N chr11 71090690 N DEL 31
A00404:156:HV37TDSXX:4:2261:26539:3897 chr11 71090515 N chr11 71090690 N DEL 32
A00404:156:HV37TDSXX:4:1323:32199:7842 chr11 71090341 N chr11 71090690 N DEL 31
A00404:155:HV27LDSXX:3:2554:17300:13291 chr11 71090515 N chr11 71090690 N DEL 28
A00404:156:HV37TDSXX:4:2506:10936:3270 chr11 71090392 N chr11 71090478 N DUP 9
A00404:155:HV27LDSXX:3:1377:3134:11584 chr11 71090500 N chr11 71090592 N DEL 6
A00404:156:HV37TDSXX:1:2374:20437:28244 chr11 71090428 N chr11 71090690 N DEL 30
A00404:155:HV27LDSXX:4:1412:19976:13416 chr11 71090691 N chr11 71090775 N DEL 11
A00297:158:HT275DSXX:2:2139:10836:10019 chr11 71090414 N chr11 71090775 N DEL 9
A00297:158:HT275DSXX:4:1173:23095:30843 chr11 71090414 N chr11 71090775 N DEL 9
A00404:155:HV27LDSXX:4:1459:26802:18537 chr11 71090414 N chr11 71090775 N DEL 9
A00404:155:HV27LDSXX:2:2459:11831:22106 chr11 71090412 N chr11 71090779 N DEL 9
A00297:158:HT275DSXX:4:1247:13584:25144 chr11 71090414 N chr11 71090775 N DEL 9
A00297:158:HT275DSXX:1:1203:4788:2895 chr11 71090414 N chr11 71090775 N DEL 9
A00404:156:HV37TDSXX:1:1240:14507:30655 chr11 71090414 N chr11 71090775 N DEL 9
A00404:156:HV37TDSXX:1:2635:7157:5556 chr11 71090414 N chr11 71090781 N DEL 9
A00404:156:HV37TDSXX:3:2219:30499:30702 chr11 71090414 N chr11 71090781 N DEL 9
A00404:155:HV27LDSXX:4:1509:12617:32737 chr11 71090415 N chr11 71090782 N DEL 9
A00404:155:HV27LDSXX:4:1509:12789:32690 chr11 71090415 N chr11 71090782 N DEL 9
A00404:156:HV37TDSXX:3:1616:28384:11193 chr11 71090420 N chr11 71090787 N DEL 7
A00404:155:HV27LDSXX:2:2337:19316:16470 chr19 18829591 N chr19 18829674 N DEL 4
A00297:158:HT275DSXX:4:2342:27787:24314 chr8 18412022 N chr8 18412225 N DEL 5
A00404:156:HV37TDSXX:2:1247:28040:19085 chr12 5812632 N chr12 5812897 N DEL 7
A00297:158:HT275DSXX:1:2632:10041:32659 chr12 5812470 N chr12 5812646 N DUP 5
A00297:158:HT275DSXX:1:1534:29677:25864 chr12 5812834 N chr12 5813149 N DEL 1
A00297:158:HT275DSXX:4:2549:10484:18302 chr12 5812834 N chr12 5813149 N DEL 1
A00404:156:HV37TDSXX:1:2225:10465:34773 chr12 5812731 N chr12 5812835 N DUP 2
A00297:158:HT275DSXX:2:1653:6198:20055 chr12 5812739 N chr12 5812845 N DUP 14
A00297:158:HT275DSXX:1:1362:30915:22498 chr12 5812724 N chr12 5813148 N DUP 9
A00404:155:HV27LDSXX:2:2305:24957:31219 chr12 5812623 N chr12 5813222 N DUP 11
A00297:158:HT275DSXX:3:1421:10954:12853 chr19 50544236 N chr19 50544537 N DEL 40
A00404:156:HV37TDSXX:2:2128:28809:20228 chr19 50544116 N chr19 50544418 N DEL 5
A00297:158:HT275DSXX:4:2561:24334:8281 chr19 50544012 N chr19 50544668 N DEL 4
A00404:155:HV27LDSXX:3:1314:3278:6355 chr1 152475895 N chr1 152476035 N DEL 29
A00297:158:HT275DSXX:2:1409:2094:5212 chr11 111358734 N chr11 111358847 N DUP 9
A00404:156:HV37TDSXX:4:1638:27733:6214 chr11 111358734 N chr11 111358847 N DUP 9
A00404:156:HV37TDSXX:1:2359:27028:3771 chr10 507336 N chr10 507466 N DEL 5
A00404:156:HV37TDSXX:1:1645:2248:9643 chr10 507375 N chr10 507595 N DEL 24
A00404:155:HV27LDSXX:2:2436:11098:28855 chr10 507417 N chr10 507637 N DEL 12
A00297:158:HT275DSXX:3:2577:22037:5932 chr10 507363 N chr10 507665 N DUP 2
A00404:155:HV27LDSXX:1:2419:31864:7639 chr10 507396 N chr10 507487 N DEL 16
A00297:158:HT275DSXX:2:1627:8802:34397 chr10 507317 N chr10 507537 N DEL 5
A00404:156:HV37TDSXX:1:2321:23294:31563 chr10 507330 N chr10 507550 N DEL 4
A00404:155:HV27LDSXX:3:1325:4381:12649 chrX 53891881 N chrX 53891953 N DEL 5
A00297:158:HT275DSXX:3:1168:22598:28260 chr11 120347348 N chr11 120347399 N DUP 9
A00297:158:HT275DSXX:4:1230:29279:14090 chr10 28262354 N chr10 28262417 N DEL 17
A00404:155:HV27LDSXX:4:1274:15492:24189 chr12 121993895 N chr12 121994252 N DEL 1
A00297:158:HT275DSXX:1:1513:19452:19586 chr12 121993858 N chr12 121994218 N DEL 65
A00297:158:HT275DSXX:2:2639:11595:21230 chr12 121993895 N chr12 121994252 N DEL 12
A00404:155:HV27LDSXX:2:2230:10149:13244 chr12 121993895 N chr12 121994252 N DEL 12
A00297:158:HT275DSXX:1:1111:1298:34334 chr12 121993895 N chr12 121994381 N DEL 11
A00404:156:HV37TDSXX:1:1315:5394:22608 chr12 121993926 N chr12 121994281 N DUP 5
A00404:155:HV27LDSXX:3:2419:30210:14387 chr12 121994013 N chr12 121994499 N DUP 6
A00404:156:HV37TDSXX:2:1439:18213:14121 chr12 121994030 N chr12 121994210 N DEL 5
A00297:158:HT275DSXX:1:2525:2908:2143 chr12 121994209 N chr12 121994339 N DEL 5
A00297:158:HT275DSXX:2:1667:8314:32957 chr12 121993998 N chr12 121994306 N DUP 7
A00404:156:HV37TDSXX:2:2519:24560:11741 chr12 121993981 N chr12 121994417 N DUP 2
A00297:158:HT275DSXX:1:2527:10131:12242 chr12 121994240 N chr12 121994370 N DEL 9
A00404:155:HV27LDSXX:4:1148:11776:13870 chr12 121993994 N chr12 121994302 N DUP 7
A00404:156:HV37TDSXX:3:1659:21224:27602 chr12 121993994 N chr12 121994299 N DUP 7
A00404:156:HV37TDSXX:4:2656:9977:8594 chr12 121994075 N chr12 121994255 N DEL 1
A00297:158:HT275DSXX:2:1522:18222:23594 chr12 121994079 N chr12 121994259 N DEL 1
A00297:158:HT275DSXX:4:1601:18231:25113 chr12 121993975 N chr12 121994284 N DEL 1
A00404:156:HV37TDSXX:1:1275:1118:19523 chr12 121993994 N chr12 121994302 N DEL 7
A00404:156:HV37TDSXX:1:1435:27905:32440 chr12 121994186 N chr12 121994316 N DEL 1
A00297:158:HT275DSXX:1:1251:4833:34194 chr1 242733851 N chr1 242733912 N DUP 15
A00297:158:HT275DSXX:1:1251:5448:32534 chr1 242733851 N chr1 242733912 N DUP 15
A00297:158:HT275DSXX:1:1439:9697:33755 chr1 242733851 N chr1 242733912 N DUP 15
A00404:156:HV37TDSXX:2:1602:19009:22232 chr1 242733851 N chr1 242733912 N DUP 15
A00404:156:HV37TDSXX:2:1602:19063:21605 chr1 242733851 N chr1 242733912 N DUP 15
A00404:156:HV37TDSXX:3:1427:29957:28541 chr1 242733851 N chr1 242733912 N DUP 15
A00404:156:HV37TDSXX:4:2133:10122:19586 chr1 242733851 N chr1 242733912 N DUP 15
A00404:155:HV27LDSXX:3:1317:20889:36479 chr1 242733851 N chr1 242733912 N DUP 15
A00297:158:HT275DSXX:2:2315:21847:22921 chr11 71124354 N chr11 71124426 N DEL 5
A00404:155:HV27LDSXX:4:1503:14525:33473 chr7 105558807 N chr7 105558942 N DUP 3
A00297:158:HT275DSXX:4:2114:27326:19163 chr2 112720052 N chr2 112720125 N DUP 8
A00297:158:HT275DSXX:3:1219:20455:2127 chr2 112720055 N chr2 112720124 N DEL 5
A00297:158:HT275DSXX:3:2677:20618:35728 chr2 112720067 N chr2 112720138 N DEL 1
A00297:158:HT275DSXX:1:1570:31458:4085 chr16 54302269 N chr16 54302462 N DUP 1
A00404:155:HV27LDSXX:1:2203:2193:32127 chr4 65574749 N chr4 65574882 N DEL 9
A00404:155:HV27LDSXX:4:2475:2338:1658 chr4 65574817 N chr4 65574878 N DUP 7
A00297:158:HT275DSXX:3:2102:20383:9111 chr4 65574782 N chr4 65574863 N DEL 6
A00297:158:HT275DSXX:2:2228:3115:2879 chr4 65574787 N chr4 65574868 N DEL 4
A00404:155:HV27LDSXX:2:1118:24523:19507 chr4 65574840 N chr4 65574893 N DEL 10
A00404:156:HV37TDSXX:1:1616:6786:23610 chr4 65574774 N chr4 65574903 N DEL 5
A00404:156:HV37TDSXX:1:1616:6949:22701 chr4 65574774 N chr4 65574903 N DEL 5
A00404:156:HV37TDSXX:4:2446:28293:14512 chr4 65574775 N chr4 65574904 N DEL 4
A00404:156:HV37TDSXX:4:2578:20573:14700 chr5 64225962 N chr5 64226122 N DUP 9
A00297:158:HT275DSXX:1:1325:19397:28667 chr3 130085447 N chr3 130085587 N DUP 10
A00404:156:HV37TDSXX:4:2432:32560:30483 chr3 130085447 N chr3 130085587 N DUP 10
A00404:155:HV27LDSXX:3:1159:19000:9659 chr3 130085469 N chr3 130085611 N DEL 12
A00404:156:HV37TDSXX:1:2272:13593:16736 chr3 130085469 N chr3 130085611 N DEL 10
A00404:156:HV37TDSXX:1:2272:15085:16219 chr3 130085469 N chr3 130085611 N DEL 10
A00404:156:HV37TDSXX:3:1264:30581:14278 chr3 130085473 N chr3 130085615 N DEL 5
A00404:155:HV27LDSXX:1:1266:14913:28009 chr3 130085482 N chr3 130085624 N DEL 2
A00297:158:HT275DSXX:2:1413:18322:29058 chr3 130085521 N chr3 130085663 N DEL 5
A00404:156:HV37TDSXX:1:2509:4797:6042 chr2 33776018 N chr2 33776138 N DEL 5
A00297:158:HT275DSXX:1:2267:20961:6104 chr2 33776018 N chr2 33776138 N DEL 5
A00297:158:HT275DSXX:1:2268:20853:4601 chr2 33776018 N chr2 33776138 N DEL 5
A00404:156:HV37TDSXX:2:2513:7374:12007 chr2 33776018 N chr2 33776138 N DEL 5
A00297:158:HT275DSXX:3:1517:23050:23500 chr2 33776018 N chr2 33776138 N DEL 5
A00404:155:HV27LDSXX:4:2509:25536:35227 chr2 33776018 N chr2 33776138 N DEL 5
A00404:155:HV27LDSXX:1:2176:25093:21652 chr2 33776018 N chr2 33776138 N DEL 5
A00297:158:HT275DSXX:2:1206:24316:29199 chr2 33776018 N chr2 33776138 N DEL 5
A00297:158:HT275DSXX:2:1206:24704:29309 chr2 33776018 N chr2 33776138 N DEL 5
A00404:155:HV27LDSXX:3:2518:15817:16736 chr2 33776018 N chr2 33776138 N DEL 5
A00404:155:HV27LDSXX:3:2537:10474:31093 chr2 33776018 N chr2 33776138 N DEL 5
A00404:156:HV37TDSXX:1:1655:11324:32534 chr2 33776018 N chr2 33776138 N DEL 5
A00297:158:HT275DSXX:3:1521:24234:16313 chr2 33776018 N chr2 33776138 N DEL 5
A00404:155:HV27LDSXX:1:1621:4164:27899 chr2 33776018 N chr2 33776138 N DEL 5
A00404:156:HV37TDSXX:4:1329:14000:10394 chr2 33776018 N chr2 33776138 N DEL 5
A00404:156:HV37TDSXX:1:2221:1615:22232 chr2 33776018 N chr2 33776138 N DEL 5
A00297:158:HT275DSXX:4:2114:26811:30921 chr14 73451305 N chr14 73451583 N DUP 3
A00404:156:HV37TDSXX:4:1421:13738:2957 chr21 14671689 N chr21 14671758 N DEL 5
A00404:155:HV27LDSXX:4:2144:27118:25191 chr21 14671690 N chr21 14671759 N DEL 5
A00404:155:HV27LDSXX:4:2144:27389:24627 chr21 14671690 N chr21 14671759 N DEL 5
A00297:158:HT275DSXX:4:1310:5077:10723 chr12 120192805 N chr12 120193110 N DEL 2
A00297:158:HT275DSXX:1:2267:9697:10238 chr12 120192603 N chr12 120193227 N DUP 5
A00404:156:HV37TDSXX:2:1123:25599:19272 chr12 120192603 N chr12 120193227 N DUP 5
A00297:158:HT275DSXX:3:2608:24740:23547 chr12 120192603 N chr12 120193227 N DUP 5
A00404:155:HV27LDSXX:1:1139:8305:28181 chr12 120192603 N chr12 120193227 N DUP 5
A00404:155:HV27LDSXX:1:1139:8323:28181 chr12 120192603 N chr12 120193227 N DUP 5
A00404:156:HV37TDSXX:1:1265:14009:18959 chr12 120192603 N chr12 120193227 N DUP 5
A00297:158:HT275DSXX:1:2406:21603:35117 chr12 120192619 N chr12 120193245 N DEL 1
A00404:155:HV27LDSXX:1:1138:30192:22279 chr1 25768413 N chr1 25768470 N DEL 16
A00404:155:HV27LDSXX:1:1138:31150:25222 chr1 25768413 N chr1 25768470 N DEL 16
A00297:158:HT275DSXX:4:2236:10050:26788 chr1 25768266 N chr1 25768431 N DEL 1
A00297:158:HT275DSXX:3:1430:9381:20212 chr1 25768242 N chr1 25768653 N DUP 5
A00297:158:HT275DSXX:4:2135:6280:10739 chr20 57896044 N chr20 57896142 N DUP 5
A00297:158:HT275DSXX:4:2135:7229:9408 chr20 57896044 N chr20 57896142 N DUP 5
A00297:158:HT275DSXX:4:2135:8567:9846 chr20 57896044 N chr20 57896142 N DUP 5
A00404:156:HV37TDSXX:3:1511:8820:11287 chr20 57896044 N chr20 57896142 N DUP 5
A00404:155:HV27LDSXX:3:1450:25364:6997 chr17 40329718 N chr17 40329853 N DEL 5
A00404:156:HV37TDSXX:1:1415:8938:3004 chr14 95066593 N chr14 95066681 N DEL 5
A00404:155:HV27LDSXX:1:1274:32253:26819 chr14 95066626 N chr14 95066813 N DEL 13
A00404:156:HV37TDSXX:2:1614:1877:31955 chr14 95066627 N chr14 95066814 N DEL 12
A00297:158:HT275DSXX:3:1154:23538:17394 chr21 44365115 N chr21 44365188 N DEL 5
A00404:155:HV27LDSXX:1:2256:15854:8970 chr5 196700 N chr5 196784 N DUP 9
A00404:155:HV27LDSXX:2:2140:3775:17237 chr5 196786 N chr5 196871 N DEL 47
A00404:155:HV27LDSXX:2:2377:27570:21715 chr5 196609 N chr5 196834 N DEL 10
A00404:156:HV37TDSXX:4:1677:11487:10708 chr5 196790 N chr5 196875 N DEL 11
A00404:156:HV37TDSXX:1:1538:5801:1266 chr20 61686740 N chr20 61686801 N DEL 9
A00404:156:HV37TDSXX:1:2349:4137:3427 chr19 2540015 N chr19 2540206 N DUP 2
A00297:158:HT275DSXX:1:1631:26928:17096 chr2 29217079 N chr2 29217184 N DEL 12
A00297:158:HT275DSXX:1:1343:17517:24909 chr2 29217079 N chr2 29217184 N DEL 14
A00297:158:HT275DSXX:1:2140:5909:18176 chr2 29217113 N chr2 29217198 N DUP 7
A00404:156:HV37TDSXX:4:2136:9805:16438 chr2 29217116 N chr2 29217201 N DUP 4
A00404:156:HV37TDSXX:4:1126:17743:28870 chr2 29217118 N chr2 29217203 N DUP 2
A00404:156:HV37TDSXX:3:2673:5909:9533 chr2 29217217 N chr2 29217289 N DUP 10
A00297:158:HT275DSXX:4:2511:27697:11788 chr5 15556137 N chr5 15556244 N DEL 5
A00404:156:HV37TDSXX:2:1652:6804:20322 chr5 15556137 N chr5 15556244 N DEL 5
A00404:155:HV27LDSXX:2:1305:4707:1188 chrX 29333333 N chrX 29333589 N DEL 4
A00404:155:HV27LDSXX:4:2635:13675:27461 chrX 29333383 N chrX 29333639 N DEL 5
A00404:156:HV37TDSXX:4:2254:5647:20447 chrX 29333403 N chrX 29334101 N DEL 5
A00297:158:HT275DSXX:1:1475:17472:25989 chrX 29333431 N chrX 29333735 N DEL 25
A00404:156:HV37TDSXX:1:1358:5584:28948 chrX 29333353 N chrX 29333482 N DEL 1
A00297:158:HT275DSXX:2:1627:19443:18317 chrX 29333536 N chrX 29334457 N DEL 10
A00404:156:HV37TDSXX:4:2250:25907:15264 chrX 29333561 N chrX 29334229 N DEL 1
A00404:155:HV27LDSXX:2:2622:14769:36558 chrX 29333468 N chrX 29333594 N DUP 8
A00297:158:HT275DSXX:2:1209:29423:6825 chrX 29333561 N chrX 29334229 N DEL 1
A00404:155:HV27LDSXX:2:2624:6931:26209 chrX 29333543 N chrX 29333943 N DUP 9
A00404:155:HV27LDSXX:4:1459:5683:8046 chrX 29333572 N chrX 29333966 N DEL 5
A00297:158:HT275DSXX:2:1624:19587:36292 chrX 29333572 N chrX 29333964 N DUP 4
A00404:156:HV37TDSXX:2:1413:17390:1329 chrX 29333576 N chrX 29333704 N DEL 5
A00404:156:HV37TDSXX:2:1354:17400:12148 chrX 29333659 N chrX 29333836 N DEL 7
A00404:156:HV37TDSXX:2:2311:15203:17519 chrX 29333839 N chrX 29334106 N DEL 2
A00404:156:HV37TDSXX:4:1150:10239:19852 chrX 29333839 N chrX 29334106 N DEL 1
A00404:156:HV37TDSXX:1:2247:1208:24533 chrX 29333470 N chrX 29333774 N DEL 7
A00297:158:HT275DSXX:2:2455:5900:11397 chrX 29333686 N chrX 29333863 N DEL 15
A00297:158:HT275DSXX:3:2618:27082:37027 chrX 29333438 N chrX 29333870 N DEL 5
A00404:156:HV37TDSXX:4:1275:7003:4194 chrX 29333594 N chrX 29333948 N DEL 7
A00404:155:HV27LDSXX:4:1304:19361:24846 chrX 29333570 N chrX 29333923 N DEL 3
A00297:158:HT275DSXX:4:2167:13991:12164 chrX 29333980 N chrX 29334508 N DEL 5
A00404:156:HV37TDSXX:2:2312:9552:6637 chrX 29333980 N chrX 29334508 N DEL 3
A00404:155:HV27LDSXX:1:1202:2058:6965 chrX 29333695 N chrX 29333872 N DEL 18
A00404:156:HV37TDSXX:1:2559:10547:33098 chrX 29333836 N chrX 29334101 N DUP 5
A00404:156:HV37TDSXX:2:1118:20076:3349 chrX 29333722 N chrX 29334114 N DUP 1
A00404:156:HV37TDSXX:4:2541:18683:31814 chrX 29334010 N chrX 29334282 N DUP 4
A00297:158:HT275DSXX:2:2455:5900:11397 chrX 29333686 N chrX 29333863 N DEL 10
A00297:158:HT275DSXX:3:1321:29532:17002 chrX 29333722 N chrX 29334114 N DUP 5
A00297:158:HT275DSXX:1:1162:14398:20979 chrX 29333722 N chrX 29334114 N DUP 5
A00404:155:HV27LDSXX:4:1626:21504:36949 chrX 29333545 N chrX 29334113 N DUP 1
A00404:156:HV37TDSXX:4:2541:18683:31814 chrX 29333697 N chrX 29334042 N DEL 10
A00297:158:HT275DSXX:4:1651:7636:14372 chrX 29333836 N chrX 29334150 N DUP 10
A00404:155:HV27LDSXX:4:1463:21450:7858 chrX 29334066 N chrX 29334163 N DUP 2
A00404:156:HV37TDSXX:2:2519:20980:34695 chrX 29334066 N chrX 29334163 N DUP 1
A00297:158:HT275DSXX:2:1214:10031:10661 chrX 29334074 N chrX 29334171 N DUP 5
A00297:158:HT275DSXX:3:2556:31439:5525 chrX 29334066 N chrX 29334163 N DUP 5
A00404:156:HV37TDSXX:2:1164:5864:3693 chrX 29333594 N chrX 29334066 N DEL 10
A00404:155:HV27LDSXX:4:2231:15835:12633 chrX 29333438 N chrX 29334136 N DEL 5
A00297:158:HT275DSXX:2:2475:15863:10739 chrX 29333594 N chrX 29334066 N DEL 2
A00297:158:HT275DSXX:3:2663:9525:3521 chrX 29333672 N chrX 29334164 N DEL 5
A00404:155:HV27LDSXX:2:2454:2193:28181 chrX 29333672 N chrX 29334164 N DEL 5
A00297:158:HT275DSXX:2:2143:9733:23954 chrX 29334130 N chrX 29334229 N DEL 5
A00404:156:HV37TDSXX:1:1271:9887:6997 chrX 29333574 N chrX 29334242 N DEL 2
A00404:155:HV27LDSXX:4:2559:16468:26725 chrX 29333541 N chrX 29334337 N DUP 18
A00297:158:HT275DSXX:3:2627:11107:24330 chrX 29333868 N chrX 29334485 N DEL 12
A00404:155:HV27LDSXX:2:2529:5466:2973 chrX 29333862 N chrX 29334479 N DEL 7
A00404:155:HV27LDSXX:2:1575:22227:11866 chrX 29333862 N chrX 29334479 N DEL 7
A00297:158:HT275DSXX:2:1473:27353:35806 chrX 29333862 N chrX 29334479 N DEL 7
A00404:156:HV37TDSXX:4:1315:31367:15452 chrX 29333410 N chrX 29334584 N DUP 1
A00404:156:HV37TDSXX:3:2651:18611:32534 chrX 29334497 N chrX 29334624 N DUP 12
A00404:155:HV27LDSXX:4:2108:1425:1799 chrX 29333910 N chrX 29334604 N DUP 6
A00404:156:HV37TDSXX:3:1615:30129:5165 chrX 29334242 N chrX 29334496 N DEL 1
A00404:155:HV27LDSXX:4:2475:22679:32377 chrX 29333460 N chrX 29334508 N DEL 10
A00297:158:HT275DSXX:1:1520:26006:4633 chrX 29333598 N chrX 29334519 N DEL 4
A00404:156:HV37TDSXX:4:2141:29568:7263 chrX 29333522 N chrX 29334570 N DEL 5
A00404:156:HV37TDSXX:1:1322:17454:30311 chrX 29333583 N chrX 29334582 N DEL 2
A00297:158:HT275DSXX:3:1641:29740:20932 chrX 29334129 N chrX 29334606 N DEL 9
A00404:155:HV27LDSXX:3:1266:21992:16814 chrX 29334128 N chrX 29334606 N DEL 7
A00404:155:HV27LDSXX:1:1402:26811:1110 chr20 49214098 N chr20 49214405 N DEL 4
A00404:156:HV37TDSXX:2:1420:31313:10911 chr20 49214128 N chr20 49214433 N DUP 5
A00404:156:HV37TDSXX:2:1374:30291:21167 chr20 49214128 N chr20 49214433 N DUP 5
A00297:158:HT275DSXX:1:2264:29179:2206 chr6 89339622 N chr6 89339796 N DEL 6
A00404:156:HV37TDSXX:3:2663:20302:2456 chr6 89339622 N chr6 89339796 N DEL 5
A00404:156:HV37TDSXX:3:1371:1597:34100 chr8 17882905 N chr8 17882972 N DEL 12
A00404:156:HV37TDSXX:4:1261:13720:30577 chr8 17883221 N chr8 17883285 N DEL 13
A00404:156:HV37TDSXX:2:1376:13250:28354 chr8 17883362 N chr8 17883433 N DEL 5
A00404:156:HV37TDSXX:2:1376:13250:28385 chr8 17883362 N chr8 17883433 N DEL 5
A00297:158:HT275DSXX:1:2230:8775:12900 chr8 17883031 N chr8 17883433 N DEL 5
A00404:156:HV37TDSXX:1:2614:21206:21684 chr8 17882996 N chr8 17883433 N DEL 5
A00404:156:HV37TDSXX:1:2511:15528:1235 chr5 135806758 N chr5 135807189 N DUP 5
A00297:158:HT275DSXX:2:2521:9742:20275 chr10 132149704 N chr10 132149787 N DUP 7
A00404:156:HV37TDSXX:4:1555:29957:26569 chr17 72783215 N chr17 72783279 N DEL 8
A00404:156:HV37TDSXX:1:2115:21676:7968 chr7 121409214 N chr7 121409266 N DUP 2
A00404:155:HV27LDSXX:4:1421:25898:15060 chr7 121409215 N chr7 121409267 N DUP 1
A00297:158:HT275DSXX:3:2135:19723:8656 chr1 55983647 N chr1 55983708 N DEL 5
A00404:156:HV37TDSXX:2:1154:30246:16454 chr4 186239011 N chr4 186239083 N DEL 2
A00297:158:HT275DSXX:2:2620:8377:22576 chr4 186239011 N chr4 186239083 N DEL 5
A00297:158:HT275DSXX:3:1257:16884:20525 chr4 186239011 N chr4 186239083 N DEL 5
A00297:158:HT275DSXX:1:1405:32570:4225 chr4 186239011 N chr4 186239083 N DEL 5
A00297:158:HT275DSXX:3:1124:13955:6308 chr4 186239011 N chr4 186239083 N DEL 5
A00404:155:HV27LDSXX:3:1338:18258:28479 chr4 186239011 N chr4 186239083 N DEL 5
A00404:155:HV27LDSXX:4:2306:16215:6464 chr4 186239011 N chr4 186239083 N DEL 5
A00297:158:HT275DSXX:4:1424:7699:14231 chr4 186239011 N chr4 186239083 N DEL 5
A00404:155:HV27LDSXX:4:1616:16089:28166 chr4 186239011 N chr4 186239083 N DEL 5
A00404:156:HV37TDSXX:4:2344:5511:13792 chr4 186239011 N chr4 186239083 N DEL 5
A00404:156:HV37TDSXX:2:1546:24080:2957 chr4 186239011 N chr4 186239083 N DEL 12
A00404:155:HV27LDSXX:2:1121:22978:18020 chr4 186239011 N chr4 186239083 N DEL 15
A00404:155:HV27LDSXX:1:1107:30129:8108 chr19 15887360 N chr19 15887537 N DUP 1
A00404:156:HV37TDSXX:3:2568:16848:26694 chr19 15887522 N chr19 15887585 N DUP 5
A00404:155:HV27LDSXX:3:2318:2618:10222 chr19 15887444 N chr19 15887685 N DUP 5
A00297:158:HT275DSXX:4:1619:25970:19570 chr19 15887531 N chr19 15887772 N DUP 9
A00404:156:HV37TDSXX:2:2245:30174:32487 chr12 8926492 N chr12 8926786 N DEL 19
A00297:158:HT275DSXX:2:1273:30671:31751 chr12 8926701 N chr12 8926996 N DEL 4
A00297:158:HT275DSXX:3:2443:4047:17926 chr17 21236032 N chr17 21236121 N DUP 1
A00404:155:HV27LDSXX:1:2654:23113:36417 chr17 21236128 N chr17 21236433 N DEL 2
A00404:156:HV37TDSXX:4:1462:15619:20149 chr20 62922261 N chr20 62922390 N DUP 5
A00404:156:HV37TDSXX:2:1106:24379:26209 chr20 62922261 N chr20 62922390 N DUP 5
A00297:158:HT275DSXX:3:1639:23873:31939 chr20 62922277 N chr20 62922406 N DEL 7
A00297:158:HT275DSXX:4:1101:32687:29418 chr15 93125811 N chr15 93125957 N DEL 7
A00404:155:HV27LDSXX:3:1528:25165:14199 chr15 93125815 N chr15 93125961 N DEL 7
A00297:158:HT275DSXX:3:2112:9914:10614 chr15 93125817 N chr15 93125963 N DEL 7
A00404:156:HV37TDSXX:4:2354:25364:6370 chr15 93125818 N chr15 93125964 N DEL 7
A00297:158:HT275DSXX:2:1613:23131:16752 chr15 93125823 N chr15 93125969 N DEL 2
A00297:158:HT275DSXX:4:1628:24786:23750 chr15 93125823 N chr15 93125969 N DEL 2
A00404:156:HV37TDSXX:2:2116:3052:24471 chr15 93125816 N chr15 93125963 N DEL 8
A00404:155:HV27LDSXX:1:2276:6668:8625 chr6 43798046 N chr6 43798123 N DEL 12
A00404:155:HV27LDSXX:2:1146:2862:5760 chr6 43798059 N chr6 43798137 N DEL 10
A00404:156:HV37TDSXX:3:1520:16703:4366 chr6 43798059 N chr6 43798137 N DEL 5
A00404:156:HV37TDSXX:4:1612:30454:28620 chr6 43798084 N chr6 43798237 N DUP 20
A00297:158:HT275DSXX:2:2555:23484:3646 chr6 43798120 N chr6 43798273 N DUP 6
A00404:155:HV27LDSXX:2:1111:29098:26647 chr6 43798183 N chr6 43798259 N DUP 40
A00297:158:HT275DSXX:1:1156:10827:35931 chr6 43798192 N chr6 43798268 N DUP 40
A00404:156:HV37TDSXX:3:2667:31656:14325 chr6 43798183 N chr6 43798259 N DUP 35
A00404:156:HV37TDSXX:1:1541:7229:18615 chr6 43798197 N chr6 43798273 N DUP 15
A00297:158:HT275DSXX:1:1456:25970:18944 chr6 43798183 N chr6 43798259 N DUP 35
A00297:158:HT275DSXX:1:2507:26142:31767 chr6 43798192 N chr6 43798268 N DUP 45
A00404:156:HV37TDSXX:3:1116:9353:28244 chr6 43798115 N chr6 43798268 N DUP 4
A00297:158:HT275DSXX:2:2160:21621:36808 chr6 43798115 N chr6 43798268 N DUP 7
A00404:155:HV27LDSXX:2:1146:2862:5760 chr6 43798192 N chr6 43798268 N DUP 10
A00404:155:HV27LDSXX:2:2146:3784:5102 chr6 43798192 N chr6 43798268 N DUP 10
A00404:156:HV37TDSXX:2:1638:14904:23641 chr6 43798192 N chr6 43798268 N DUP 11
A00297:158:HT275DSXX:3:1350:29297:17221 chr6 43798192 N chr6 43798268 N DUP 22
A00404:156:HV37TDSXX:2:2652:10547:5666 chr6 43798192 N chr6 43798268 N DUP 25
A00297:158:HT275DSXX:1:1543:25635:29669 chr6 43798192 N chr6 43798268 N DUP 26
A00404:155:HV27LDSXX:3:1418:8486:6856 chr6 43798183 N chr6 43798259 N DUP 39
A00297:158:HT275DSXX:2:1213:30563:29904 chr6 43798192 N chr6 43798268 N DUP 35
A00404:156:HV37TDSXX:2:1223:10890:30248 chr6 43798192 N chr6 43798268 N DUP 35
A00297:158:HT275DSXX:1:2232:12255:33144 chr6 43798197 N chr6 43798273 N DUP 5
A00297:158:HT275DSXX:2:2505:28917:4445 chr6 43798197 N chr6 43798273 N DUP 6
A00404:155:HV27LDSXX:2:2635:6316:26772 chr6 43798183 N chr6 43798259 N DUP 31
A00297:158:HT275DSXX:3:2667:24840:12978 chr6 43798192 N chr6 43798268 N DUP 42
A00297:158:HT275DSXX:2:1557:9959:2268 chr6 43798192 N chr6 43798268 N DUP 42
A00404:156:HV37TDSXX:4:2333:17761:2597 chr6 43798192 N chr6 43798268 N DUP 37
A00404:155:HV27LDSXX:4:2555:16523:28792 chr6 43798192 N chr6 43798268 N DUP 37
A00404:156:HV37TDSXX:2:1223:10890:30248 chr6 43798119 N chr6 43798348 N DUP 3
A00404:156:HV37TDSXX:1:2130:22625:32597 chr6 43798253 N chr6 43798330 N DEL 37
A00404:156:HV37TDSXX:4:2666:13693:13056 chr6 43798238 N chr6 43798315 N DEL 37
A00404:155:HV27LDSXX:2:2571:19135:16000 chr6 43798089 N chr6 43798434 N DEL 5
A00404:156:HV37TDSXX:2:1659:12093:9064 chr6 154397868 N chr6 154397990 N DEL 2
A00404:156:HV37TDSXX:1:2119:10456:35258 chr8 51231316 N chr8 51231434 N DUP 5
A00404:156:HV37TDSXX:4:2461:13494:24236 chr5 14793141 N chr5 14793190 N DUP 9
A00297:158:HT275DSXX:3:1416:23502:29230 chr5 14793141 N chr5 14793190 N DUP 10
A00297:158:HT275DSXX:3:1416:24361:30373 chr5 14793141 N chr5 14793190 N DUP 6
A00297:158:HT275DSXX:3:1316:16351:3129 chr5 14793165 N chr5 14793218 N DEL 13
A00297:158:HT275DSXX:1:1565:3269:7654 chr4 49152705 N chr4 49152838 N DUP 4
A00404:155:HV27LDSXX:3:2571:9399:25285 chr4 49152767 N chr4 49152919 N DUP 3
A00404:156:HV37TDSXX:2:1207:26115:1532 chr4 49152689 N chr4 49152871 N DUP 10
A00297:158:HT275DSXX:2:2504:14995:15530 chr7 88266696 N chr7 88266793 N DUP 10
A00404:156:HV37TDSXX:4:2441:20934:8563 chr7 88266935 N chr7 88267016 N DEL 5
A00404:155:HV27LDSXX:3:1230:4896:30264 chr7 88266943 N chr7 88267024 N DEL 5
A00404:155:HV27LDSXX:2:1274:27434:2848 chr6 69467828 N chr6 69468105 N DUP 5
A00404:155:HV27LDSXX:4:1267:5095:3521 chr7 71798220 N chr7 71798285 N DEL 5
A00404:155:HV27LDSXX:3:1638:27552:12665 chr10 10033523 N chr10 10033624 N DUP 2
A00404:155:HV27LDSXX:3:1638:27670:12868 chr10 10033523 N chr10 10033624 N DUP 2
A00404:156:HV37TDSXX:2:1638:14226:25316 chr10 10033523 N chr10 10033624 N DUP 2
A00297:158:HT275DSXX:3:2202:21187:7874 chr10 10033523 N chr10 10033624 N DUP 3
A00297:158:HT275DSXX:4:2663:23384:18035 chr10 10033543 N chr10 10033644 N DUP 13
A00297:158:HT275DSXX:1:2238:19081:21793 chr10 10033593 N chr10 10033644 N DUP 22
A00404:155:HV27LDSXX:1:2516:12988:35258 chr10 10033593 N chr10 10033644 N DUP 25
A00404:156:HV37TDSXX:2:2569:24361:34945 chr10 10033551 N chr10 10033602 N DUP 14
A00404:156:HV37TDSXX:2:2569:24514:35618 chr10 10033593 N chr10 10033644 N DUP 19
A00404:156:HV37TDSXX:2:2378:17273:1188 chr10 10033593 N chr10 10033644 N DUP 19
A00404:155:HV27LDSXX:3:2425:20835:23390 chr10 10033593 N chr10 10033644 N DUP 14
A00404:156:HV37TDSXX:4:2275:22281:31563 chr10 10033593 N chr10 10033644 N DUP 14
A00404:155:HV27LDSXX:2:1219:14651:1438 chr10 10033593 N chr10 10033644 N DUP 14
A00404:155:HV27LDSXX:2:1404:31304:6136 chr10 10033546 N chr10 10033625 N DEL 10
A00297:158:HT275DSXX:1:2177:4408:29512 chr10 10033583 N chr10 10033636 N DEL 4
A00404:155:HV27LDSXX:2:2263:27959:30780 chr22 50686542 N chr22 50686689 N DUP 5
A00404:156:HV37TDSXX:3:1457:22453:29168 chr22 50686587 N chr22 50686854 N DEL 5
A00404:156:HV37TDSXX:3:2457:23972:35900 chr22 50686676 N chr22 50686943 N DEL 5
A00404:156:HV37TDSXX:3:2457:23972:35900 chr22 50686676 N chr22 50686943 N DEL 5
A00404:156:HV37TDSXX:3:2213:26332:21042 chr22 50686625 N chr22 50686949 N DUP 5
A00404:155:HV27LDSXX:3:2315:24849:17973 chr22 50686677 N chr22 50686942 N DUP 5
A00404:155:HV27LDSXX:1:2218:32298:16438 chr6 167514431 N chr6 167514591 N DUP 5
A00404:156:HV37TDSXX:2:1619:16568:23234 chr6 167514492 N chr6 167514594 N DUP 5
A00404:156:HV37TDSXX:4:1126:4797:14747 chr6 167514539 N chr6 167514643 N DEL 5
A00297:158:HT275DSXX:1:1427:26096:3192 chr6 167514539 N chr6 167514643 N DEL 5
A00297:158:HT275DSXX:1:1122:17237:35728 chr6 167514539 N chr6 167514643 N DEL 5
A00297:158:HT275DSXX:4:2653:5846:30154 chr6 167514539 N chr6 167514643 N DEL 5
A00297:158:HT275DSXX:1:2665:1895:20400 chr6 167514541 N chr6 167514645 N DEL 5
A00404:156:HV37TDSXX:3:2123:10285:16454 chr6 167514541 N chr6 167514645 N DEL 5
A00297:158:HT275DSXX:1:1633:6460:11616 chr4 89802770 N chr4 89802907 N DEL 7
A00404:155:HV27LDSXX:4:2112:4417:34131 chr3 175119938 N chr3 175120026 N DEL 9
A00404:155:HV27LDSXX:3:1673:22372:31000 chr14 54203722 N chr14 54204076 N DEL 11
A00404:155:HV27LDSXX:2:2165:15076:24909 chr14 54203801 N chr14 54203977 N DEL 5
A00404:156:HV37TDSXX:1:1372:14290:16407 chr14 54203801 N chr14 54203977 N DEL 5
A00297:158:HT275DSXX:3:1353:1570:1360 chr14 54203801 N chr14 54203977 N DEL 5
A00404:155:HV27LDSXX:2:1157:14525:2472 chr14 54203801 N chr14 54203977 N DEL 6
A00404:155:HV27LDSXX:1:1554:2844:26522 chr14 54203840 N chr14 54204014 N DUP 11
A00404:155:HV27LDSXX:3:1403:6985:32252 chr14 54203755 N chr14 54204057 N DUP 5
A00404:155:HV27LDSXX:4:2415:7771:17957 chr14 54203803 N chr14 54203928 N DUP 18
A00404:155:HV27LDSXX:3:1642:29758:16736 chr14 54203839 N chr14 54204241 N DEL 12
A00404:156:HV37TDSXX:1:2470:16333:3912 chr14 54203767 N chr14 54204119 N DUP 5
A00404:156:HV37TDSXX:4:2205:3423:15374 chr14 54203766 N chr14 54203892 N DUP 8
A00404:155:HV27LDSXX:3:1642:29758:16736 chr14 54203839 N chr14 54204241 N DEL 12
A00404:155:HV27LDSXX:4:2336:2564:1016 chr14 54203898 N chr14 54204076 N DEL 5
A00297:158:HT275DSXX:3:1353:1570:1360 chr14 54203803 N chr14 54203928 N DUP 6
A00404:155:HV27LDSXX:3:1403:6985:32252 chr14 54203840 N chr14 54204014 N DUP 7
A00297:158:HT275DSXX:3:1362:28149:21809 chr14 54203947 N chr14 54204076 N DEL 1
A00404:155:HV27LDSXX:2:2378:25292:16705 chr14 54203752 N chr14 54203929 N DEL 14
A00297:158:HT275DSXX:4:2644:28348:36276 chr14 54203686 N chr14 54203959 N DEL 9
A00404:155:HV27LDSXX:2:2378:25292:16705 chr14 54203989 N chr14 54204216 N DEL 5
A00404:155:HV27LDSXX:2:1141:19190:35102 chr14 54203598 N chr14 54204047 N DUP 7
A00404:156:HV37TDSXX:4:2662:19560:17550 chr14 54203995 N chr14 54204220 N DUP 3
A00404:155:HV27LDSXX:3:2372:21612:33191 chr14 54203868 N chr14 54204093 N DUP 15
A00404:155:HV27LDSXX:2:2437:18728:35556 chr14 54203537 N chr14 54204212 N DUP 3
A00404:156:HV37TDSXX:3:1469:7491:6073 chr14 54203680 N chr14 54204132 N DEL 5
A00297:158:HT275DSXX:3:2136:30364:23140 chr14 54204238 N chr14 54204493 N DEL 1
A00404:156:HV37TDSXX:2:2531:25482:31031 chr14 54204238 N chr14 54204493 N DEL 3
A00404:156:HV37TDSXX:3:2406:27706:31250 chr14 54203648 N chr14 54204198 N DEL 5
A00404:155:HV27LDSXX:3:2224:17951:29763 chr14 54204274 N chr14 54204402 N DEL 5
A00404:155:HV27LDSXX:3:2120:23583:35164 chr14 54204326 N chr14 54204405 N DEL 8
A00297:158:HT275DSXX:4:2115:5999:30044 chr14 54204196 N chr14 54204322 N DUP 5
A00297:158:HT275DSXX:4:2102:17264:15577 chr14 54203762 N chr14 54203888 N DUP 28
A00404:155:HV27LDSXX:1:2542:32588:9204 chr14 54204191 N chr14 54204446 N DEL 15
A00404:155:HV27LDSXX:1:2542:32588:9204 chr14 54204191 N chr14 54204446 N DEL 10
A00404:156:HV37TDSXX:2:2531:25482:31031 chr14 54203837 N chr14 54204493 N DEL 5
A00404:156:HV37TDSXX:2:2531:25979:31328 chr14 54204365 N chr14 54204493 N DEL 10
A00404:156:HV37TDSXX:3:1565:14823:25128 chr11 69733868 N chr11 69733936 N DEL 5
A00297:158:HT275DSXX:3:1319:10972:30796 chr11 69733868 N chr11 69733936 N DEL 13
A00297:158:HT275DSXX:4:2456:32154:12712 chr11 69733884 N chr11 69733952 N DEL 8
A00404:155:HV27LDSXX:2:2574:6849:31485 chr11 69733829 N chr11 69733962 N DEL 3
A00404:156:HV37TDSXX:2:2627:3405:2628 chrX 2253512 N chrX 2253613 N DEL 5
A00404:155:HV27LDSXX:4:2416:19144:28134 chrX 2253423 N chrX 2253474 N DEL 31
A00404:155:HV27LDSXX:4:1430:14009:19398 chrX 2253500 N chrX 2253549 N DUP 5
A00404:156:HV37TDSXX:4:2634:22372:35102 chrX 2253425 N chrX 2253476 N DEL 20
A00297:158:HT275DSXX:1:1173:10185:22639 chrX 2253474 N chrX 2253573 N DUP 14
A00297:158:HT275DSXX:3:1163:5909:16235 chrX 2253474 N chrX 2253573 N DUP 13
A00297:158:HT275DSXX:1:2645:30382:28557 chrX 2253476 N chrX 2253525 N DUP 7
A00297:158:HT275DSXX:4:2430:13440:8703 chrX 2253474 N chrX 2253573 N DUP 11
A00297:158:HT275DSXX:1:2418:5276:31798 chrX 2253477 N chrX 2253576 N DUP 12
A00404:155:HV27LDSXX:3:2261:10122:12696 chrX 2253340 N chrX 2253488 N DEL 1
A00404:155:HV27LDSXX:3:1616:5285:33442 chrX 2253477 N chrX 2253576 N DUP 20
A00404:155:HV27LDSXX:1:2609:19090:22467 chrX 2253497 N chrX 2253596 N DUP 10
A00297:158:HT275DSXX:2:1524:23601:2440 chrX 2253477 N chrX 2253576 N DUP 22
A00297:158:HT275DSXX:4:1422:28637:22341 chrX 2253523 N chrX 2253622 N DUP 10
A00404:155:HV27LDSXX:4:1417:25301:10739 chrX 2253377 N chrX 2253528 N DEL 5
A00404:156:HV37TDSXX:2:2660:5656:2331 chrX 2253450 N chrX 2253551 N DEL 5
A00297:158:HT275DSXX:3:1524:10999:24330 chrX 2253496 N chrX 2253597 N DEL 5
A00297:158:HT275DSXX:3:2371:22263:12900 chrX 2253512 N chrX 2253613 N DEL 5
A00297:158:HT275DSXX:4:1214:2230:29183 chr18 51050517 N chr18 51050821 N DUP 3
A00404:155:HV27LDSXX:1:2162:3486:26882 chr1 197770780 N chr1 197770933 N DEL 3
A00297:158:HT275DSXX:1:1504:18240:33238 chr14 38837537 N chr14 38837678 N DEL 13
A00297:158:HT275DSXX:4:1261:29306:3239 chr7 157461427 N chr7 157461606 N DEL 20
A00404:155:HV27LDSXX:1:1510:9399:12633 chr7 157461482 N chr7 157461609 N DEL 1
A00297:158:HT275DSXX:2:1171:23583:4601 chr7 157461484 N chr7 157461629 N DEL 4
A00404:156:HV37TDSXX:4:1610:21956:5134 chr7 157461484 N chr7 157461629 N DEL 5
A00297:158:HT275DSXX:2:1613:32606:10989 chr7 157461489 N chr7 157461620 N DEL 14
A00297:158:HT275DSXX:3:2361:12020:32769 chr7 157461491 N chr7 157461594 N DEL 17
A00297:158:HT275DSXX:4:2114:10402:34413 chr7 157461412 N chr7 157461701 N DUP 32
A00404:155:HV27LDSXX:3:1577:16143:20807 chr7 157461448 N chr7 157461583 N DUP 16
A00297:158:HT275DSXX:2:2317:15619:20964 chr7 157461420 N chr7 157461479 N DUP 10
A00404:155:HV27LDSXX:4:2157:25156:11553 chr7 157461416 N chr7 157461637 N DUP 11
A00404:155:HV27LDSXX:1:1512:6343:24878 chr7 157461539 N chr7 157461626 N DEL 13
A00404:155:HV27LDSXX:1:1512:6533:27085 chr7 157461539 N chr7 157461626 N DEL 13
A00404:156:HV37TDSXX:2:1348:15474:25128 chr7 157461525 N chr7 157461638 N DEL 20
A00404:155:HV27LDSXX:2:2316:22110:20744 chr7 157461525 N chr7 157461638 N DEL 23
A00297:158:HT275DSXX:4:2374:19569:21543 chr7 157461495 N chr7 157461718 N DUP 13
A00404:156:HV37TDSXX:1:1404:9353:36072 chr7 157461437 N chr7 157461540 N DUP 9
A00297:158:HT275DSXX:2:2644:22815:8531 chr7 157461441 N chr7 157461726 N DUP 4
A00404:155:HV27LDSXX:3:1633:23502:28980 chr7 157461525 N chr7 157461638 N DEL 25
A00297:158:HT275DSXX:4:1222:21088:2660 chr7 157461525 N chr7 157461576 N DEL 22
A00404:156:HV37TDSXX:1:1446:16785:18349 chr7 157461531 N chr7 157461626 N DEL 18
A00297:158:HT275DSXX:3:1426:9896:28463 chr7 157461541 N chr7 157461620 N DEL 15
A00297:158:HT275DSXX:4:1222:21088:2660 chr7 157461560 N chr7 157461821 N DUP 19
A00404:156:HV37TDSXX:2:1302:30924:15280 chr7 157461440 N chr7 157461505 N DEL 8
A00404:156:HV37TDSXX:3:1537:32524:3239 chr7 157461530 N chr7 157461655 N DUP 15
A00404:155:HV27LDSXX:4:2253:20193:11694 chr7 157461608 N chr7 157461677 N DUP 20
A00297:158:HT275DSXX:4:1246:22498:6292 chr7 157461467 N chr7 157461532 N DEL 5
A00297:158:HT275DSXX:4:2246:18412:3161 chr7 157461467 N chr7 157461532 N DEL 5
A00404:156:HV37TDSXX:3:1465:30228:33019 chr7 157461564 N chr7 157461713 N DUP 9
A00404:156:HV37TDSXX:3:1318:18882:11835 chr7 157461510 N chr7 157461575 N DUP 17
A00404:156:HV37TDSXX:4:2618:7988:36245 chr7 157461552 N chr7 157461635 N DUP 17
A00404:155:HV27LDSXX:4:2104:27751:16924 chr7 157461608 N chr7 157461677 N DUP 23
A00297:158:HT275DSXX:1:2240:12120:8985 chr7 157461439 N chr7 157461554 N DEL 11
A00404:155:HV27LDSXX:4:1559:6777:23876 chr7 157461445 N chr7 157461552 N DEL 5
A00404:155:HV27LDSXX:3:1604:2537:12618 chr7 157461511 N chr7 157461586 N DEL 10
A00404:155:HV27LDSXX:1:2349:23285:11443 chr7 157461567 N chr7 157461754 N DEL 8
A00297:158:HT275DSXX:3:1548:27742:21355 chr7 157461642 N chr7 157461709 N DUP 20
A00404:156:HV37TDSXX:4:2220:16902:29450 chr7 157461433 N chr7 157461564 N DEL 3
A00297:158:HT275DSXX:3:1356:8223:24158 chr7 157461445 N chr7 157461650 N DUP 4
A00404:155:HV27LDSXX:1:1665:31250:21261 chr7 157461508 N chr7 157461711 N DUP 15
A00404:156:HV37TDSXX:3:1352:17996:20008 chr7 157461414 N chr7 157461673 N DUP 13
A00404:155:HV27LDSXX:2:1117:25780:36276 chr7 157461529 N chr7 157461624 N DEL 20
A00297:158:HT275DSXX:4:1562:25988:30592 chr7 157461489 N chr7 157461594 N DEL 16
A00404:155:HV27LDSXX:4:1140:24415:34945 chr7 157461606 N chr7 157461827 N DUP 18
A00404:155:HV27LDSXX:1:2613:24894:20149 chr7 157461575 N chr7 157461668 N DEL 19
A00297:158:HT275DSXX:2:2444:26594:29543 chr7 157461600 N chr7 157461653 N DUP 20
A00297:158:HT275DSXX:3:2330:3495:31344 chr7 157461482 N chr7 157461563 N DUP 14
A00404:155:HV27LDSXX:3:1170:24840:13542 chr7 157461531 N chr7 157461712 N DUP 12
A00297:158:HT275DSXX:2:1417:21621:32863 chr7 157461642 N chr7 157461721 N DUP 17
A00404:155:HV27LDSXX:3:1315:8504:15436 chr7 157461531 N chr7 157461712 N DUP 12
A00404:155:HV27LDSXX:3:2315:6289:35117 chr7 157461530 N chr7 157461589 N DUP 10
A00404:155:HV27LDSXX:3:2333:21215:2503 chr7 157461531 N chr7 157461712 N DUP 12
A00404:156:HV37TDSXX:3:1122:3441:18850 chr7 157461639 N chr7 157461702 N DUP 11
A00404:156:HV37TDSXX:2:2639:19153:6104 chr7 157461642 N chr7 157461721 N DUP 16
A00297:158:HT275DSXX:2:2668:18412:13495 chr7 157461530 N chr7 157461647 N DUP 18
A00297:158:HT275DSXX:2:2654:24334:17926 chr7 157461641 N chr7 157461708 N DUP 4
A00297:158:HT275DSXX:3:2361:12020:32769 chr7 157461607 N chr7 157461718 N DUP 16
A00404:155:HV27LDSXX:2:1119:10438:22232 chr7 157461466 N chr7 157461693 N DUP 1
A00404:155:HV27LDSXX:3:1567:8865:31219 chr7 157461608 N chr7 157461677 N DUP 21
A00297:158:HT275DSXX:4:2374:19569:21543 chr7 157461414 N chr7 157461703 N DUP 20
A00297:158:HT275DSXX:3:1678:19199:2957 chr7 157461594 N chr7 157461693 N DUP 13
A00404:155:HV27LDSXX:1:1407:8043:6402 chr7 157461642 N chr7 157461709 N DUP 21
A00404:155:HV27LDSXX:3:2465:23032:18270 chr7 157461614 N chr7 157461665 N DUP 6
A00404:156:HV37TDSXX:1:1132:27444:18677 chr7 157461531 N chr7 157461618 N DUP 9
A00404:155:HV27LDSXX:3:1573:23764:25457 chr7 157461531 N chr7 157461618 N DUP 16
A00404:155:HV27LDSXX:2:2577:30020:7795 chr7 157461525 N chr7 157461578 N DEL 17
A00297:158:HT275DSXX:2:1227:14561:26710 chr7 157461436 N chr7 157461651 N DEL 7
A00297:158:HT275DSXX:2:1339:12337:24173 chr7 157461547 N chr7 157461678 N DEL 17
A00404:156:HV37TDSXX:3:2518:9751:19225 chr7 157461547 N chr7 157461678 N DEL 21
A00404:155:HV27LDSXX:1:2349:23285:11443 chr7 157461460 N chr7 157461647 N DEL 8
A00404:155:HV27LDSXX:4:1474:1353:24909 chr7 157461495 N chr7 157461764 N DUP 16
A00404:156:HV37TDSXX:2:1302:30924:15280 chr7 157461694 N chr7 157461837 N DUP 15
A00297:158:HT275DSXX:4:1577:23086:35430 chr7 157461442 N chr7 157461727 N DEL 10
A00297:158:HT275DSXX:2:2317:15619:20964 chr7 157461745 N chr7 157461834 N DUP 15
A00404:156:HV37TDSXX:2:1616:28049:30436 chr7 157461457 N chr7 157461784 N DEL 20
A00404:155:HV27LDSXX:4:2162:5412:5760 chr7 157461781 N chr7 157461834 N DUP 15
A00404:156:HV37TDSXX:4:1156:25364:31579 chr7 157461429 N chr7 157461786 N DEL 5
A00297:158:HT275DSXX:2:2375:16758:31955 chr7 157461758 N chr7 157461819 N DEL 5
A00404:156:HV37TDSXX:2:1225:13096:33317 chr4 73757857 N chr4 73757994 N DUP 5
A00404:155:HV27LDSXX:1:1567:25825:34726 chr9 64939140 N chr9 64939358 N DUP 5
A00297:158:HT275DSXX:3:2218:1262:17613 chr7 72766676 N chr7 72766988 N DUP 4
A00297:158:HT275DSXX:3:2218:1750:16297 chr7 72766676 N chr7 72766988 N DUP 4
A00404:155:HV27LDSXX:3:2472:5638:17644 chr7 72766677 N chr7 72766989 N DUP 3
A00404:156:HV37TDSXX:1:1656:24144:35070 chr1 228438416 N chr1 228438666 N DUP 5
A00404:155:HV27LDSXX:3:2226:17842:10942 chr1 228438777 N chr1 228438983 N DEL 5
A00404:156:HV37TDSXX:1:1656:24144:35070 chr1 228438514 N chr1 228438766 N DEL 10
A00404:155:HV27LDSXX:2:2309:13675:19382 chr1 228438799 N chr1 228438964 N DEL 50
A00404:156:HV37TDSXX:2:1578:20066:15201 chr4 49546163 N chr4 49546607 N DEL 5
A00404:156:HV37TDSXX:3:2239:13078:35102 chr4 49546289 N chr4 49546581 N DUP 2
A00404:155:HV27LDSXX:3:1161:6352:31751 chr19 48342438 N chr19 48342492 N DEL 5
A00404:155:HV27LDSXX:4:2174:26784:21136 chr19 48342438 N chr19 48342492 N DEL 9
A00404:155:HV27LDSXX:4:2515:5249:28933 chr19 48342438 N chr19 48342492 N DEL 12
A00297:158:HT275DSXX:1:2367:16866:22874 chr12 129817996 N chr12 129818188 N DUP 5
A00404:156:HV37TDSXX:4:2560:18448:8140 chr12 131259393 N chr12 131259450 N DEL 5
A00404:155:HV27LDSXX:3:2116:23375:25504 chr12 131259393 N chr12 131259450 N DEL 5
A00404:155:HV27LDSXX:1:2457:27489:24643 chr12 131259397 N chr12 131259454 N DEL 5
A00404:156:HV37TDSXX:4:2468:22254:1830 chr12 131259430 N chr12 131259487 N DEL 10
A00404:155:HV27LDSXX:1:1610:12915:37043 chr12 131259483 N chr12 131259614 N DUP 3
A00404:155:HV27LDSXX:2:1657:9842:36041 chr12 131259521 N chr12 131259594 N DEL 9
A00297:158:HT275DSXX:4:2102:22101:36104 chr12 131259714 N chr12 131260095 N DEL 2
A00297:158:HT275DSXX:2:1254:11550:27853 chr12 131259427 N chr12 131259860 N DEL 24
A00297:158:HT275DSXX:4:1667:22887:5055 chr12 131259798 N chr12 131260035 N DEL 5
A00404:155:HV27LDSXX:2:2363:8910:9721 chr12 131259400 N chr12 131259741 N DEL 5
A00297:158:HT275DSXX:1:1576:14633:5071 chr12 131259798 N chr12 131260035 N DEL 3
A00297:158:HT275DSXX:1:2426:28040:12226 chr12 131259826 N chr12 131260035 N DEL 6
A00404:155:HV27LDSXX:3:2510:11785:32111 chr12 131259826 N chr12 131260035 N DEL 10
A00297:158:HT275DSXX:2:2466:6668:2613 chr12 131259826 N chr12 131260035 N DEL 5
A00404:155:HV27LDSXX:1:2636:30996:21699 chr12 131259826 N chr12 131260035 N DEL 5
A00297:158:HT275DSXX:4:1518:25753:8422 chr12 131259418 N chr12 131260153 N DUP 8
A00404:156:HV37TDSXX:3:2214:30337:6089 chr12 131259409 N chr12 131260146 N DEL 15
A00404:156:HV37TDSXX:4:2217:21694:36495 chr1 50710782 N chr1 50711090 N DEL 5
A00404:156:HV37TDSXX:3:1475:7771:11350 chr8 43195630 N chr8 43195850 N DEL 5
A00404:155:HV27LDSXX:4:1323:6632:31892 chr8 43195637 N chr8 43195887 N DEL 5
A00404:155:HV27LDSXX:4:1239:2609:36323 chr8 43195680 N chr8 43195808 N DUP 4
A00404:156:HV37TDSXX:4:2123:25238:29637 chr8 43195687 N chr8 43195907 N DEL 7
A00404:156:HV37TDSXX:4:2123:25283:30655 chr8 43195687 N chr8 43195907 N DEL 7
A00404:155:HV27LDSXX:2:1218:29405:27054 chr10 1010186 N chr10 1010343 N DEL 8
A00404:155:HV27LDSXX:4:1504:18466:20854 chr10 1010196 N chr10 1010353 N DEL 5
A00404:155:HV27LDSXX:4:1647:22869:12132 chr2 241815449 N chr2 241815577 N DUP 18
A00404:155:HV27LDSXX:1:1571:11605:35837 chr2 241815425 N chr2 241815510 N DUP 4
A00404:155:HV27LDSXX:1:1451:20193:18803 chr2 241815444 N chr2 241815572 N DUP 15
A00297:158:HT275DSXX:3:1407:5737:29935 chr2 241815451 N chr2 241815536 N DUP 6
A00297:158:HT275DSXX:3:1407:6397:28510 chr2 241815451 N chr2 241815536 N DUP 6
A00404:156:HV37TDSXX:2:1678:22245:22639 chr2 241815487 N chr2 241815572 N DUP 12
A00404:156:HV37TDSXX:2:2525:17635:15718 chr2 241815444 N chr2 241815572 N DUP 28
A00404:156:HV37TDSXX:2:2345:15501:16376 chr19 15887392 N chr19 15887813 N DEL 4
A00297:158:HT275DSXX:3:1353:14091:6261 chr19 15887392 N chr19 15887813 N DEL 5
A00404:155:HV27LDSXX:3:2546:9344:8719 chr19 15887522 N chr19 15887941 N DUP 5
A00404:156:HV37TDSXX:3:1273:27615:6762 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:3:1371:15790:24674 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:1:1106:31421:30138 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:4:1549:31078:16203 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:4:1549:31087:16219 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:1:2530:25997:28635 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:3:2160:27905:17973 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:3:1133:17616:13307 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:4:1641:21685:14653 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:4:2641:20934:14011 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:1:2104:31882:6731 chr19 15887522 N chr19 15887941 N DUP 5
A00404:156:HV37TDSXX:1:2524:4942:30718 chr19 15887556 N chr19 15887977 N DEL 4
A00404:156:HV37TDSXX:4:1641:21450:29528 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:2:2251:1904:7545 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:4:1215:15338:8516 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:3:1505:16604:31532 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:1:1657:21359:27273 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:1:2657:21423:2487 chr19 15887522 N chr19 15887941 N DUP 5
A00404:156:HV37TDSXX:2:1427:7283:1673 chr19 15887522 N chr19 15887941 N DUP 5
A00404:156:HV37TDSXX:3:2568:16848:26694 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:4:1411:6741:9940 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:4:2421:13711:33974 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:2:1272:25554:6292 chr19 15887522 N chr19 15887941 N DUP 5
A00297:158:HT275DSXX:1:1434:22860:33880 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:3:2431:23800:21136 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:3:2431:24062:21966 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:2:1521:28881:27179 chr19 15887522 N chr19 15887941 N DUP 5
A00404:155:HV27LDSXX:2:1637:18656:6433 chr19 15887522 N chr19 15887941 N DUP 5
A00404:156:HV37TDSXX:2:1421:6524:3114 chr19 15887523 N chr19 15887942 N DUP 5
A00297:158:HT275DSXX:3:1604:16080:23077 chr19 15887528 N chr19 15887947 N DUP 5
A00297:158:HT275DSXX:1:2448:18900:15530 chr19 15887534 N chr19 15887953 N DUP 3
A00297:158:HT275DSXX:4:2273:5873:26694 chr19 15887535 N chr19 15887954 N DUP 2
A00404:156:HV37TDSXX:2:2509:2555:31970 chr19 15887535 N chr19 15887954 N DUP 2
A00297:158:HT275DSXX:3:1231:28348:8970 chr19 15887224 N chr19 15887674 N DUP 1
A00404:155:HV27LDSXX:3:2318:2618:10222 chr19 15887444 N chr19 15887685 N DUP 5
A00404:155:HV27LDSXX:3:1133:17616:13307 chr19 15887684 N chr19 15887863 N DEL 15
A00297:158:HT275DSXX:4:1619:25970:19570 chr19 15887723 N chr19 15888062 N DEL 9
A00404:156:HV37TDSXX:3:1231:32208:17942 chr19 15887418 N chr19 15887839 N DEL 1
A00404:156:HV37TDSXX:2:2509:2555:31970 chr19 15887940 N chr19 15888870 N DUP 5
A00404:155:HV27LDSXX:3:1103:18267:16689 chr19 15887437 N chr19 15888106 N DUP 5
A00404:155:HV27LDSXX:3:2322:23493:27461 chr19 15888271 N chr19 15888432 N DEL 5
A00297:158:HT275DSXX:4:1619:25970:19570 chr19 15887407 N chr19 15888166 N DEL 4
A00404:155:HV27LDSXX:2:2156:12879:26083 chr19 15888323 N chr19 15888648 N DUP 5
A00404:155:HV27LDSXX:2:2204:30364:25895 chr19 15887381 N chr19 15888470 N DUP 5
A00404:156:HV37TDSXX:1:2229:6271:18208 chr19 15887564 N chr19 15888643 N DEL 5
A00404:155:HV27LDSXX:4:1505:21748:5087 chr19 15888253 N chr19 15888664 N DEL 5
A00404:156:HV37TDSXX:3:2347:9100:12493 chr16 80411123 N chr16 80411200 N DEL 5
A00404:156:HV37TDSXX:4:2502:20085:20400 chr16 80411123 N chr16 80411200 N DEL 5
A00404:156:HV37TDSXX:2:2216:14371:1611 chr16 80411121 N chr16 80411200 N DEL 12
A00404:155:HV27LDSXX:2:1315:8621:23719 chr16 80411163 N chr16 80411238 N DUP 27
A00404:156:HV37TDSXX:1:2619:22019:20055 chr16 80411163 N chr16 80411238 N DUP 26
A00404:155:HV27LDSXX:2:1473:4598:14559 chr16 80411177 N chr16 80411238 N DUP 43
A00297:158:HT275DSXX:2:1667:6976:3583 chr16 80411124 N chr16 80411237 N DUP 15
A00297:158:HT275DSXX:1:2135:4535:5525 chr16 80411163 N chr16 80411238 N DUP 12
A00297:158:HT275DSXX:1:2135:4535:5556 chr16 80411163 N chr16 80411238 N DUP 12
A00297:158:HT275DSXX:2:2123:26332:4977 chr16 80411124 N chr16 80411237 N DUP 17
A00297:158:HT275DSXX:2:2206:1172:28103 chr16 80411177 N chr16 80411238 N DUP 30
A00404:156:HV37TDSXX:4:1405:9444:15280 chr16 80411163 N chr16 80411238 N DUP 7
A00297:158:HT275DSXX:2:2330:21305:29997 chr16 80411124 N chr16 80411237 N DUP 15
A00404:156:HV37TDSXX:1:1478:7609:9596 chr16 80411134 N chr16 80411209 N DUP 5
A00404:156:HV37TDSXX:4:2266:16631:26130 chr16 80411163 N chr16 80411238 N DUP 19
A00404:155:HV27LDSXX:4:1255:13530:33630 chr16 80411163 N chr16 80411238 N DUP 19
A00297:158:HT275DSXX:2:1169:23520:1141 chr16 80411163 N chr16 80411238 N DUP 20
A00404:155:HV27LDSXX:2:1243:29333:29121 chr16 80411163 N chr16 80411238 N DUP 21
A00297:158:HT275DSXX:2:2469:3441:10864 chr16 80411163 N chr16 80411238 N DUP 22
A00404:156:HV37TDSXX:2:2131:16495:23829 chr16 80411163 N chr16 80411238 N DUP 23
A00404:155:HV27LDSXX:4:2161:1669:25300 chr16 80411163 N chr16 80411238 N DUP 25
A00404:156:HV37TDSXX:2:1352:24677:21402 chr16 80411190 N chr16 80411248 N DUP 9
A00297:158:HT275DSXX:2:2641:2085:22451 chr16 80411163 N chr16 80411238 N DUP 27
A00297:158:HT275DSXX:1:1639:22516:19507 chr10 132651447 N chr10 132651676 N DUP 1
A00297:158:HT275DSXX:4:2573:2672:3521 chr10 132651474 N chr10 132651613 N DEL 5
A00297:158:HT275DSXX:1:1340:21549:16078 chr10 132651445 N chr10 132651630 N DEL 15
A00404:156:HV37TDSXX:4:1378:28085:16188 chr3 123607550 N chr3 123607679 N DEL 2
A00404:155:HV27LDSXX:2:1406:25934:6042 chr3 123607733 N chr3 123607906 N DUP 7
A00404:155:HV27LDSXX:2:2246:1280:4773 chr3 123607539 N chr3 123607948 N DEL 7
A00404:155:HV27LDSXX:2:2645:9263:18756 chr7 5538878 N chr7 5538981 N DEL 33
A00297:158:HT275DSXX:1:1205:20148:10582 chr13 18614717 N chr13 18615175 N DUP 5
A00297:158:HT275DSXX:1:1205:21359:29528 chr13 18614717 N chr13 18615175 N DUP 5
A00404:155:HV27LDSXX:3:2411:13964:24580 chr13 18614718 N chr13 18615072 N DUP 5
A00404:156:HV37TDSXX:2:1266:23647:22686 chr13 18614720 N chr13 18615481 N DUP 5
A00404:156:HV37TDSXX:4:2458:7175:13260 chr13 113375366 N chr13 113375967 N DEL 10
A00404:156:HV37TDSXX:2:1610:10429:17049 chr13 113375305 N chr13 113375416 N DEL 5
A00297:158:HT275DSXX:2:2216:19434:6089 chr13 113375438 N chr13 113375517 N DUP 5
A00404:155:HV27LDSXX:3:2317:1353:16767 chr13 113375440 N chr13 113375919 N DUP 5
A00297:158:HT275DSXX:3:2445:32805:16908 chr13 113375580 N chr13 113376001 N DEL 5
A00404:156:HV37TDSXX:4:2118:10827:30232 chr13 113376001 N chr13 113376080 N DUP 17
A00297:158:HT275DSXX:3:1429:6551:7138 chr13 113375580 N chr13 113376001 N DEL 9
A00404:155:HV27LDSXX:4:1434:17029:29074 chr13 113375580 N chr13 113376001 N DEL 10
A00404:156:HV37TDSXX:1:2155:15338:9455 chr13 113375340 N chr13 113376001 N DEL 10
A00404:156:HV37TDSXX:1:2643:1380:31062 chr13 113375856 N chr13 113375935 N DUP 5
A00297:158:HT275DSXX:4:1531:29405:13933 chr13 113375535 N chr13 113375856 N DEL 1
A00297:158:HT275DSXX:3:1144:25807:19914 chr13 113375341 N chr13 113376082 N DEL 1
A00297:158:HT275DSXX:2:2236:28492:20243 chr13 113375679 N chr13 113376018 N DUP 5
A00297:158:HT275DSXX:2:2218:28284:10551 chr13 113375340 N chr13 113376001 N DEL 10
A00297:158:HT275DSXX:4:1529:22733:9455 chr13 113375346 N chr13 113376007 N DEL 5
A00404:156:HV37TDSXX:4:1217:9643:4789 chr13 113376001 N chr13 113376080 N DUP 15
A00404:155:HV27LDSXX:3:1605:2220:23782 chr13 113375341 N chr13 113376082 N DEL 4
A00404:156:HV37TDSXX:3:1478:5050:6543 chr13 113376130 N chr13 113376358 N DEL 25
A00404:156:HV37TDSXX:1:2249:29478:4726 chr13 113375561 N chr13 113376241 N DEL 1
A00404:156:HV37TDSXX:1:1648:21088:32127 chr12 110173183 N chr12 110173309 N DUP 5
A00404:156:HV37TDSXX:1:1648:21106:32095 chr12 110173183 N chr12 110173309 N DUP 5
A00297:158:HT275DSXX:1:2264:9896:17315 chr12 110173266 N chr12 110173362 N DUP 10
A00297:158:HT275DSXX:3:1231:11577:10269 chr3 49938856 N chr3 49939019 N DEL 23
A00404:156:HV37TDSXX:4:1436:25934:25019 chr18 72354569 N chr18 72354650 N DEL 39
A00404:156:HV37TDSXX:3:1108:5556:28933 chr18 72354535 N chr18 72354614 N DUP 17
A00404:156:HV37TDSXX:2:1166:3242:37012 chr18 72354593 N chr18 72354658 N DEL 15
A00297:158:HT275DSXX:4:2170:14398:24424 chr18 72354594 N chr18 72354667 N DEL 5
A00297:158:HT275DSXX:4:2171:19416:15201 chr18 72354594 N chr18 72354667 N DEL 5
A00404:155:HV27LDSXX:3:1225:17761:34413 chr10 34010312 N chr10 34010541 N DEL 6
A00297:158:HT275DSXX:2:2245:18376:9111 chr10 34010312 N chr10 34010541 N DEL 7
A00404:155:HV27LDSXX:3:1340:12744:35556 chr10 34010312 N chr10 34010541 N DEL 7
A00404:156:HV37TDSXX:4:1260:4761:33755 chr10 34010375 N chr10 34010460 N DUP 12
A00297:158:HT275DSXX:3:1126:14226:6308 chr10 34010375 N chr10 34010460 N DUP 13
A00404:156:HV37TDSXX:4:2106:28537:21418 chr10 34010397 N chr10 34010466 N DUP 13
A00297:158:HT275DSXX:1:2603:30463:4617 chr10 34010397 N chr10 34010466 N DUP 13
A00404:156:HV37TDSXX:4:2131:30761:19194 chr10 34010397 N chr10 34010466 N DUP 13
A00297:158:HT275DSXX:1:1347:2094:31548 chr10 34010397 N chr10 34010466 N DUP 13
A00404:155:HV27LDSXX:3:2623:27751:16297 chr10 34010397 N chr10 34010466 N DUP 13
A00404:156:HV37TDSXX:2:2266:25599:16736 chr10 34010397 N chr10 34010466 N DUP 13
A00297:158:HT275DSXX:2:2124:21341:28025 chr10 34010397 N chr10 34010466 N DUP 13
A00404:155:HV27LDSXX:2:2225:27498:17989 chr10 34010397 N chr10 34010466 N DUP 13
A00404:156:HV37TDSXX:1:1219:20003:32565 chr10 34010397 N chr10 34010466 N DUP 13
A00404:155:HV27LDSXX:3:1320:9155:10113 chr10 34010397 N chr10 34010466 N DUP 13
A00297:158:HT275DSXX:3:1117:4399:28902 chr10 34010442 N chr10 34010512 N DEL 8
A00404:155:HV27LDSXX:3:1421:29017:1423 chr10 34010442 N chr10 34010512 N DEL 8
A00297:158:HT275DSXX:2:1304:5312:3677 chr10 34010442 N chr10 34010512 N DEL 8
A00404:155:HV27LDSXX:2:1649:4237:14904 chr10 34010442 N chr10 34010512 N DEL 8
A00297:158:HT275DSXX:3:1314:20166:17785 chr10 34010442 N chr10 34010512 N DEL 8
A00404:156:HV37TDSXX:2:2475:13539:34303 chr10 34010442 N chr10 34010512 N DEL 8
A00297:158:HT275DSXX:2:2125:5746:30859 chr11 126259774 N chr11 126260070 N DEL 4
A00297:158:HT275DSXX:1:2111:21251:14058 chr11 126259790 N chr11 126260086 N DEL 1
A00297:158:HT275DSXX:1:1406:9977:31955 chr3 196334966 N chr3 196335037 N DEL 5
A00404:155:HV27LDSXX:1:2507:21386:33552 chr3 196334967 N chr3 196335108 N DEL 1
A00404:155:HV27LDSXX:4:2202:30400:11522 chr3 196334967 N chr3 196335108 N DEL 7
A00404:155:HV27LDSXX:2:2166:11162:7764 chr3 196334967 N chr3 196335108 N DEL 7
A00297:158:HT275DSXX:2:1338:15411:6230 chr3 196335115 N chr3 196335185 N DUP 7
A00404:155:HV27LDSXX:2:2448:27299:29168 chr3 196335118 N chr3 196335188 N DUP 7
A00404:155:HV27LDSXX:3:2610:2175:12273 chr3 196335115 N chr3 196335185 N DUP 5
A00297:158:HT275DSXX:1:2455:5412:17597 chr3 196335115 N chr3 196335185 N DUP 1
A00297:158:HT275DSXX:1:1606:13919:29575 chr3 196335201 N chr3 196335551 N DEL 21
A00404:156:HV37TDSXX:4:1244:5068:33004 chr3 196335480 N chr3 196335551 N DEL 12
A00404:156:HV37TDSXX:1:1136:10827:4335 chr3 196335027 N chr3 196335657 N DEL 2
A00404:155:HV27LDSXX:3:1511:24469:33191 chr3 196335577 N chr3 196335683 N DEL 20
A00297:158:HT275DSXX:1:2422:27064:8625 chr21 45141950 N chr21 45142183 N DUP 5
A00297:158:HT275DSXX:4:2418:13214:14575 chr4 126101423 N chr4 126101580 N DUP 4
A00297:158:HT275DSXX:4:2418:13376:14231 chr4 126101423 N chr4 126101580 N DUP 4
A00404:155:HV27LDSXX:3:1356:31295:20901 chr4 126101393 N chr4 126101580 N DUP 4
A00404:156:HV37TDSXX:2:1263:24442:28416 chr4 126101389 N chr4 126101538 N DEL 7
A00404:155:HV27LDSXX:1:1557:21197:31626 chr4 126101524 N chr4 126101593 N DEL 6
A00297:158:HT275DSXX:1:2607:3794:22999 chr5 46434985 N chr5 46436050 N DEL 15
A00404:156:HV37TDSXX:3:1429:25816:25755 chr5 46434991 N chr5 46436048 N DEL 15
A00404:155:HV27LDSXX:3:1108:5701:26741 chr5 46434994 N chr5 46436050 N DEL 15
A00404:155:HV27LDSXX:2:1626:2799:7435 chr5 46434996 N chr5 46436049 N DEL 15
A00297:158:HT275DSXX:3:2628:24939:8703 chr5 46434999 N chr5 46436050 N DEL 15
A00297:158:HT275DSXX:1:1444:20039:16971 chr5 46435002 N chr5 46436049 N DEL 15
A00297:158:HT275DSXX:1:2444:17870:16376 chr5 46435002 N chr5 46436049 N DEL 15
A00297:158:HT275DSXX:3:2651:26684:7435 chr5 46435052 N chr5 46436049 N DEL 10
A00297:158:HT275DSXX:4:1648:11180:1908 chr5 46435052 N chr5 46436049 N DEL 5
A00404:155:HV27LDSXX:4:1507:30843:13135 chr5 46435052 N chr5 46436049 N DEL 10
A00404:155:HV27LDSXX:1:1163:24912:20650 chr5 46435054 N chr5 46436049 N DEL 5
A00404:155:HV27LDSXX:1:2373:3531:35196 chr5 46435054 N chr5 46436049 N DEL 5
A00404:156:HV37TDSXX:2:1630:4878:26256 chr5 46435054 N chr5 46436049 N DEL 13
A00404:156:HV37TDSXX:2:2467:22327:5087 chr5 46435057 N chr5 46436050 N DEL 15
A00404:156:HV37TDSXX:3:1669:27389:23844 chr5 46435059 N chr5 46436049 N DEL 5
A00297:158:HT275DSXX:4:2416:18258:1266 chr5 46435059 N chr5 46436049 N DEL 5
A00297:158:HT275DSXX:4:2119:17119:16861 chr5 46435060 N chr5 46436049 N DEL 19
A00404:155:HV27LDSXX:2:1238:10773:21057 chr5 46435065 N chr5 46436050 N DEL 6
A00404:156:HV37TDSXX:1:2523:17616:30029 chr5 46435065 N chr5 46436050 N DEL 6
A00297:158:HT275DSXX:3:2355:7464:13667 chr5 46435069 N chr5 46436049 N DEL 10
A00404:156:HV37TDSXX:1:2117:26503:9251 chr5 46435071 N chr5 46436050 N DEL 10
A00297:158:HT275DSXX:2:1201:23466:17581 chr5 46435129 N chr5 46436049 N DEL 20
A00404:156:HV37TDSXX:4:2405:29903:26130 chr5 46435138 N chr5 46436050 N DEL 20
A00404:155:HV27LDSXX:4:2407:8431:23015 chr5 46435140 N chr5 46436050 N DEL 25
A00404:156:HV37TDSXX:3:1442:2049:22044 chr5 46435140 N chr5 46436050 N DEL 25
A00404:156:HV37TDSXX:3:2516:30553:13698 chr5 46435140 N chr5 46436050 N DEL 25
A00404:155:HV27LDSXX:3:2546:21088:22701 chr5 46435149 N chr5 46436049 N DEL 25
A00297:158:HT275DSXX:3:1140:32904:8030 chr5 46435151 N chr5 46436050 N DEL 20
A00297:158:HT275DSXX:3:2139:30861:34084 chr5 46435151 N chr5 46436050 N DEL 20
A00297:158:HT275DSXX:3:2628:24939:8703 chr5 46435157 N chr5 46436048 N DEL 30
A00404:156:HV37TDSXX:1:1415:9218:8844 chr5 46435161 N chr5 46436048 N DEL 27
A00404:156:HV37TDSXX:2:2101:17291:18255 chr5 46435166 N chr5 46436050 N DEL 35
A00404:156:HV37TDSXX:2:2423:18936:5603 chr5 46435166 N chr5 46436050 N DEL 35
A00404:156:HV37TDSXX:2:2412:7021:29089 chr7 333907 N chr7 334062 N DEL 16
A00297:158:HT275DSXX:3:1311:6831:20713 chr7 333999 N chr7 334314 N DEL 1
A00297:158:HT275DSXX:3:2217:22200:35931 chr7 333918 N chr7 334125 N DUP 5
A00404:155:HV27LDSXX:4:1663:22896:14121 chr7 334047 N chr7 334458 N DEL 9
A00404:156:HV37TDSXX:4:2134:13792:13322 chr7 334077 N chr7 334444 N DEL 12
A00404:155:HV27LDSXX:2:1239:24135:27978 chr7 333914 N chr7 334173 N DUP 4
A00404:155:HV27LDSXX:2:1122:23565:30686 chr7 334068 N chr7 334479 N DUP 9
A00297:158:HT275DSXX:3:2150:4960:16971 chr7 333958 N chr7 334173 N DUP 5
A00297:158:HT275DSXX:2:1516:27633:1720 chr7 333960 N chr7 334175 N DUP 5
A00404:156:HV37TDSXX:1:2637:20663:27226 chr7 333958 N chr7 334173 N DUP 5
A00297:158:HT275DSXX:2:2602:4490:36072 chr7 333928 N chr7 334189 N DEL 5
A00404:156:HV37TDSXX:3:1135:12029:19319 chr7 334013 N chr7 334230 N DEL 3
A00404:156:HV37TDSXX:4:2220:5213:6543 chr7 334313 N chr7 334522 N DEL 25
A00297:158:HT275DSXX:2:2316:15881:5603 chr7 333940 N chr7 334299 N DEL 4
A00404:156:HV37TDSXX:2:2145:31512:36714 chr7 334475 N chr7 334596 N DEL 7
A00404:155:HV27LDSXX:2:2164:27724:19038 chr7 334465 N chr7 334522 N DEL 28
A00297:158:HT275DSXX:2:1620:30219:15060 chr7 334527 N chr7 334646 N DEL 5
A00404:156:HV37TDSXX:3:1476:5484:30718 chr8 11026289 N chr8 11026425 N DEL 16
A00404:155:HV27LDSXX:2:2359:24623:28260 chr8 11026395 N chr8 11026695 N DEL 5
A00404:155:HV27LDSXX:2:2359:24623:28260 chr8 11026307 N chr8 11026607 N DEL 15
A00404:156:HV37TDSXX:3:2177:23194:15702 chr8 11026396 N chr8 11026569 N DUP 5
A00404:155:HV27LDSXX:3:2347:11903:8609 chr8 11026356 N chr8 11026407 N DEL 5
A00404:155:HV27LDSXX:3:2674:7093:11240 chr8 11026325 N chr8 11026401 N DEL 5
A00404:155:HV27LDSXX:3:2608:1163:5196 chr8 11026544 N chr8 11026595 N DEL 2
A00297:158:HT275DSXX:3:1517:14488:19257 chr8 11026339 N chr8 11026589 N DEL 5
A00404:155:HV27LDSXX:2:1213:11966:18145 chr8 11026595 N chr8 11026743 N DUP 15
A00404:156:HV37TDSXX:2:1673:30174:10755 chr8 11026396 N chr8 11026596 N DEL 5
A00404:155:HV27LDSXX:3:2674:7093:11240 chr8 11026323 N chr8 11026598 N DEL 7
A00404:156:HV37TDSXX:4:2667:6804:12900 chr8 11026328 N chr8 11026603 N DEL 6
A00404:155:HV27LDSXX:1:1239:9435:18709 chr8 11026396 N chr8 11026694 N DUP 5
A00297:158:HT275DSXX:3:1657:11442:1861 chr8 11026517 N chr8 11026740 N DUP 5
A00404:156:HV37TDSXX:1:1111:20826:12915 chr8 11026750 N chr8 11026950 N DEL 5
A00297:158:HT275DSXX:3:2103:30671:13463 chr8 11026595 N chr8 11026743 N DUP 5
A00297:158:HT275DSXX:4:2342:1298:1423 chr8 11026595 N chr8 11026743 N DUP 5
A00297:158:HT275DSXX:3:1374:8015:22514 chr8 11026723 N chr8 11026998 N DEL 8
A00404:156:HV37TDSXX:4:2551:11568:4492 chr8 11026642 N chr8 11027139 N DUP 4
A00404:155:HV27LDSXX:1:2605:6370:32127 chr8 11026595 N chr8 11026743 N DUP 4
A00404:155:HV27LDSXX:1:1635:30969:11287 chr8 11026595 N chr8 11026743 N DUP 5
A00404:155:HV27LDSXX:1:1401:31955:1846 chr8 11026595 N chr8 11026743 N DUP 5
A00297:158:HT275DSXX:2:2529:25364:22874 chr8 11026595 N chr8 11026743 N DUP 13
A00297:158:HT275DSXX:2:2455:25771:9612 chr8 11026595 N chr8 11026743 N DUP 27
A00404:155:HV27LDSXX:4:1248:32181:34147 chr8 11026595 N chr8 11026743 N DUP 30
A00404:155:HV27LDSXX:2:1358:31638:36839 chr8 11026595 N chr8 11026743 N DUP 20
A00404:156:HV37TDSXX:2:2153:20419:26647 chr8 11026687 N chr8 11026911 N DEL 5
A00404:156:HV37TDSXX:1:1516:25418:20744 chr8 11026327 N chr8 11026923 N DUP 10
A00404:156:HV37TDSXX:1:1111:20826:12915 chr8 11026537 N chr8 11026959 N DUP 10
A00297:158:HT275DSXX:3:1230:20654:19257 chr8 11026595 N chr8 11026967 N DUP 10
A00404:155:HV27LDSXX:3:2274:20600:7106 chr8 11026595 N chr8 11026967 N DUP 10
A00404:156:HV37TDSXX:3:2575:9209:6480 chr8 11026587 N chr8 11026959 N DUP 10
A00404:156:HV37TDSXX:1:1541:22851:29919 chr8 11026321 N chr8 11027067 N DUP 1
A00404:156:HV37TDSXX:4:2667:6804:12900 chr8 11026355 N chr8 11027003 N DEL 10
A00297:158:HT275DSXX:4:2531:5339:10238 chr8 11026347 N chr8 11026995 N DEL 10
A00297:158:HT275DSXX:2:1620:19605:16689 chr8 11026328 N chr8 11027001 N DEL 9
A00297:158:HT275DSXX:4:1522:9236:16986 chr8 11026336 N chr8 11027009 N DEL 1
A00404:155:HV27LDSXX:2:1636:31448:26490 chr8 11026366 N chr8 11027114 N DEL 5
A00297:158:HT275DSXX:3:1513:22761:36683 chr8 11026366 N chr8 11027114 N DEL 5
A00297:158:HT275DSXX:4:1301:30327:35947 chr3 48734085 N chr3 48734242 N DEL 4
A00404:155:HV27LDSXX:3:2210:11089:20040 chr3 48734058 N chr3 48734175 N DEL 34
A00404:155:HV27LDSXX:3:2210:14281:22060 chr3 48734058 N chr3 48734175 N DEL 34
A00297:158:HT275DSXX:4:1301:30327:35947 chr3 48734085 N chr3 48734242 N DEL 15
A00404:156:HV37TDSXX:2:1359:31186:1329 chr3 48734225 N chr3 48734340 N DUP 10
A00297:158:HT275DSXX:4:1126:5846:36198 chr3 48734138 N chr3 48734332 N DEL 10
A00297:158:HT275DSXX:1:1246:25409:32095 chr3 48734074 N chr3 48734347 N DEL 18
A00297:158:HT275DSXX:3:1313:18313:28416 chrX 76218656 N chrX 76218851 N DUP 5
A00404:155:HV27LDSXX:2:1118:8449:6699 chr2 202215769 N chr2 202216113 N DEL 5
A00404:156:HV37TDSXX:1:2665:25120:7326 chr2 202215769 N chr2 202216113 N DEL 5
A00297:158:HT275DSXX:3:1221:29378:31297 chr2 202215782 N chr2 202215917 N DUP 5
A00404:156:HV37TDSXX:3:1437:21630:24048 chr2 202215786 N chr2 202216128 N DUP 3
A00297:158:HT275DSXX:2:1222:26702:22686 chr2 202216046 N chr2 202216385 N DEL 1
A00404:155:HV27LDSXX:2:2477:18050:35164 chr15 74334467 N chr15 74334612 N DEL 10
A00297:158:HT275DSXX:2:2136:30110:30624 chr15 74334449 N chr15 74334642 N DEL 20
A00404:156:HV37TDSXX:4:1272:3396:24784 chr15 74334336 N chr15 74334457 N DEL 5
A00404:156:HV37TDSXX:1:1620:26512:19445 chr15 74334274 N chr15 74334467 N DEL 4
A00404:156:HV37TDSXX:3:1627:8567:24439 chr15 74334585 N chr15 74334706 N DEL 10
A00404:155:HV27LDSXX:2:2142:21856:7279 chr15 74334543 N chr15 74334831 N DEL 21
A00297:158:HT275DSXX:4:1413:32434:36902 chr15 74334436 N chr15 74334844 N DEL 2
A00297:158:HT275DSXX:3:2621:3432:9064 chr7 102512799 N chr7 102512906 N DUP 7
A00297:158:HT275DSXX:3:1122:26268:1830 chr7 102512937 N chr7 102513010 N DUP 6
A00404:156:HV37TDSXX:2:2551:9480:27305 chr7 102512946 N chr7 102513007 N DEL 30
A00404:156:HV37TDSXX:1:2543:5132:6433 chr8 78524041 N chr8 78524098 N DUP 5
A00404:155:HV27LDSXX:4:2243:29903:2080 chr7 107680001 N chr7 107680052 N DEL 11
A00404:155:HV27LDSXX:4:1526:7844:19586 chr7 107679961 N chr7 107680053 N DEL 11
A00404:155:HV27LDSXX:3:1322:21802:17989 chr7 107679966 N chr7 107680058 N DEL 9
A00404:155:HV27LDSXX:2:2629:27326:12680 chr7 107679967 N chr7 107680059 N DEL 8
A00404:156:HV37TDSXX:2:1427:4137:18333 chr7 107680160 N chr7 107680266 N DEL 10
A00404:156:HV37TDSXX:4:2463:28501:34632 chr7 107679998 N chr7 107680274 N DEL 4
A00404:155:HV27LDSXX:1:2236:25319:2722 chr7 107680092 N chr7 107680272 N DEL 6
A00297:158:HT275DSXX:4:1558:15664:30311 chr7 107680332 N chr7 107680403 N DUP 1
A00297:158:HT275DSXX:1:2655:11632:35822 chr7 107679970 N chr7 107680444 N DUP 10
A00404:156:HV37TDSXX:3:2466:23213:2362 chr7 107680434 N chr7 107680530 N DEL 10
A00404:156:HV37TDSXX:1:1149:15040:26287 chr7 107680434 N chr7 107680530 N DEL 10
A00404:156:HV37TDSXX:3:2318:31647:20509 chr7 107679987 N chr7 107680450 N DEL 15
A00404:156:HV37TDSXX:2:1164:9073:5932 chr7 107679987 N chr7 107680450 N DEL 15
A00297:158:HT275DSXX:1:1260:29080:21699 chr7 107679987 N chr7 107680450 N DEL 15
A00297:158:HT275DSXX:1:1260:29369:22608 chr7 107679987 N chr7 107680450 N DEL 15
A00297:158:HT275DSXX:1:1261:29803:2973 chr7 107679987 N chr7 107680450 N DEL 15
A00297:158:HT275DSXX:1:2163:11062:32988 chr7 107679987 N chr7 107680450 N DEL 15
A00404:156:HV37TDSXX:1:2172:13838:8672 chr7 107679965 N chr7 107680451 N DEL 14
A00297:158:HT275DSXX:1:2507:9607:25175 chr7 107679968 N chr7 107680454 N DEL 11
A00404:155:HV27LDSXX:4:1471:16929:30968 chr7 107680001 N chr7 107680464 N DEL 1
A00404:155:HV27LDSXX:1:1535:10556:3959 chr7 107680000 N chr7 107680481 N DEL 5
A00297:158:HT275DSXX:3:2228:31087:1188 chr19 4185152 N chr19 4185370 N DEL 14
A00404:156:HV37TDSXX:2:2233:13178:18615 chrX 31067067 N chrX 31067384 N DEL 5
A00297:158:HT275DSXX:1:1268:4679:23500 chrX 31067018 N chrX 31067079 N DUP 5
A00404:155:HV27LDSXX:3:1360:5520:13933 chrX 31067018 N chrX 31067079 N DUP 5
A00404:155:HV27LDSXX:1:1468:14443:16047 chrX 31067018 N chrX 31067079 N DUP 5
A00404:155:HV27LDSXX:1:1468:6922:31735 chrX 31067018 N chrX 31067079 N DUP 5
A00297:158:HT275DSXX:1:2460:23113:17879 chrX 31066900 N chrX 31067163 N DEL 17
A00404:155:HV27LDSXX:1:1207:19741:16579 chrX 31067036 N chrX 31067165 N DEL 13
A00404:155:HV27LDSXX:4:1120:17562:25927 chrX 31066900 N chrX 31067163 N DEL 18
A00297:158:HT275DSXX:3:2410:10059:11772 chrX 31067035 N chrX 31067166 N DEL 13
A00297:158:HT275DSXX:3:1536:13856:14935 chrX 31067164 N chrX 31067289 N DUP 9
A00404:155:HV27LDSXX:2:1531:18096:36839 chrX 31067008 N chrX 31067295 N DUP 18
A00404:156:HV37TDSXX:1:1247:22652:35243 chrX 31067036 N chrX 31067167 N DEL 12
A00297:158:HT275DSXX:3:1324:30436:26459 chrX 31067200 N chrX 31067417 N DUP 9
A00404:155:HV27LDSXX:3:2659:11315:20243 chrX 31067164 N chrX 31067289 N DUP 13
A00404:155:HV27LDSXX:3:2109:9272:18020 chrX 31066941 N chrX 31067254 N DEL 10
A00297:158:HT275DSXX:3:1374:32407:5102 chrX 31067004 N chrX 31067373 N DUP 9
A00297:158:HT275DSXX:4:1309:22254:25128 chrX 31066998 N chrX 31067163 N DEL 16
A00297:158:HT275DSXX:4:2657:3224:9079 chrX 31066881 N chrX 31067332 N DEL 7
A00297:158:HT275DSXX:2:1174:20555:22247 chrX 31067084 N chrX 31067335 N DEL 7
A00404:155:HV27LDSXX:1:1652:18267:26490 chr20 24980639 N chr20 24980826 N DEL 30
A00404:155:HV27LDSXX:1:1652:18267:26490 chr20 24980639 N chr20 24980826 N DEL 40
A00404:156:HV37TDSXX:2:2276:15266:24111 chr22 48679099 N chr22 48679315 N DEL 1
A00404:156:HV37TDSXX:2:2544:31593:31970 chr22 48679099 N chr22 48679315 N DEL 6
A00404:155:HV27LDSXX:1:1302:8034:17002 chr22 48679099 N chr22 48679315 N DEL 10
A00297:158:HT275DSXX:2:2177:2184:4930 chr22 48679106 N chr22 48679251 N DUP 10
A00404:155:HV27LDSXX:1:2550:3314:9549 chr22 48679258 N chr22 48679403 N DUP 25
A00297:158:HT275DSXX:3:2523:32461:17253 chr22 48679063 N chr22 48679293 N DUP 41
A00297:158:HT275DSXX:4:2143:32678:2785 chr22 48679063 N chr22 48679293 N DUP 42
A00404:155:HV27LDSXX:4:2106:6334:25238 chr22 48679248 N chr22 48679485 N DUP 17
A00404:155:HV27LDSXX:1:2249:17870:6793 chr22 48679315 N chr22 48679462 N DEL 9
A00404:155:HV27LDSXX:1:2556:8486:34976 chr22 48679052 N chr22 48679290 N DUP 45
A00297:158:HT275DSXX:2:2445:10899:16485 chr22 48679316 N chr22 48679392 N DUP 15
A00404:156:HV37TDSXX:2:2601:15609:20541 chr22 48679249 N chr22 48679342 N DEL 5
A00404:155:HV27LDSXX:3:1131:28791:1658 chr22 48679183 N chr22 48679290 N DUP 11
A00297:158:HT275DSXX:2:2567:1407:27477 chr22 48679271 N chr22 48679393 N DUP 10
A00404:155:HV27LDSXX:4:1411:24370:28729 chr22 48679456 N chr22 48679825 N DEL 10
A00297:158:HT275DSXX:3:1150:8693:16705 chr22 48679385 N chr22 48679593 N DEL 15
A00404:156:HV37TDSXX:3:2626:25852:32863 chr22 48679593 N chr22 48679661 N DUP 5
A00404:155:HV27LDSXX:4:1407:32488:1078 chr22 48679239 N chr22 48679593 N DEL 8
A00297:158:HT275DSXX:3:1267:30183:36824 chr22 48679061 N chr22 48679600 N DEL 5
A00404:155:HV27LDSXX:2:1545:19072:9846 chr22 48679162 N chr22 48679639 N DEL 5
A00404:156:HV37TDSXX:4:2449:27932:9314 chr22 48679686 N chr22 48679825 N DEL 10
A00297:158:HT275DSXX:1:1566:6497:22138 chr22 48679162 N chr22 48679455 N DEL 5
A00404:156:HV37TDSXX:3:2626:25852:32863 chr22 48679477 N chr22 48679593 N DEL 5
A00404:156:HV37TDSXX:2:1502:14434:12179 chr22 48679523 N chr22 48679708 N DEL 5
A00297:158:HT275DSXX:4:2151:27697:21809 chr22 48679523 N chr22 48679708 N DEL 5
A00404:156:HV37TDSXX:2:2437:29152:20040 chr22 48679454 N chr22 48679708 N DEL 5
A00404:156:HV37TDSXX:2:2437:30110:18255 chr22 48679454 N chr22 48679708 N DEL 5
A00404:155:HV27LDSXX:4:1407:32488:1078 chr22 48679454 N chr22 48679708 N DEL 5
A00297:158:HT275DSXX:4:1556:20708:6417 chr22 48679546 N chr22 48679754 N DEL 10
A00297:158:HT275DSXX:1:1355:31412:29590 chr22 48679686 N chr22 48679825 N DEL 10
A00404:155:HV27LDSXX:4:2320:29107:3270 chr22 48679435 N chr22 48679735 N DEL 10
A00297:158:HT275DSXX:2:2160:5728:26443 chr22 48679150 N chr22 48679742 N DEL 4
A00297:158:HT275DSXX:2:1667:5936:12649 chr22 48679846 N chr22 48679901 N DEL 33
A00297:158:HT275DSXX:2:1667:6081:13526 chr22 48679669 N chr22 48679931 N DEL 28
A00404:155:HV27LDSXX:4:1542:3848:24878 chr22 48679569 N chr22 48679946 N DEL 38
A00297:158:HT275DSXX:2:2318:16288:6089 chr22 48679846 N chr22 48679901 N DEL 26
A00297:158:HT275DSXX:2:2318:17463:13291 chr22 48679846 N chr22 48679901 N DEL 26
A00297:158:HT275DSXX:4:2448:21441:35243 chr22 48679140 N chr22 48679901 N DEL 23
A00297:158:HT275DSXX:2:1622:9227:35540 chr22 48679055 N chr22 48679901 N DEL 16
A00404:155:HV27LDSXX:2:1556:3622:18537 chr22 48679152 N chr22 48679913 N DEL 3
A00404:155:HV27LDSXX:1:2445:30246:19961 chr1 13982884 N chr1 13983044 N DUP 5
A00297:158:HT275DSXX:2:1531:27046:25066 chr2 10587240 N chr2 10587299 N DUP 18
A00404:156:HV37TDSXX:2:2646:19497:4100 chr2 10587236 N chr2 10587341 N DUP 6
A00297:158:HT275DSXX:3:2225:13404:15436 chr2 10587271 N chr2 10587368 N DEL 12
A00297:158:HT275DSXX:3:1667:20663:9001 chr2 10587212 N chr2 10587387 N DEL 7
A00297:158:HT275DSXX:2:1203:15094:19648 chr22 44884516 N chr22 44884583 N DEL 1
A00297:158:HT275DSXX:2:2456:28646:1251 chr22 44884516 N chr22 44884583 N DEL 19
A00404:156:HV37TDSXX:1:2373:8169:12571 chr22 44884516 N chr22 44884583 N DEL 20
A00404:156:HV37TDSXX:1:2373:8431:11522 chr22 44884516 N chr22 44884583 N DEL 20
A00404:155:HV27LDSXX:1:1358:20121:18865 chr22 44884516 N chr22 44884583 N DEL 14
A00404:156:HV37TDSXX:4:1470:1090:16501 chr22 44884529 N chr22 44884596 N DEL 2
A00404:156:HV37TDSXX:2:1363:7979:24424 chr22 44884449 N chr22 44884718 N DUP 11
A00297:158:HT275DSXX:4:2254:25880:14935 chr22 44884449 N chr22 44884718 N DUP 11
A00297:158:HT275DSXX:1:1468:9607:32440 chr7 99518991 N chr7 99519292 N DEL 3
A00404:155:HV27LDSXX:2:2273:14832:34882 chr7 99518953 N chr7 99519254 N DEL 24
A00297:158:HT275DSXX:4:2378:20220:17159 chr7 99518820 N chr7 99519420 N DUP 5
A00404:156:HV37TDSXX:4:1173:25518:6386 chr7 99518820 N chr7 99519420 N DUP 5
A00404:155:HV27LDSXX:3:1201:17707:36417 chr7 99518820 N chr7 99519420 N DUP 5
A00404:156:HV37TDSXX:1:2263:22562:36839 chr7 99518820 N chr7 99519420 N DUP 5
A00404:156:HV37TDSXX:3:1308:1334:5650 chr7 99518820 N chr7 99519420 N DUP 5
A00404:155:HV27LDSXX:3:2106:12961:25285 chr7 99518820 N chr7 99519420 N DUP 5
A00297:158:HT275DSXX:4:1460:2130:14043 chr5 58563186 N chr5 58564288 N DEL 5
A00297:158:HT275DSXX:4:1460:2130:14043 chr5 58563206 N chr5 58563854 N DEL 9
A00297:158:HT275DSXX:3:2433:13340:13510 chr5 58563225 N chr5 58564790 N DEL 10
A00404:156:HV37TDSXX:4:1623:5873:4930 chr5 58563358 N chr5 58564042 N DEL 6
A00404:156:HV37TDSXX:3:1216:3016:7467 chr5 58563215 N chr5 58563369 N DEL 10
A00297:158:HT275DSXX:3:1522:16667:12070 chr5 58563684 N chr5 58563951 N DEL 15
A00404:155:HV27LDSXX:2:1448:18828:16783 chr5 58563209 N chr5 58563665 N DEL 2
A00404:156:HV37TDSXX:1:2261:11451:33692 chr5 58563305 N chr5 58563795 N DUP 1
A00297:158:HT275DSXX:2:1528:14552:21934 chr5 58563613 N chr5 58563689 N DEL 25
A00297:158:HT275DSXX:3:1667:32199:17331 chr5 58563490 N chr5 58563872 N DEL 46
A00297:158:HT275DSXX:3:1667:32199:17331 chr5 58563481 N chr5 58563863 N DEL 34
A00404:156:HV37TDSXX:4:2302:21052:35070 chr5 58563988 N chr5 58564102 N DUP 4
A00404:155:HV27LDSXX:4:1542:3070:26193 chr5 58563718 N chr5 58564024 N DEL 4
A00404:156:HV37TDSXX:2:1127:17363:3818 chr5 58564164 N chr5 58564393 N DEL 5
A00404:156:HV37TDSXX:4:2371:29749:22388 chr5 58563327 N chr5 58564161 N DEL 5
A00404:156:HV37TDSXX:4:2278:3152:18944 chr5 58564437 N chr5 58564862 N DEL 22
A00404:156:HV37TDSXX:1:2377:20320:30232 chr5 58564173 N chr5 58564402 N DEL 17
A00404:155:HV27LDSXX:1:2216:24885:18380 chr5 58563738 N chr5 58564537 N DUP 3
A00404:155:HV27LDSXX:2:2417:27814:12868 chr5 58564677 N chr5 58564797 N DEL 12
A00404:156:HV37TDSXX:1:1654:17363:7921 chr5 58563241 N chr5 58564650 N DEL 3
A00404:156:HV37TDSXX:4:1568:21079:33113 chr5 58564420 N chr5 58564843 N DUP 3
A00404:156:HV37TDSXX:3:2153:22634:20807 chr5 58563443 N chr5 58564853 N DUP 5
A00404:156:HV37TDSXX:4:2567:16134:1470 chr5 58563443 N chr5 58564853 N DUP 5
A00404:156:HV37TDSXX:4:1139:13349:4664 chr5 58563443 N chr5 58564853 N DUP 5
A00297:158:HT275DSXX:4:2605:21377:1407 chr5 58564787 N chr5 58564902 N DUP 5
A00404:155:HV27LDSXX:1:2226:22516:7388 chr5 58564184 N chr5 58564800 N DEL 10
A00404:156:HV37TDSXX:4:2278:3152:18944 chr5 58564383 N chr5 58564808 N DEL 5
A00297:158:HT275DSXX:2:2535:6027:35822 chr5 58564437 N chr5 58564862 N DEL 5
A00297:158:HT275DSXX:3:2107:8079:13761 chr9 66249826 N chr9 66249900 N DUP 27
A00404:156:HV37TDSXX:3:1178:3875:17284 chr9 66249792 N chr9 66249843 N DEL 19
A00297:158:HT275DSXX:4:1116:10782:16783 chr9 66249722 N chr9 66249900 N DUP 10
A00297:158:HT275DSXX:4:1116:8513:14638 chr9 66249722 N chr9 66249900 N DUP 10
A00297:158:HT275DSXX:3:1422:25635:2769 chr4 176723651 N chr4 176723721 N DEL 5
A00404:155:HV27LDSXX:4:1348:29161:10160 chr4 176723568 N chr4 176723656 N DUP 5
A00404:155:HV27LDSXX:1:2175:8314:3583 chr4 176723568 N chr4 176723656 N DUP 5
A00404:156:HV37TDSXX:4:2518:26377:27539 chr4 176723568 N chr4 176723656 N DUP 5
A00297:158:HT275DSXX:1:1450:10194:35556 chr4 176723568 N chr4 176723656 N DUP 5
A00404:156:HV37TDSXX:3:2443:29939:17957 chr20 16035196 N chr20 16035263 N DEL 5
A00404:156:HV37TDSXX:3:2443:30038:17973 chr20 16035196 N chr20 16035263 N DEL 5
A00297:158:HT275DSXX:4:1416:29170:32095 chr20 16035246 N chr20 16035315 N DUP 11
A00404:155:HV27LDSXX:3:1117:32217:11130 chr20 16035246 N chr20 16035315 N DUP 15
A00404:156:HV37TDSXX:2:2331:14000:15843 chr20 16035224 N chr20 16035279 N DUP 17
A00404:155:HV27LDSXX:1:2468:20428:19554 chr20 16035273 N chr20 16035347 N DEL 20
A00297:158:HT275DSXX:1:2345:12518:1971 chr20 16035273 N chr20 16035347 N DEL 19
A00404:156:HV37TDSXX:2:1607:30147:30154 chr20 16035273 N chr20 16035347 N DEL 16
A00297:158:HT275DSXX:1:1239:10963:31281 chr20 16035275 N chr20 16035349 N DEL 12
A00404:155:HV27LDSXX:3:1641:24126:18818 chr20 16035274 N chr20 16035348 N DEL 13
A00404:156:HV37TDSXX:2:2107:28438:32581 chr20 16035278 N chr20 16035352 N DEL 10
A00404:155:HV27LDSXX:1:2102:28583:12665 chr20 16035278 N chr20 16035352 N DEL 10
A00404:156:HV37TDSXX:4:2361:4282:9659 chr20 48664890 N chr20 48665169 N DEL 5
A00404:155:HV27LDSXX:2:2111:2772:7701 chr20 48665051 N chr20 48665274 N DEL 4
A00297:158:HT275DSXX:3:1253:26467:3020 chr20 48664968 N chr20 48665026 N DEL 6
A00297:158:HT275DSXX:4:2149:13449:9157 chr20 48664968 N chr20 48665026 N DEL 6
A00404:156:HV37TDSXX:3:1252:4752:4742 chr20 48664968 N chr20 48665026 N DEL 6
A00404:155:HV27LDSXX:3:1534:31819:9721 chr20 48665079 N chr20 48665134 N DUP 9
A00404:156:HV37TDSXX:2:1170:22182:25755 chr20 48664888 N chr20 48665165 N DUP 5
A00404:156:HV37TDSXX:3:2563:30798:36135 chr20 48665069 N chr20 48665320 N DEL 5
A00404:155:HV27LDSXX:3:1422:27606:33771 chr20 48664914 N chr20 48665412 N DUP 4
A00297:158:HT275DSXX:1:2162:31150:14418 chr20 48664914 N chr20 48665412 N DUP 9
A00297:158:HT275DSXX:1:2162:31358:13620 chr20 48664914 N chr20 48665412 N DUP 9
A00404:156:HV37TDSXX:4:1517:1380:18693 chr20 48665412 N chr20 48665469 N DEL 20
A00404:155:HV27LDSXX:3:1668:9769:10895 chr20 48664914 N chr20 48665412 N DUP 10
A00404:155:HV27LDSXX:3:2667:7455:26929 chr20 48664914 N chr20 48665412 N DUP 10
A00404:155:HV27LDSXX:3:2668:3188:2754 chr20 48664914 N chr20 48665412 N DUP 10
A00404:156:HV37TDSXX:3:2113:27407:4523 chr20 48664914 N chr20 48665412 N DUP 5
A00297:158:HT275DSXX:2:2315:11993:3693 chr20 48664968 N chr20 48665468 N DEL 10
A00404:155:HV27LDSXX:2:1660:8522:19883 chr20 48664968 N chr20 48665468 N DEL 10
A00404:155:HV27LDSXX:2:1660:8540:19914 chr20 48664968 N chr20 48665468 N DEL 10
A00297:158:HT275DSXX:4:2405:17056:34820 chr3 95588253 N chr3 95588412 N DUP 10
A00297:158:HT275DSXX:3:1623:12952:31469 chr3 95588288 N chr3 95588449 N DEL 5
A00404:155:HV27LDSXX:3:2128:17571:29387 chr3 95588288 N chr3 95588449 N DEL 5
A00404:156:HV37TDSXX:3:1166:30761:35509 chr3 95588288 N chr3 95588449 N DEL 5
A00404:156:HV37TDSXX:2:2654:9353:33661 chr3 95588286 N chr3 95588447 N DEL 10
A00404:155:HV27LDSXX:4:2230:28203:2769 chr3 95588286 N chr3 95588447 N DEL 10
A00404:155:HV27LDSXX:2:2340:9968:28839 chr20 47951398 N chr20 47951478 N DEL 20
A00297:158:HT275DSXX:2:2233:9182:10379 chr20 47951398 N chr20 47951478 N DEL 22
A00404:155:HV27LDSXX:4:2508:25192:24862 chr20 47951398 N chr20 47951478 N DEL 15
A00297:158:HT275DSXX:2:2226:16098:21042 chr20 47951398 N chr20 47951478 N DEL 15
A00297:158:HT275DSXX:1:2660:17960:13307 chr20 47951398 N chr20 47951478 N DEL 16
A00297:158:HT275DSXX:1:2660:17978:13338 chr20 47951398 N chr20 47951478 N DEL 16
A00297:158:HT275DSXX:3:1549:14606:8249 chr20 47951469 N chr20 47951557 N DEL 2
A00404:156:HV37TDSXX:3:1611:23737:28228 chr20 47951398 N chr20 47951478 N DEL 12
A00297:158:HT275DSXX:3:2560:32380:16454 chr20 47951398 N chr20 47951478 N DEL 17
A00297:158:HT275DSXX:3:1540:1814:35352 chr20 47951398 N chr20 47951478 N DEL 17
A00297:158:HT275DSXX:2:2367:14705:26897 chr20 47951398 N chr20 47951478 N DEL 17
A00404:156:HV37TDSXX:4:2678:28664:3255 chr20 47951398 N chr20 47951478 N DEL 17
A00297:158:HT275DSXX:3:1635:18846:22827 chr20 47951312 N chr20 47951549 N DUP 5
A00297:158:HT275DSXX:2:1564:12653:33082 chr20 47951398 N chr20 47951478 N DEL 17
A00404:155:HV27LDSXX:1:2166:24587:7874 chr20 47951398 N chr20 47951478 N DEL 17
A00404:156:HV37TDSXX:4:2372:4607:23813 chr20 47951398 N chr20 47951478 N DEL 17
A00297:158:HT275DSXX:2:1321:32353:5916 chr20 47951401 N chr20 47951481 N DEL 10
A00404:155:HV27LDSXX:4:1225:29179:25097 chr20 47951407 N chr20 47951487 N DEL 7
A00404:155:HV27LDSXX:4:2121:24668:17722 chr20 47951535 N chr20 47951621 N DUP 5
A00404:155:HV27LDSXX:2:2678:10031:8187 chr20 47951407 N chr20 47951487 N DEL 6
A00404:155:HV27LDSXX:1:2366:12970:18349 chr20 47951410 N chr20 47951490 N DEL 3
A00404:155:HV27LDSXX:2:2158:27769:26224 chr20 47951535 N chr20 47951621 N DUP 5
A00297:158:HT275DSXX:3:1621:9534:6042 chr20 47951301 N chr20 47951504 N DEL 5
A00297:158:HT275DSXX:3:1549:14606:8249 chr20 47951535 N chr20 47951621 N DUP 5
A00297:158:HT275DSXX:2:2158:25229:21418 chr20 47951535 N chr20 47951621 N DUP 5
A00297:158:HT275DSXX:2:1352:1244:21245 chr20 47951535 N chr20 47951621 N DUP 5
A00404:156:HV37TDSXX:1:2526:18629:32910 chr20 47951535 N chr20 47951621 N DUP 5
A00404:155:HV27LDSXX:3:1461:17960:10708 chr20 47951210 N chr20 47951535 N DEL 5
A00297:158:HT275DSXX:2:1510:10339:16047 chr20 47951210 N chr20 47951535 N DEL 5
A00404:155:HV27LDSXX:4:1310:11767:12446 chr20 47951248 N chr20 47951539 N DEL 5
A00404:155:HV27LDSXX:4:2507:11577:25488 chr13 79801321 N chr13 79801382 N DUP 5
A00297:158:HT275DSXX:4:1564:29550:16595 chr13 79801321 N chr13 79801382 N DUP 5
A00404:155:HV27LDSXX:4:1675:8865:27586 chr13 79801321 N chr13 79801382 N DUP 5
A00404:156:HV37TDSXX:4:2433:26639:20509 chr13 79801337 N chr13 79801400 N DEL 5
A00404:156:HV37TDSXX:4:2433:26793:20650 chr13 79801337 N chr13 79801400 N DEL 5
A00297:158:HT275DSXX:1:1173:11785:1736 chr13 79801380 N chr13 79801441 N DEL 5
A00404:155:HV27LDSXX:3:2156:32289:27853 chr10 116728152 N chr10 116728284 N DUP 5
A00297:158:HT275DSXX:4:1466:11749:32769 chr10 116728156 N chr10 116728290 N DEL 5
A00297:158:HT275DSXX:1:2530:16423:36292 chr10 116728166 N chr10 116728300 N DEL 1
A00404:155:HV27LDSXX:4:2372:4607:24878 chr2 142906155 N chr2 142906206 N DUP 7
A00404:155:HV27LDSXX:2:2221:30074:34663 chr12 74951594 N chr12 74951734 N DEL 4
A00404:155:HV27LDSXX:4:2177:5132:36652 chr12 74951594 N chr12 74951734 N DEL 4
A00404:155:HV27LDSXX:4:2177:5692:36620 chr12 74951594 N chr12 74951734 N DEL 4
A00404:156:HV37TDSXX:2:2609:20934:10723 chr12 74951594 N chr12 74951734 N DEL 5
A00404:156:HV37TDSXX:4:1338:7428:25128 chr12 74951594 N chr12 74951734 N DEL 7
A00404:156:HV37TDSXX:3:1522:4580:26616 chr12 74951594 N chr12 74951734 N DEL 7
A00404:155:HV27LDSXX:3:2334:17273:23484 chr12 74951594 N chr12 74951734 N DEL 7
A00404:155:HV27LDSXX:1:2355:29948:12399 chr12 74951621 N chr12 74951670 N DUP 5
A00404:155:HV27LDSXX:4:1454:14425:31986 chr12 74951650 N chr12 74951724 N DEL 20
A00297:158:HT275DSXX:3:1540:20790:6684 chr12 74951625 N chr12 74951724 N DEL 17
A00297:158:HT275DSXX:3:2539:19479:25426 chr12 74951625 N chr12 74951724 N DEL 17
A00297:158:HT275DSXX:2:2141:12843:8860 chr12 74951627 N chr12 74951726 N DEL 13
A00404:156:HV37TDSXX:2:2271:11369:2801 chr12 74951622 N chr12 74951770 N DEL 8
A00404:156:HV37TDSXX:4:2210:7455:15280 chr7 13102575 N chr7 13103052 N DEL 5
A00404:155:HV27LDSXX:1:1207:12038:14105 chr7 13102575 N chr7 13103052 N DEL 5
A00404:155:HV27LDSXX:1:1513:9055:12915 chr7 13102552 N chr7 13102629 N DEL 5
A00404:155:HV27LDSXX:3:1338:3432:25504 chr7 13102653 N chr7 13102770 N DEL 14
A00404:156:HV37TDSXX:3:1407:20717:12571 chr4 142246067 N chr4 142246126 N DEL 25
A00404:156:HV37TDSXX:3:2126:9191:1564 chr4 142246067 N chr4 142246126 N DEL 25
A00297:158:HT275DSXX:3:2517:27398:7482 chr4 142246067 N chr4 142246126 N DEL 25
A00404:155:HV27LDSXX:4:1453:27208:12915 chr4 142246067 N chr4 142246126 N DEL 25
A00297:158:HT275DSXX:1:2277:32624:12680 chr4 142246067 N chr4 142246126 N DEL 22
A00404:156:HV37TDSXX:1:2321:25211:13714 chr4 142246078 N chr4 142246137 N DEL 22
A00404:156:HV37TDSXX:4:1125:13982:28933 chr4 142246067 N chr4 142246126 N DEL 21
A00297:158:HT275DSXX:2:1205:18511:22623 chr4 142246029 N chr4 142246126 N DEL 15
A00404:155:HV27LDSXX:4:1453:2537:3787 chr4 142246036 N chr4 142246133 N DEL 8
A00297:158:HT275DSXX:1:1647:5945:10661 chrX 113299937 N chrX 113300115 N DEL 11
A00404:155:HV27LDSXX:1:2529:7003:4194 chrX 113299937 N chrX 113300115 N DEL 12
A00404:155:HV27LDSXX:4:1307:20482:6558 chr19 689258 N chr19 689335 N DUP 18
A00404:155:HV27LDSXX:3:1358:8775:22075 chr19 689277 N chr19 689423 N DUP 5
A00297:158:HT275DSXX:1:1174:26775:29731 chr19 689354 N chr19 689422 N DUP 25
A00404:156:HV37TDSXX:1:1352:5204:33990 chr19 689354 N chr19 689422 N DUP 25
A00404:156:HV37TDSXX:2:1612:6388:22858 chr19 689354 N chr19 689422 N DUP 25
A00404:156:HV37TDSXX:4:2273:30879:15233 chr19 689302 N chr19 689372 N DEL 33
A00404:156:HV37TDSXX:3:1378:4227:21089 chr19 689302 N chr19 689372 N DEL 33
A00404:156:HV37TDSXX:4:1611:4029:10567 chr19 689302 N chr19 689372 N DEL 33
A00404:156:HV37TDSXX:1:1317:30680:9533 chr19 689302 N chr19 689372 N DEL 29
A00297:158:HT275DSXX:2:2245:11252:20478 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:4:2601:2935:26303 chr16 46397308 N chr16 46397477 N DUP 5
A00404:156:HV37TDSXX:1:2154:26467:6026 chr16 46397235 N chr16 46397301 N DEL 5
A00297:158:HT275DSXX:4:2523:2908:2143 chr16 46397195 N chr16 46397380 N DUP 1
A00297:158:HT275DSXX:1:1243:5791:30874 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:2:1256:25807:13244 chr16 46397317 N chr16 46397486 N DUP 5
A00297:158:HT275DSXX:3:2363:29306:15796 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:1:2305:10113:21261 chr16 46397237 N chr16 46397471 N DUP 7
A00404:155:HV27LDSXX:1:1550:16477:5447 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:3:2404:25681:19194 chr16 46397195 N chr16 46397380 N DUP 1
A00297:158:HT275DSXX:1:2131:27941:28839 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:4:2220:1895:23218 chr16 46397195 N chr16 46397380 N DUP 1
A00297:158:HT275DSXX:3:2317:5159:14403 chr16 46397369 N chr16 46397440 N DUP 4
A00297:158:HT275DSXX:2:2129:10203:25582 chr16 46397195 N chr16 46397380 N DUP 1
A00297:158:HT275DSXX:4:1365:3540:27007 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:2:2170:10538:11068 chr16 46397195 N chr16 46397380 N DUP 1
A00404:155:HV27LDSXX:4:2575:9887:28103 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:2:1140:7084:7999 chr16 46397313 N chr16 46397482 N DUP 5
A00404:156:HV37TDSXX:2:2214:4716:24095 chr16 46397195 N chr16 46397380 N DUP 1
A00404:155:HV27LDSXX:1:2614:10484:13416 chr16 46397369 N chr16 46397440 N DUP 3
A00297:158:HT275DSXX:1:2365:31530:8656 chr16 46397195 N chr16 46397380 N DUP 1
A00297:158:HT275DSXX:4:2228:1461:19366 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:4:2251:7961:25457 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:1:1170:29894:22294 chr16 46397195 N chr16 46397380 N DUP 1
A00297:158:HT275DSXX:2:1571:19732:30342 chr16 46397342 N chr16 46397488 N DUP 3
A00404:155:HV27LDSXX:1:1609:18069:26960 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:4:2343:2465:15906 chr16 46397195 N chr16 46397380 N DUP 1
A00404:155:HV27LDSXX:3:2178:27995:2503 chr16 46397195 N chr16 46397380 N DUP 1
A00404:156:HV37TDSXX:3:1303:3251:15890 chr16 46397195 N chr16 46397380 N DUP 1
A00404:155:HV27LDSXX:3:1633:27353:17675 chr16 13126949 N chr16 13127050 N DUP 1
A00404:156:HV37TDSXX:1:1451:14109:7388 chr4 147798892 N chr4 147798943 N DEL 17
A00404:156:HV37TDSXX:3:1304:6940:19022 chr22 40687187 N chr22 40687350 N DEL 15
A00404:156:HV37TDSXX:1:1524:6994:28635 chr1 41425549 N chr1 41425820 N DUP 6
A00297:158:HT275DSXX:2:1611:32253:10629 chr1 41425546 N chr1 41425817 N DUP 9
A00297:158:HT275DSXX:3:2337:6732:9424 chr1 41425549 N chr1 41425820 N DUP 6
A00404:156:HV37TDSXX:1:1448:7997:20635 chr4 1537252 N chr4 1537311 N DEL 4
A00404:155:HV27LDSXX:2:1643:14217:10958 chr22 39563908 N chr22 39564019 N DEL 9
A00404:155:HV27LDSXX:3:2361:32434:11851 chr22 39563908 N chr22 39564019 N DEL 9
A00404:155:HV27LDSXX:4:2261:19831:13542 chr22 39563865 N chr22 39564019 N DEL 9
A00404:155:HV27LDSXX:2:1543:14877:17738 chr22 39563865 N chr22 39564019 N DEL 9
A00404:155:HV27LDSXX:1:2644:17806:31986 chr22 39563909 N chr22 39564020 N DEL 9
A00404:156:HV37TDSXX:1:1610:26530:35039 chr22 39563911 N chr22 39564022 N DEL 9
A00297:158:HT275DSXX:1:1219:8205:32675 chr1 86215760 N chr1 86215957 N DEL 3
A00297:158:HT275DSXX:2:1620:18141:27242 chr1 86215733 N chr1 86215927 N DEL 5
A00404:155:HV27LDSXX:2:1217:27290:31970 chr6 32595661 N chr6 32595758 N DUP 5
A00404:156:HV37TDSXX:1:1638:20835:4319 chr6 32595653 N chr6 32595751 N DUP 5
A00404:155:HV27LDSXX:4:1137:12509:14325 chr6 32595666 N chr6 32596167 N DUP 6
A00404:156:HV37TDSXX:3:2266:2546:11193 chr6 32595631 N chr6 32595728 N DUP 11
A00404:156:HV37TDSXX:3:2266:2844:11209 chr6 32595631 N chr6 32595728 N DUP 5
A00404:155:HV27LDSXX:4:1424:30373:32706 chr6 32595776 N chr6 32595902 N DUP 3
A00404:155:HV27LDSXX:1:2332:26521:35086 chr6 32595890 N chr6 32596069 N DEL 5
A00404:155:HV27LDSXX:4:2343:31259:8500 chr6 32595780 N chr6 32595906 N DUP 2
A00404:156:HV37TDSXX:1:2361:15709:22654 chr6 32595890 N chr6 32596118 N DEL 5
A00404:156:HV37TDSXX:1:2670:30436:35321 chr6 32595902 N chr6 32596130 N DEL 1
A00404:156:HV37TDSXX:4:2132:18792:36573 chr6 32595890 N chr6 32596069 N DEL 5
A00297:158:HT275DSXX:3:1253:13386:5290 chr6 32595890 N chr6 32596069 N DEL 5
A00404:155:HV27LDSXX:3:2667:24966:32550 chr6 32595890 N chr6 32596069 N DEL 5
A00297:158:HT275DSXX:2:2159:24316:29136 chr6 32595845 N chr6 32595971 N DUP 2
A00404:156:HV37TDSXX:2:2429:14886:5228 chr6 32595631 N chr6 32595905 N DUP 19
A00404:155:HV27LDSXX:2:1340:26811:18490 chr6 32595883 N chr6 32596009 N DUP 5
A00404:155:HV27LDSXX:2:1340:27001:18568 chr6 32595883 N chr6 32596009 N DUP 5
A00404:156:HV37TDSXX:2:2351:13150:8735 chr6 32595883 N chr6 32596009 N DUP 5
A00404:155:HV27LDSXX:4:1606:32624:3568 chr17 1247476 N chr17 1247593 N DEL 12
A00297:158:HT275DSXX:2:2159:26133:7795 chr1 3471001 N chr1 3471124 N DEL 1
A00404:156:HV37TDSXX:1:1124:24089:3756 chr1 3471052 N chr1 3471171 N DEL 5
A00404:155:HV27LDSXX:1:2248:28131:16266 chr1 3471013 N chr1 3471226 N DEL 28
A00404:155:HV27LDSXX:1:2248:28131:16266 chr1 3470839 N chr1 3471231 N DEL 7
A00297:158:HT275DSXX:1:1330:30933:23719 chr1 3471025 N chr1 3471238 N DEL 3
A00404:155:HV27LDSXX:2:2555:6081:15937 chr15 70279783 N chr15 70279974 N DEL 2
A00404:155:HV27LDSXX:2:2555:7157:19398 chr15 70279783 N chr15 70279974 N DEL 2
A00404:156:HV37TDSXX:2:2437:25418:24345 chr15 70279785 N chr15 70279976 N DEL 5
A00404:155:HV27LDSXX:3:2509:5412:8202 chr15 70279790 N chr15 70280175 N DEL 19
A00404:156:HV37TDSXX:4:2202:28926:20619 chr15 70279813 N chr15 70280002 N DUP 5
A00404:156:HV37TDSXX:4:2473:4291:16752 chr15 70279813 N chr15 70280002 N DUP 5
A00404:156:HV37TDSXX:4:2473:4815:18255 chr15 70279813 N chr15 70280002 N DUP 5
A00404:155:HV27LDSXX:2:2217:19759:30483 chr15 70279813 N chr15 70280002 N DUP 5
A00404:155:HV27LDSXX:1:2213:26874:14810 chr15 70279815 N chr15 70280004 N DUP 5
A00297:158:HT275DSXX:3:2337:21802:36652 chr15 70279896 N chr15 70279961 N DEL 5
A00404:156:HV37TDSXX:1:1610:24478:8030 chr15 70279896 N chr15 70279961 N DEL 2
A00404:155:HV27LDSXX:3:1459:4508:1908 chr15 70279896 N chr15 70279961 N DEL 13
A00404:156:HV37TDSXX:3:2307:7862:17707 chr15 70279896 N chr15 70279961 N DEL 10
A00404:156:HV37TDSXX:4:1239:18683:27993 chr15 70279896 N chr15 70279961 N DEL 5
A00404:155:HV27LDSXX:3:1451:10899:28823 chr15 70279832 N chr15 70279961 N DEL 5
A00404:156:HV37TDSXX:4:1537:20455:12931 chr15 70279835 N chr15 70280158 N DEL 5
A00404:156:HV37TDSXX:4:1339:6225:7639 chr15 70279837 N chr15 70280160 N DEL 5
A00404:155:HV27LDSXX:3:1544:8305:32910 chr15 70279908 N chr15 70280167 N DEL 5
A00404:156:HV37TDSXX:3:2478:1714:4679 chr15 70280029 N chr15 70280158 N DEL 5
A00404:155:HV27LDSXX:2:1344:4200:19946 chr15 70280029 N chr15 70280158 N DEL 5
A00404:155:HV27LDSXX:2:2217:19759:30483 chr15 70280029 N chr15 70280158 N DEL 5
A00297:158:HT275DSXX:2:2219:6831:19930 chr15 70280029 N chr15 70280158 N DEL 5
A00404:155:HV27LDSXX:3:1528:9399:36965 chr15 70280029 N chr15 70280158 N DEL 5
A00404:155:HV27LDSXX:3:1529:9869:1485 chr15 70280029 N chr15 70280158 N DEL 5
A00297:158:HT275DSXX:1:2147:20772:20682 chr15 70280029 N chr15 70280158 N DEL 5
A00404:155:HV27LDSXX:2:2327:21558:8484 chr15 70280029 N chr15 70280158 N DEL 5
A00404:156:HV37TDSXX:2:1360:25545:32643 chr15 70279839 N chr15 70280158 N DEL 5
A00297:158:HT275DSXX:2:1669:4426:25160 chr15 70279848 N chr15 70280169 N DEL 4
A00297:158:HT275DSXX:4:1216:14082:14011 chr15 70280029 N chr15 70280158 N DEL 8
A00404:156:HV37TDSXX:2:1324:19533:32690 chr15 70280029 N chr15 70280158 N DEL 7
A00297:158:HT275DSXX:3:2633:12120:7795 chr15 70280029 N chr15 70280158 N DEL 5
A00404:156:HV37TDSXX:2:1232:29577:21840 chr15 70280029 N chr15 70280158 N DEL 5
A00404:156:HV37TDSXX:1:1610:24641:7999 chr15 70279904 N chr15 70280425 N DEL 18
A00297:158:HT275DSXX:2:2211:11749:24283 chr14 105622612 N chr14 105622671 N DEL 8
A00297:158:HT275DSXX:4:2413:24089:13870 chr18 69894594 N chr18 69894686 N DEL 7
A00404:155:HV27LDSXX:4:1375:22833:28855 chr18 69894671 N chr18 69894796 N DEL 2
A00404:156:HV37TDSXX:3:1518:21187:31328 chr20 60500528 N chr20 60500885 N DEL 6
A00297:158:HT275DSXX:1:2622:30662:15264 chr20 60500888 N chr20 60501258 N DEL 9
A00297:158:HT275DSXX:1:1635:10673:12148 chr20 60500896 N chr20 60501354 N DEL 6
A00404:155:HV27LDSXX:1:1305:32362:17206 chr20 60500659 N chr20 60501002 N DUP 5
A00404:155:HV27LDSXX:2:1505:22101:28119 chr20 60500619 N chr20 60500977 N DEL 11
A00404:156:HV37TDSXX:2:2547:28980:8688 chr20 60500860 N chr20 60501053 N DUP 1
A00404:156:HV37TDSXX:3:1451:25753:20008 chr20 60500664 N chr20 60501028 N DEL 5
A00297:158:HT275DSXX:4:1457:19949:16971 chr20 60500814 N chr20 60501159 N DEL 1
A00404:155:HV27LDSXX:1:2168:25563:25441 chr20 60500428 N chr20 60501335 N DEL 5
A00404:155:HV27LDSXX:1:2522:11993:27179 chr20 60501428 N chr20 60501655 N DEL 5
A00404:155:HV27LDSXX:3:1121:2582:15452 chr20 60501302 N chr20 60501749 N DUP 5
A00404:155:HV27LDSXX:3:1630:23891:18129 chr2 231955018 N chr2 231955089 N DEL 4
A00404:155:HV27LDSXX:3:1630:24334:18427 chr2 231955018 N chr2 231955089 N DEL 4
A00404:156:HV37TDSXX:1:1359:12346:12101 chr2 231955048 N chr2 231955121 N DUP 5
A00404:156:HV37TDSXX:1:1426:24126:13025 chr2 231955053 N chr2 231955126 N DUP 5
A00404:155:HV27LDSXX:2:2350:16342:22498 chr4 2210771 N chr4 2211450 N DUP 5
A00297:158:HT275DSXX:4:1349:27814:22263 chr22 16254710 N chr22 16254891 N DUP 1
A00297:158:HT275DSXX:2:1666:18810:9330 chr8 62870817 N chr8 62870870 N DEL 1
A00404:156:HV37TDSXX:1:1635:16233:12759 chrY 13380148 N chrY 13380221 N DEL 5
A00297:158:HT275DSXX:4:2118:21721:18568 chr3 139802762 N chr3 139802845 N DUP 5
A00404:156:HV37TDSXX:4:2604:26323:21966 chr3 139802762 N chr3 139802845 N DUP 5
A00404:156:HV37TDSXX:1:2540:16405:31469 chr3 154136361 N chr3 154136428 N DUP 8
A00297:158:HT275DSXX:3:2420:7202:34882 chr3 154136361 N chr3 154136428 N DUP 9
A00297:158:HT275DSXX:1:1432:9977:35744 chr14 105083412 N chr14 105083564 N DEL 28
A00404:155:HV27LDSXX:3:1526:3396:34460 chr14 105083379 N chr14 105083682 N DEL 5
A00404:156:HV37TDSXX:3:1245:30472:4883 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:4:1316:28122:17691 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:2319:13720:3302 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:1:1431:3775:31735 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:3:1162:17336:3709 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:3:2371:17879:1485 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:1:2242:31756:13182 chr2 32866889 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:1:2567:29948:7889 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:4:1570:5927:2268 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:4:1410:6063:3411 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:2:1569:24596:20635 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:2576:13286:35399 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:1:2528:18584:25974 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:1:2543:15302:33317 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:1174:8757:19163 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:1:1225:20509:19006 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:1:1338:14678:25598 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:4:1639:20392:14857 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:4:2413:22625:22451 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:1:1323:30101:22686 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:4:1368:21450:36573 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:3:1231:5511:23625 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:4:1207:29324:30138 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:2:2560:14244:7341 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:4:1414:15501:8641 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:1:2415:16432:16579 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:4:2455:4101:17769 chr2 32866896 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:1:2305:7473:12649 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:2:2276:29749:12806 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:1:1174:9317:27868 chr2 32866892 N chr2 32867280 N DEL 1
A00404:155:HV27LDSXX:4:2144:18484:26772 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:2:1251:25238:30796 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:4:1165:3161:13636 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:1:1648:14787:30702 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:2:2608:11975:16125 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:4:2662:24297:2018 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:2:1445:29731:11992 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:2:1465:9100:29966 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:1:2509:21468:24424 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:1328:21739:4820 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:1606:29586:34006 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:1:1321:11568:22060 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:3:1272:18991:5697 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:2:2102:26160:10441 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:3:1451:6632:23531 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:2:2424:1434:32221 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:4:2247:6777:1642 chr2 32866897 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:4:1677:28293:2801 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:1:1170:5204:11945 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:3:2172:14344:12273 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:2:1473:20528:29496 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:3:1448:15329:2080 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:2:1157:2926:2206 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:4:1354:11785:9064 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:1:1154:28628:20729 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:1:2443:30282:33051 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:1:1353:2230:18568 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:1510:23194:35055 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:1628:2962:24972 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:2:2135:29857:28808 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:4:1414:7554:1705 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:1377:31548:20400 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:2:2566:12237:23907 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:4:1425:3676:2065 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:4:1616:7862:35963 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:3:2602:7798:34632 chr2 32866894 N chr2 32867280 N DEL 2
A00297:158:HT275DSXX:3:1678:31991:24706 chr2 32866894 N chr2 32867280 N DEL 2
A00404:155:HV27LDSXX:3:1665:9308:18427 chr2 32866894 N chr2 32867280 N DEL 2
A00404:156:HV37TDSXX:2:2615:30138:14700 chr3 42798006 N chr3 42798102 N DUP 5
A00404:156:HV37TDSXX:2:2313:22797:3583 chr1 73390675 N chr1 73390799 N DEL 10
A00404:155:HV27LDSXX:4:1536:10511:7701 chr11 468887 N chr11 469321 N DEL 27
A00404:156:HV37TDSXX:2:1133:16920:5869 chr11 469021 N chr11 469299 N DEL 36
A00404:156:HV37TDSXX:4:2277:29405:27680 chr11 468961 N chr11 469572 N DUP 5
A00404:156:HV37TDSXX:4:2574:31873:34773 chr11 468990 N chr11 469578 N DUP 5
A00404:156:HV37TDSXX:2:2575:24297:7780 chr11 469032 N chr11 469216 N DUP 2
A00297:158:HT275DSXX:3:2256:26964:20102 chr11 469113 N chr11 469208 N DUP 5
A00297:158:HT275DSXX:4:1654:12717:33160 chr11 469444 N chr11 469553 N DEL 4
A00297:158:HT275DSXX:1:1674:3558:22936 chr11 469444 N chr11 469553 N DEL 19
A00297:158:HT275DSXX:2:2444:4679:2300 chr11 469444 N chr11 469553 N DEL 19
A00404:156:HV37TDSXX:4:1116:19027:21292 chr11 469444 N chr11 469553 N DEL 19
A00404:155:HV27LDSXX:3:2530:14922:24893 chr11 469444 N chr11 469553 N DEL 23
A00404:156:HV37TDSXX:2:1521:24062:20400 chr11 469444 N chr11 469553 N DEL 24
A00297:158:HT275DSXX:3:1345:26865:35556 chr11 469444 N chr11 469553 N DEL 22
A00404:156:HV37TDSXX:4:2201:22399:17550 chr11 469444 N chr11 469553 N DEL 22
A00404:156:HV37TDSXX:2:2675:17065:35900 chrX 147152544 N chrX 147152603 N DEL 9
A00404:155:HV27LDSXX:2:2559:12201:13072 chrX 147152502 N chrX 147152579 N DUP 36
A00404:155:HV27LDSXX:3:1446:12264:24392 chrX 147152530 N chrX 147152587 N DUP 29
A00404:155:HV27LDSXX:1:1537:27507:11052 chrX 147152503 N chrX 147152554 N DEL 5
A00404:155:HV27LDSXX:4:2276:3549:22921 chrX 147152504 N chrX 147152555 N DEL 5
A00404:156:HV37TDSXX:3:2359:11017:14309 chrX 147152493 N chrX 147152562 N DEL 5
A00404:155:HV27LDSXX:2:2351:28772:6668 chr6 15415817 N chr6 15415943 N DUP 5
A00404:156:HV37TDSXX:1:1515:4164:23735 chr6 15415817 N chr6 15415943 N DUP 5
A00404:156:HV37TDSXX:3:1624:4029:13510 chr6 15415817 N chr6 15415943 N DUP 5
A00404:155:HV27LDSXX:3:1675:4661:10160 chr6 15415817 N chr6 15415943 N DUP 5
A00404:156:HV37TDSXX:2:2274:18864:11240 chr6 15415801 N chr6 15415984 N DUP 12
A00404:155:HV27LDSXX:3:1110:3830:2080 chr6 15415955 N chr6 15416088 N DUP 5
A00297:158:HT275DSXX:2:1272:31801:2863 chr6 15415833 N chr6 15415961 N DEL 5
A00404:155:HV27LDSXX:3:1563:19506:8249 chr6 15415857 N chr6 15415977 N DEL 21
A00404:156:HV37TDSXX:4:1232:12129:4523 chr6 15415847 N chr6 15415974 N DEL 7
A00297:158:HT275DSXX:2:2435:14859:3302 chr6 15415857 N chr6 15415977 N DEL 21
A00404:155:HV27LDSXX:3:2425:8540:34695 chr6 15415832 N chr6 15416009 N DEL 10
A00404:156:HV37TDSXX:4:2101:2971:15655 chr6 15415813 N chr6 15416036 N DEL 1
A00297:158:HT275DSXX:2:1636:20826:23782 chr6 15415802 N chr6 15416025 N DEL 7
A00297:158:HT275DSXX:1:2338:4237:32941 chr1 195841338 N chr1 195841393 N DEL 7
A00404:156:HV37TDSXX:2:1349:26485:5995 chr1 195841338 N chr1 195841393 N DEL 11
A00404:156:HV37TDSXX:2:1534:6216:35368 chr4 706309 N chr4 706908 N DEL 5
A00404:155:HV27LDSXX:3:2630:16902:23531 chr4 706347 N chr4 707152 N DEL 5
A00404:156:HV37TDSXX:2:2401:18530:24878 chr4 706386 N chr4 706488 N DEL 5
A00404:155:HV27LDSXX:3:1668:31665:36699 chr4 706386 N chr4 706488 N DEL 5
A00404:156:HV37TDSXX:4:2668:26549:35603 chr4 706386 N chr4 706488 N DEL 5
A00404:156:HV37TDSXX:4:2668:26612:34898 chr4 706386 N chr4 706488 N DEL 5
A00404:156:HV37TDSXX:3:1401:31593:19977 chr4 706386 N chr4 706488 N DEL 5
A00297:158:HT275DSXX:4:2153:25319:8140 chr4 706390 N chr4 706525 N DEL 5
A00404:156:HV37TDSXX:2:1641:26820:1908 chr4 706390 N chr4 706525 N DEL 5
A00404:156:HV37TDSXX:2:1641:27751:4147 chr4 706390 N chr4 706525 N DEL 5
A00404:156:HV37TDSXX:3:2455:12084:2691 chr4 706390 N chr4 706525 N DEL 5
A00297:158:HT275DSXX:1:1464:26404:23954 chr4 706390 N chr4 706525 N DEL 5
A00404:155:HV27LDSXX:4:1517:2645:31939 chr4 706390 N chr4 706525 N DEL 5
A00404:155:HV27LDSXX:1:2114:10592:13855 chr4 706390 N chr4 706525 N DEL 5
A00297:158:HT275DSXX:1:2417:3748:34538 chr4 706390 N chr4 706525 N DEL 5
A00404:156:HV37TDSXX:4:1173:30789:20494 chr4 706390 N chr4 706525 N DEL 5
A00404:156:HV37TDSXX:1:2573:3441:18881 chr4 706390 N chr4 706525 N DEL 5
A00404:156:HV37TDSXX:3:1676:27145:29590 chr4 706396 N chr4 706501 N DUP 14
A00404:155:HV27LDSXX:4:1125:20754:18333 chr4 706481 N chr4 706614 N DUP 5
A00404:156:HV37TDSXX:4:1133:10149:31219 chr4 706637 N chr4 706808 N DEL 20
A00404:155:HV27LDSXX:2:2328:3775:33207 chr4 706266 N chr4 706727 N DUP 5
A00404:155:HV27LDSXX:4:2442:22309:12571 chr4 706750 N chr4 707127 N DEL 2
A00404:156:HV37TDSXX:4:1133:10149:31219 chr4 706637 N chr4 706808 N DEL 10
A00404:155:HV27LDSXX:4:1442:22173:33755 chr4 706699 N chr4 707075 N DEL 5
A00404:156:HV37TDSXX:3:1664:4417:9392 chr4 1452910 N chr4 1453085 N DUP 10
A00404:155:HV27LDSXX:4:2641:21576:30530 chr4 1452908 N chr4 1453432 N DUP 12
A00404:155:HV27LDSXX:3:1574:27570:1329 chr4 1453164 N chr4 1453282 N DUP 5
A00404:156:HV37TDSXX:4:1242:15031:35916 chr10 3290924 N chr10 3291044 N DEL 5
A00404:155:HV27LDSXX:3:2359:11234:32784 chr10 3290895 N chr10 3290945 N DUP 5
A00297:158:HT275DSXX:4:2351:14705:17315 chr10 3290914 N chr10 3291034 N DEL 5
A00297:158:HT275DSXX:1:2249:17662:32017 chr22 44640086 N chr22 44640198 N DEL 7
A00297:158:HT275DSXX:1:2249:18710:30138 chr22 44640086 N chr22 44640198 N DEL 7
A00297:158:HT275DSXX:1:2249:17662:32017 chr22 44640094 N chr22 44640317 N DEL 15
A00404:156:HV37TDSXX:3:2211:22652:26349 chr22 44640119 N chr22 44640342 N DEL 17
A00404:156:HV37TDSXX:2:2223:30110:26522 chr22 44640139 N chr22 44640325 N DEL 35
A00404:156:HV37TDSXX:2:2223:30246:26349 chr22 44640126 N chr22 44640312 N DEL 40
A00404:156:HV37TDSXX:2:2618:24831:3568 chr22 44640089 N chr22 44640236 N DUP 5
A00297:158:HT275DSXX:1:2628:23194:7153 chr22 44640207 N chr22 44640319 N DEL 5
A00404:155:HV27LDSXX:3:2477:15863:17566 chr22 44640255 N chr22 44640404 N DEL 40
A00404:156:HV37TDSXX:1:1410:1967:23249 chr22 44640328 N chr22 44640403 N DEL 20
A00404:156:HV37TDSXX:3:2211:22652:26349 chr22 44640125 N chr22 44640348 N DEL 8
A00297:158:HT275DSXX:1:1315:18150:9909 chr22 44640218 N chr22 44640404 N DEL 10
A00297:158:HT275DSXX:2:1656:30083:20619 chr11 72268719 N chr11 72268784 N DUP 8
A00297:158:HT275DSXX:1:2556:22272:8625 chr11 72268784 N chr11 72268848 N DEL 8
A00404:155:HV27LDSXX:4:1171:31611:8735 chr11 72268704 N chr11 72268856 N DEL 4
A00404:156:HV37TDSXX:4:1353:28574:7388 chr11 72268995 N chr11 72269116 N DEL 11
A00297:158:HT275DSXX:1:2605:32298:22764 chr11 72268995 N chr11 72269116 N DEL 11
A00404:156:HV37TDSXX:2:2631:2537:18161 chr11 72268970 N chr11 72269116 N DEL 11
A00404:156:HV37TDSXX:4:2658:5565:1736 chr11 72268970 N chr11 72269116 N DEL 11
A00404:156:HV37TDSXX:2:1436:17038:33379 chr2 241572900 N chr2 241573306 N DEL 11
A00297:158:HT275DSXX:1:2171:23791:15295 chr2 241572884 N chr2 241573169 N DEL 6
A00297:158:HT275DSXX:1:2171:23791:15295 chr2 241572884 N chr2 241573169 N DEL 6
A00404:156:HV37TDSXX:2:1157:27127:26897 chr2 241572933 N chr2 241573055 N DEL 5
A00297:158:HT275DSXX:2:1436:19596:4523 chr2 241572899 N chr2 241573020 N DUP 5
A00404:156:HV37TDSXX:4:2266:27769:17519 chr2 241572997 N chr2 241573319 N DUP 5
A00404:156:HV37TDSXX:4:2266:27769:17519 chr2 241572996 N chr2 241573199 N DEL 9
A00297:158:HT275DSXX:1:2340:19370:15468 chr2 241573015 N chr2 241573178 N DEL 5
A00404:156:HV37TDSXX:2:1137:32542:34679 chr2 241573024 N chr2 241573187 N DEL 5
A00297:158:HT275DSXX:4:2639:21811:29590 chr2 241572933 N chr2 241573178 N DEL 5
A00404:155:HV27LDSXX:3:2551:23149:5948 chr2 241572919 N chr2 241573040 N DUP 5
A00404:155:HV27LDSXX:2:2651:2121:35853 chr2 241573007 N chr2 241573127 N DUP 2
A00404:156:HV37TDSXX:2:2464:29568:27085 chr2 241573023 N chr2 241573186 N DEL 5
A00297:158:HT275DSXX:4:2478:9001:33833 chr2 241573002 N chr2 241573284 N DUP 5
A00404:155:HV27LDSXX:2:2108:3857:3286 chr2 241573002 N chr2 241573284 N DUP 5
A00404:156:HV37TDSXX:1:2356:26693:20979 chr2 241573002 N chr2 241573284 N DUP 5
A00404:156:HV37TDSXX:4:1341:28854:16579 chr2 241573002 N chr2 241573284 N DUP 5
A00404:156:HV37TDSXX:2:2465:12834:32643 chr2 241573002 N chr2 241573284 N DUP 5
A00297:158:HT275DSXX:2:1436:19596:4523 chr2 241573002 N chr2 241573284 N DUP 5
A00404:156:HV37TDSXX:3:1619:22670:1172 chr2 241573215 N chr2 241573375 N DUP 4
A00404:156:HV37TDSXX:1:2259:26946:11240 chr2 241573254 N chr2 241573374 N DUP 5
A00404:155:HV27LDSXX:4:2657:16333:17221 chr2 241573002 N chr2 241573284 N DUP 5
A00404:156:HV37TDSXX:3:1561:13964:8547 chr2 241572952 N chr2 241573357 N DEL 5
A00404:156:HV37TDSXX:2:1555:10122:13886 chr2 241572975 N chr2 241573297 N DUP 10
A00404:156:HV37TDSXX:2:1302:8169:34334 chr2 241573062 N chr2 241573306 N DEL 11
A00404:155:HV27LDSXX:4:1501:3495:9862 chr2 241573285 N chr2 241573364 N DUP 5
A00297:158:HT275DSXX:2:2672:32054:25160 chr2 241573062 N chr2 241573306 N DEL 10
A00404:156:HV37TDSXX:3:1641:32714:1658 chr2 241573062 N chr2 241573306 N DEL 10
A00404:155:HV27LDSXX:1:2516:7048:23406 chr2 241573062 N chr2 241573306 N DEL 10
A00297:158:HT275DSXX:1:1313:19144:15421 chr2 241573022 N chr2 241573306 N DEL 8
A00297:158:HT275DSXX:2:1420:28438:30827 chr2 241573022 N chr2 241573306 N DEL 5
A00404:155:HV27LDSXX:3:2468:23158:29951 chr2 241573025 N chr2 241573309 N DEL 5
A00404:155:HV27LDSXX:2:2423:32108:8594 chr2 241573026 N chr2 241573310 N DEL 5
A00404:156:HV37TDSXX:1:1319:24288:2722 chr2 241573026 N chr2 241573310 N DEL 5
A00404:155:HV27LDSXX:2:2376:2456:24690 chr2 241573284 N chr2 241573405 N DEL 10
A00404:156:HV37TDSXX:2:2619:4571:20776 chr2 241572943 N chr2 241573428 N DEL 12
A00297:158:HT275DSXX:2:2512:4010:14481 chr1 119783969 N chr1 119784034 N DEL 4
A00404:155:HV27LDSXX:4:2478:25048:8453 chrX 76218211 N chrX 76218338 N DUP 1
A00404:155:HV27LDSXX:1:1312:26648:18740 chrX 76218165 N chrX 76218422 N DEL 11
A00404:156:HV37TDSXX:4:2439:11478:34679 chr10 1944671 N chr10 1944725 N DEL 14
A00404:156:HV37TDSXX:2:2367:20925:9142 chr10 1944803 N chr10 1944855 N DUP 15
A00404:155:HV27LDSXX:3:2512:10574:29199 chr10 1944872 N chr10 1944977 N DUP 10
A00404:156:HV37TDSXX:1:1118:10556:9095 chr10 1944669 N chr10 1944877 N DEL 4
A00297:158:HT275DSXX:2:2277:20410:3145 chr10 1944824 N chr10 1944878 N DEL 6
A00297:158:HT275DSXX:1:1172:25319:6324 chr10 1944831 N chr10 1944885 N DEL 10
A00404:155:HV27LDSXX:2:1264:18656:15139 chr10 1944689 N chr10 1944950 N DEL 50
A00404:155:HV27LDSXX:2:1264:18656:15139 chr10 1944699 N chr10 1944960 N DEL 5
A00297:158:HT275DSXX:2:1536:19741:6621 chr10 1944712 N chr10 1944973 N DEL 10
A00404:155:HV27LDSXX:4:2615:1823:16423 chr3 8046528 N chr3 8046617 N DUP 8
A00404:156:HV37TDSXX:1:1406:12500:7889 chr9 2722250 N chr9 2722556 N DEL 5
A00404:156:HV37TDSXX:4:1530:23493:7106 chr9 2722162 N chr9 2722499 N DUP 5
A00297:158:HT275DSXX:1:2245:9697:30874 chr9 2722537 N chr9 2722600 N DUP 5
A00404:155:HV27LDSXX:3:1436:30816:4257 chr12 34535207 N chr12 34535969 N DUP 7
A00404:155:HV27LDSXX:3:2436:28122:6950 chr12 34535207 N chr12 34535969 N DUP 7
A00404:155:HV27LDSXX:1:2475:16179:34491 chr12 34535215 N chr12 34535557 N DUP 7
A00404:155:HV27LDSXX:4:1533:23430:29575 chr12 34535137 N chr12 34535650 N DUP 2
A00404:156:HV37TDSXX:4:1140:12264:22169 chr12 34535151 N chr12 34535665 N DEL 2
A00297:158:HT275DSXX:1:2547:32768:26960 chr12 34535152 N chr12 34535666 N DEL 2
A00404:156:HV37TDSXX:3:1118:12246:23985 chr12 34535152 N chr12 34535666 N DEL 2
A00404:155:HV27LDSXX:3:1657:9525:12258 chr18 559410 N chr18 559499 N DEL 1
A00404:156:HV37TDSXX:2:1640:14534:14732 chr7 56168144 N chr7 56168419 N DUP 8
A00404:156:HV37TDSXX:4:1364:7527:21230 chr7 56168144 N chr7 56168419 N DUP 8
A00404:155:HV27LDSXX:1:1425:23032:35587 chr7 56168134 N chr7 56168351 N DUP 2
A00404:155:HV27LDSXX:4:1164:8404:23782 chr7 56168298 N chr7 56168351 N DUP 5
A00297:158:HT275DSXX:3:2613:2193:36292 chr7 56168314 N chr7 56168367 N DEL 8
A00404:155:HV27LDSXX:1:2523:4571:20118 chr7 56168315 N chr7 56168368 N DEL 7
A00404:156:HV37TDSXX:3:1469:15655:15264 chr7 56168315 N chr7 56168368 N DEL 7
A00404:155:HV27LDSXX:2:2204:2917:12587 chr2 130758110 N chr2 130758336 N DUP 1
A00404:156:HV37TDSXX:4:1215:17381:27837 chr2 130758153 N chr2 130758384 N DEL 18
A00404:156:HV37TDSXX:3:1556:2202:29136 chr2 130758156 N chr2 130758387 N DEL 15
A00404:156:HV37TDSXX:1:2502:30138:4930 chr6 116800414 N chr6 116800514 N DEL 1
A00404:156:HV37TDSXX:4:1665:26295:12054 chr14 76539032 N chr14 76539295 N DEL 6
A00404:155:HV27LDSXX:2:1403:11632:17440 chr14 76539042 N chr14 76539412 N DEL 8
A00404:156:HV37TDSXX:4:2455:17797:35133 chr3 146635237 N chr3 146635296 N DEL 5
A00404:156:HV37TDSXX:2:1632:27923:34914 chr3 146635237 N chr3 146635296 N DEL 5
A00297:158:HT275DSXX:3:2610:17481:16736 chr3 146635469 N chr3 146635534 N DUP 15
A00404:155:HV27LDSXX:4:1532:4806:36088 chr3 146635489 N chr3 146635556 N DUP 3
A00404:156:HV37TDSXX:3:2459:21133:13197 chr11 122575082 N chr11 122575218 N DEL 21
A00297:158:HT275DSXX:1:1620:27570:6621 chr7 64856566 N chr7 64856867 N DEL 4
A00404:156:HV37TDSXX:1:1463:3486:5400 chr5 194295 N chr5 194346 N DEL 5
A00404:155:HV27LDSXX:2:1144:20907:6042 chr5 194307 N chr5 194358 N DEL 3
A00297:158:HT275DSXX:4:1218:11903:28651 chr5 194309 N chr5 194410 N DEL 1
A00404:155:HV27LDSXX:2:2216:14208:5494 chr15 96135568 N chr15 96135696 N DUP 1
A00404:156:HV37TDSXX:2:1604:6696:21637 chr15 96135711 N chr15 96135812 N DEL 5
A00297:158:HT275DSXX:1:1440:29469:20776 chr15 96135711 N chr15 96135812 N DEL 5
A00297:158:HT275DSXX:3:1530:3070:14043 chr15 96135711 N chr15 96135812 N DEL 5
A00404:156:HV37TDSXX:1:2178:18945:25254 chr9 36306027 N chr9 36306335 N DEL 5
A00404:155:HV27LDSXX:3:2503:31367:22216 chr9 36306034 N chr9 36306342 N DEL 5
A00404:155:HV27LDSXX:1:1543:25346:9001 chr9 36306039 N chr9 36306347 N DEL 1
A00404:156:HV37TDSXX:1:2673:3260:29058 chr8 144687022 N chr8 144687806 N DEL 1
A00404:155:HV27LDSXX:2:2612:25907:13009 chr8 144687028 N chr8 144687812 N DEL 8
A00404:156:HV37TDSXX:3:2339:5448:13213 chr8 144687028 N chr8 144687812 N DEL 12
A00297:158:HT275DSXX:1:1140:12237:31046 chr8 144687028 N chr8 144687812 N DEL 13
A00404:155:HV27LDSXX:1:1310:16107:32643 chr8 144687028 N chr8 144687812 N DEL 15
A00404:155:HV27LDSXX:2:2176:13991:19460 chr8 144687028 N chr8 144687812 N DEL 14
A00297:158:HT275DSXX:3:2576:29116:8046 chr8 144687028 N chr8 144687812 N DEL 15
A00404:156:HV37TDSXX:3:1315:3947:12148 chr8 144687028 N chr8 144687812 N DEL 15
A00404:155:HV27LDSXX:2:2612:17571:10410 chr8 144687028 N chr8 144687812 N DEL 8
A00404:155:HV27LDSXX:2:2147:4915:30608 chr8 144687051 N chr8 144687303 N DEL 17
A00404:156:HV37TDSXX:1:1549:13666:34741 chr8 144687051 N chr8 144687303 N DEL 18
A00404:155:HV27LDSXX:3:1218:3911:18568 chr8 144687051 N chr8 144687303 N DEL 20
A00404:155:HV27LDSXX:3:2117:30725:31845 chr8 144687051 N chr8 144687303 N DEL 20
A00297:158:HT275DSXX:4:2420:3341:33301 chr8 144687051 N chr8 144687303 N DEL 20
A00404:155:HV27LDSXX:2:1442:15094:30733 chr8 144687051 N chr8 144687303 N DEL 20
A00404:155:HV27LDSXX:1:1410:12545:3364 chr8 144687051 N chr8 144687303 N DEL 23
A00404:156:HV37TDSXX:2:1327:4869:31939 chr8 144687051 N chr8 144687303 N DEL 25
A00404:155:HV27LDSXX:3:2525:6488:11851 chr8 144687051 N chr8 144687303 N DEL 30
A00404:156:HV37TDSXX:1:1238:21233:24580 chr8 144687051 N chr8 144687303 N DEL 25
A00297:158:HT275DSXX:4:1571:29098:35289 chr8 144687072 N chr8 144687855 N DEL 39
A00404:155:HV27LDSXX:1:2176:13856:11616 chr8 144687256 N chr8 144687401 N DEL 17
A00404:155:HV27LDSXX:3:2113:12201:29450 chr8 144687198 N chr8 144687413 N DEL 5
A00404:155:HV27LDSXX:3:2503:6632:12007 chr8 144687126 N chr8 144687413 N DEL 11
A00404:155:HV27LDSXX:1:1132:3278:5916 chr8 144687126 N chr8 144687413 N DEL 14
A00404:155:HV27LDSXX:1:1132:3296:5102 chr8 144687126 N chr8 144687413 N DEL 14
A00404:156:HV37TDSXX:3:1317:14931:29105 chr8 144687222 N chr8 144687718 N DUP 25
A00297:158:HT275DSXX:1:1669:12680:22200 chr8 144687222 N chr8 144687577 N DUP 16
A00404:155:HV27LDSXX:3:2356:25527:25003 chr8 144687029 N chr8 144687917 N DUP 28
A00404:156:HV37TDSXX:3:1237:32768:14372 chr8 144687246 N chr8 144687319 N DEL 4
A00404:155:HV27LDSXX:2:2147:4915:30608 chr8 144687097 N chr8 144687239 N DUP 15
A00404:156:HV37TDSXX:1:2340:18340:22075 chr8 144687256 N chr8 144687401 N DEL 21
A00404:156:HV37TDSXX:4:2539:11577:34632 chr8 144687314 N chr8 144687915 N DUP 4
A00404:155:HV27LDSXX:4:2263:32009:6918 chr8 144687504 N chr8 144687823 N DEL 24
A00297:158:HT275DSXX:3:2528:31015:22795 chr8 144687470 N chr8 144687754 N DEL 15
A00297:158:HT275DSXX:2:1429:12888:33270 chr8 144687163 N chr8 144687233 N DUP 17
A00404:155:HV27LDSXX:2:2176:13991:19460 chr8 144687163 N chr8 144687482 N DUP 11
A00404:155:HV27LDSXX:1:1104:1633:4758 chr8 144687163 N chr8 144687482 N DUP 11
A00404:155:HV27LDSXX:4:2413:17192:15984 chr8 144687103 N chr8 144687744 N DEL 18
A00404:155:HV27LDSXX:2:1123:22309:8750 chr8 144687164 N chr8 144687805 N DEL 3
A00404:156:HV37TDSXX:4:2373:1868:31187 chr8 144687113 N chr8 144687754 N DEL 29
A00297:158:HT275DSXX:1:2408:17381:1031 chr8 144687591 N chr8 144687804 N DEL 11
A00297:158:HT275DSXX:4:2318:32497:6136 chr8 144687269 N chr8 144688050 N DEL 10
A00404:155:HV27LDSXX:3:1577:18249:32095 chr8 144687582 N chr8 144688042 N DEL 15
A00297:158:HT275DSXX:1:2664:16324:21433 chr8 144687630 N chr8 144687699 N DUP 5
A00404:156:HV37TDSXX:4:2432:32108:19554 chr8 144687630 N chr8 144687699 N DUP 5
A00404:155:HV27LDSXX:4:2319:32470:30201 chr8 144687652 N chr8 144688109 N DUP 15
A00404:155:HV27LDSXX:1:1270:8386:15577 chr8 144687630 N chr8 144687699 N DUP 5
A00297:158:HT275DSXX:4:2115:24569:5995 chr8 144687592 N chr8 144687802 N DUP 7
A00404:155:HV27LDSXX:3:1149:16116:4100 chr8 144687412 N chr8 144687731 N DEL 5
A00404:156:HV37TDSXX:3:2357:10375:19460 chr8 144687240 N chr8 144687738 N DEL 2
A00297:158:HT275DSXX:1:1249:5095:3333 chr8 144687678 N chr8 144687855 N DEL 10
A00404:155:HV27LDSXX:2:2534:1045:28729 chr8 144687808 N chr8 144688054 N DUP 10
A00404:155:HV27LDSXX:4:2669:18692:22561 chr8 144687802 N chr8 144687906 N DUP 11
A00404:155:HV27LDSXX:4:1239:12264:29935 chr8 144687752 N chr8 144688034 N DUP 22
A00297:158:HT275DSXX:3:2237:7355:4742 chr8 144687802 N chr8 144687906 N DUP 17
A00404:156:HV37TDSXX:1:2122:7762:32064 chr8 144687222 N chr8 144687965 N DUP 7
A00404:156:HV37TDSXX:2:2506:23647:1579 chr8 144687701 N chr8 144687843 N DEL 8
A00297:158:HT275DSXX:1:1646:10899:7936 chr8 144687099 N chr8 144687952 N DEL 7
A00404:155:HV27LDSXX:4:1121:26693:8797 chr19 57087943 N chr19 57088078 N DUP 2
A00404:155:HV27LDSXX:4:1121:27778:9987 chr19 57087943 N chr19 57088078 N DUP 2
A00297:158:HT275DSXX:2:2220:27019:35196 chr16 86932414 N chr16 86932580 N DUP 2
A00297:158:HT275DSXX:2:1314:16731:19257 chr16 86932582 N chr16 86932660 N DEL 5
A00404:156:HV37TDSXX:3:2521:2148:17487 chr16 86932582 N chr16 86932660 N DEL 5
A00404:156:HV37TDSXX:1:1130:17562:23954 chr16 84965781 N chr16 84965856 N DUP 5
A00297:158:HT275DSXX:1:1342:27615:36229 chr16 84965781 N chr16 84965856 N DUP 6
A00404:156:HV37TDSXX:1:1258:23339:7560 chr16 84965797 N chr16 84965866 N DEL 6
A00404:155:HV27LDSXX:1:1270:17065:31203 chr16 84965798 N chr16 84965867 N DEL 6
A00297:158:HT275DSXX:1:1113:27118:36933 chr15 20444608 N chr15 20444933 N DEL 10
A00404:156:HV37TDSXX:2:1461:2573:28244 chr15 20444659 N chr15 20444930 N DEL 5
A00297:158:HT275DSXX:4:1305:15573:17942 chr15 20444614 N chr15 20444885 N DEL 5
A00297:158:HT275DSXX:3:1606:11107:23923 chr15 20444659 N chr15 20444930 N DEL 5
A00297:158:HT275DSXX:4:1671:28763:32174 chr15 20444691 N chr15 20444908 N DEL 5
A00297:158:HT275DSXX:2:2173:1913:6590 chr15 20444664 N chr15 20444881 N DEL 5
A00297:158:HT275DSXX:4:1305:15573:17942 chr15 20444867 N chr15 20444976 N DEL 5
A00404:156:HV37TDSXX:2:1426:25120:4695 chr15 20444691 N chr15 20444962 N DEL 15
A00297:158:HT275DSXX:1:1255:15763:16172 chr17 79528401 N chr17 79528470 N DUP 5
A00404:156:HV37TDSXX:3:1245:28718:26522 chr17 79528295 N chr17 79528565 N DEL 10
A00297:158:HT275DSXX:2:1158:1606:11694 chr17 79528304 N chr17 79528574 N DEL 5
A00404:155:HV27LDSXX:2:2642:14606:12352 chr17 16939450 N chr17 16939503 N DEL 17
A00404:155:HV27LDSXX:2:1128:16107:2143 chr17 16939539 N chr17 16939611 N DEL 8
A00404:156:HV37TDSXX:3:1368:15826:36323 chr2 79982445 N chr2 79982515 N DEL 5
A00404:155:HV27LDSXX:1:2247:6813:16391 chr11 56179151 N chr11 56179210 N DEL 3
A00297:158:HT275DSXX:3:1212:3369:32597 chr16 286054 N chr16 286123 N DUP 18
A00404:155:HV27LDSXX:2:2533:14787:7780 chr16 286080 N chr16 286133 N DEL 16
A00297:158:HT275DSXX:3:1433:1877:32612 chr11 34885322 N chr11 34885390 N DUP 5
A00404:155:HV27LDSXX:1:2143:29993:1830 chr11 55616493 N chr11 55616558 N DUP 5
A00404:155:HV27LDSXX:3:1560:32344:7247 chr11 55616466 N chr11 55616529 N DEL 3
A00404:155:HV27LDSXX:4:2641:27769:27727 chr11 55616463 N chr11 55616530 N DEL 2
A00404:156:HV37TDSXX:2:2502:21305:32440 chr11 55616463 N chr11 55616530 N DEL 2
A00404:155:HV27LDSXX:2:2356:24288:12774 chr17 14431909 N chr17 14431989 N DUP 5
A00404:156:HV37TDSXX:2:2528:19849:20964 chr11 134092961 N chr11 134093106 N DUP 10
A00297:158:HT275DSXX:4:2520:31765:11788 chr11 134092887 N chr11 134093180 N DEL 5
A00404:156:HV37TDSXX:4:1528:3613:10379 chr11 68892713 N chr11 68892792 N DUP 5
A00404:155:HV27LDSXX:1:2465:24225:13917 chr11 68892713 N chr11 68892792 N DUP 5
A00404:156:HV37TDSXX:4:1159:10827:4460 chr11 68892699 N chr11 68892820 N DEL 2
A00404:156:HV37TDSXX:2:1674:25934:36918 chr11 68892721 N chr11 68892842 N DEL 15
A00404:156:HV37TDSXX:3:1130:17508:13683 chr17 41041373 N chr17 41041512 N DEL 1
A00297:158:HT275DSXX:4:1632:29975:7373 chr17 41041397 N chr17 41041536 N DEL 12
A00404:155:HV27LDSXX:1:2641:27398:35728 chr17 41041383 N chr17 41041520 N DUP 4
A00297:158:HT275DSXX:2:1172:10366:23516 chr17 41041383 N chr17 41041520 N DUP 5
A00404:156:HV37TDSXX:1:2216:31891:23343 chr17 41041397 N chr17 41041536 N DEL 45
A00404:155:HV27LDSXX:4:2361:25952:2503 chr17 41041397 N chr17 41041536 N DEL 45
A00404:155:HV27LDSXX:3:1126:26467:9064 chr17 41041397 N chr17 41041536 N DEL 45
A00404:155:HV27LDSXX:3:1126:26901:9157 chr17 41041397 N chr17 41041536 N DEL 45
A00297:158:HT275DSXX:3:1540:23113:32471 chr1 58730006 N chr1 58730226 N DUP 8
A00404:155:HV27LDSXX:3:2161:17282:26349 chr1 58730006 N chr1 58730226 N DUP 6
A00404:155:HV27LDSXX:3:2404:26802:10238 chr1 58730048 N chr1 58730144 N DEL 5
A00404:156:HV37TDSXX:4:1414:11171:11381 chr1 58730048 N chr1 58730144 N DEL 5
A00404:155:HV27LDSXX:1:2645:26567:3662 chr1 58730048 N chr1 58730144 N DEL 5
A00297:158:HT275DSXX:3:2471:1307:22388 chr1 58730048 N chr1 58730144 N DEL 5
A00297:158:HT275DSXX:3:2471:1380:22420 chr1 58730048 N chr1 58730144 N DEL 5
A00404:156:HV37TDSXX:3:1217:5059:10003 chr1 58730048 N chr1 58730144 N DEL 5
A00404:156:HV37TDSXX:3:1475:6262:14184 chr1 58730000 N chr1 58730069 N DEL 10
A00404:156:HV37TDSXX:1:2429:30725:12994 chr1 58730000 N chr1 58730069 N DEL 10
A00297:158:HT275DSXX:4:1320:25699:7451 chr1 58730000 N chr1 58730069 N DEL 10
A00404:155:HV27LDSXX:3:1553:13738:14512 chr1 58730000 N chr1 58730069 N DEL 10
A00404:155:HV27LDSXX:2:2453:14262:9064 chr1 58729956 N chr1 58730147 N DUP 3
A00404:156:HV37TDSXX:1:2159:18584:16548 chr1 58729956 N chr1 58730147 N DUP 5
A00297:158:HT275DSXX:3:1152:18204:14418 chr1 58729956 N chr1 58730147 N DUP 5
A00297:158:HT275DSXX:4:1451:5981:28009 chr1 58729956 N chr1 58730147 N DUP 5
A00404:155:HV27LDSXX:3:2629:4607:24001 chr1 58729956 N chr1 58730147 N DUP 5
A00404:156:HV37TDSXX:1:2410:24786:12007 chr1 58729956 N chr1 58730147 N DUP 5
A00404:155:HV27LDSXX:2:1273:12400:33552 chr1 58729956 N chr1 58730147 N DUP 5
A00404:156:HV37TDSXX:1:2146:29062:12273 chr1 58729956 N chr1 58730147 N DUP 5
A00404:155:HV27LDSXX:3:1171:3721:30890 chr1 58729956 N chr1 58730147 N DUP 5
A00404:155:HV27LDSXX:3:1227:23466:21089 chr1 58729956 N chr1 58730147 N DUP 5
A00297:158:HT275DSXX:1:2503:5855:35931 chr1 58729956 N chr1 58730147 N DUP 5
A00404:155:HV27LDSXX:2:2333:5258:13166 chr1 58729956 N chr1 58730147 N DUP 5
A00404:156:HV37TDSXX:1:1307:29821:13839 chr1 58729956 N chr1 58730147 N DUP 5
A00404:155:HV27LDSXX:4:1422:4291:5008 chr1 58729956 N chr1 58730147 N DUP 5
A00404:155:HV27LDSXX:4:1422:8124:6762 chr1 58729956 N chr1 58730147 N DUP 5
A00297:158:HT275DSXX:2:2654:27543:3724 chr1 58729972 N chr1 58730226 N DUP 5
A00404:156:HV37TDSXX:4:2471:9254:8594 chr1 58729972 N chr1 58730226 N DUP 5
A00404:156:HV37TDSXX:1:1122:32651:34679 chr1 58730044 N chr1 58730237 N DEL 5
A00404:155:HV27LDSXX:1:1138:8811:31187 chr1 58730044 N chr1 58730237 N DEL 5
A00404:156:HV37TDSXX:1:2533:8757:11992 chr1 58730044 N chr1 58730237 N DEL 5
A00404:155:HV27LDSXX:3:2103:3197:5431 chr1 58730044 N chr1 58730237 N DEL 5
A00404:156:HV37TDSXX:2:1227:21414:35665 chr1 58730044 N chr1 58730237 N DEL 5
A00404:156:HV37TDSXX:4:2510:23963:16845 chr1 58730044 N chr1 58730237 N DEL 5
A00404:155:HV27LDSXX:3:1206:23936:36558 chr1 58730044 N chr1 58730237 N DEL 5
A00297:158:HT275DSXX:1:1547:2682:18129 chr1 58730044 N chr1 58730237 N DEL 5
A00297:158:HT275DSXX:2:1552:20175:17049 chr1 58730044 N chr1 58730237 N DEL 5
A00404:155:HV27LDSXX:1:1459:32398:14575 chr2 89773515 N chr2 89773715 N DEL 10
A00404:156:HV37TDSXX:3:1310:32235:10786 chrX 27210670 N chrX 27210790 N DUP 7
A00404:156:HV37TDSXX:3:2315:20256:15154 chrX 27210670 N chrX 27210749 N DUP 7
A00404:156:HV37TDSXX:4:1230:9543:9345 chrX 27210670 N chrX 27210790 N DUP 7
A00404:156:HV37TDSXX:1:1634:2175:35321 chrX 27210670 N chrX 27210790 N DUP 7
A00404:155:HV27LDSXX:4:1126:24080:35900 chrX 27210670 N chrX 27210749 N DUP 7
A00404:156:HV37TDSXX:1:2362:30120:24314 chrX 27210670 N chrX 27210790 N DUP 7
A00297:158:HT275DSXX:4:1514:9670:17769 chrX 27210670 N chrX 27210749 N DUP 7
A00297:158:HT275DSXX:2:1349:30373:34867 chrX 27210670 N chrX 27210790 N DUP 7
A00404:155:HV27LDSXX:1:1326:2926:21214 chrX 27210670 N chrX 27210749 N DUP 7
A00404:156:HV37TDSXX:2:1602:28031:28933 chrX 27210670 N chrX 27210790 N DUP 7
A00404:156:HV37TDSXX:2:2374:4508:2566 chrX 27210670 N chrX 27210790 N DUP 7
A00404:156:HV37TDSXX:2:2374:3766:3317 chrX 27210670 N chrX 27210790 N DUP 7
A00404:156:HV37TDSXX:3:1176:4453:12524 chrX 27210670 N chrX 27210749 N DUP 7
A00404:156:HV37TDSXX:3:1463:20654:26303 chrX 27210670 N chrX 27210749 N DUP 7
A00404:155:HV27LDSXX:1:2453:11559:11334 chrX 27210670 N chrX 27210790 N DUP 7
A00404:156:HV37TDSXX:1:1629:18005:26443 chrX 27210670 N chrX 27210749 N DUP 7
A00297:158:HT275DSXX:3:2253:18358:17315 chrX 27210670 N chrX 27210749 N DUP 7
A00297:158:HT275DSXX:3:2253:18475:17487 chrX 27210670 N chrX 27210749 N DUP 7
A00404:156:HV37TDSXX:2:2549:26503:3176 chrX 27210670 N chrX 27210749 N DUP 7
A00404:156:HV37TDSXX:1:1137:12165:8124 chrX 27210670 N chrX 27210790 N DUP 7
A00404:155:HV27LDSXX:3:2251:6207:21073 chrX 27210670 N chrX 27210749 N DUP 7
A00297:158:HT275DSXX:1:2650:32425:30311 chrX 27210749 N chrX 27211363 N DEL 25
A00404:155:HV27LDSXX:1:2453:11559:11334 chrX 27210749 N chrX 27211363 N DEL 16
A00404:156:HV37TDSXX:2:1602:28031:28933 chrX 27210708 N chrX 27211363 N DEL 16
A00404:156:HV37TDSXX:1:2268:9878:25520 chrX 27210708 N chrX 27211363 N DEL 16
A00297:158:HT275DSXX:3:1324:4101:15890 chrX 27210709 N chrX 27211364 N DEL 13
A00404:156:HV37TDSXX:2:2374:3766:3317 chrX 27210708 N chrX 27211363 N DEL 12
A00404:156:HV37TDSXX:2:2374:4508:2566 chrX 27210708 N chrX 27211363 N DEL 12
A00404:155:HV27LDSXX:4:1511:19054:25535 chr9 41778964 N chr9 41779044 N DEL 5
A00404:155:HV27LDSXX:3:2131:10013:11162 chr9 41778964 N chr9 41779044 N DEL 9
A00404:155:HV27LDSXX:2:1205:28854:11130 chr9 41778964 N chr9 41779044 N DEL 12
A00404:155:HV27LDSXX:3:2643:26765:29747 chr9 41778938 N chr9 41779017 N DEL 2
A00404:156:HV37TDSXX:2:2101:1262:31015 chr9 41779090 N chr9 41779169 N DEL 5
A00297:158:HT275DSXX:4:2407:5828:19163 chr8 99850066 N chr8 99850305 N DEL 5
A00297:158:HT275DSXX:4:2143:29044:10050 chr8 99850305 N chr8 99850406 N DUP 5
A00404:155:HV27LDSXX:1:2507:24985:33771 chr8 99850134 N chr8 99850467 N DEL 5
A00404:155:HV27LDSXX:1:2317:6262:25958 chr8 99850134 N chr8 99850467 N DEL 5
A00404:156:HV37TDSXX:2:1516:18521:5321 chr8 99850134 N chr8 99850467 N DEL 5
A00297:158:HT275DSXX:4:2511:10899:27508 chr8 99850061 N chr8 99850430 N DUP 5
A00404:156:HV37TDSXX:1:1572:18349:19993 chr8 99850339 N chr8 99850406 N DUP 5
A00404:155:HV27LDSXX:1:1366:19271:25974 chr8 99850073 N chr8 99850380 N DEL 5
A00404:156:HV37TDSXX:4:2332:15664:18223 chr8 99850073 N chr8 99850380 N DEL 5
A00297:158:HT275DSXX:1:2226:9543:15859 chr13 113859023 N chr13 113859109 N DUP 13
A00404:156:HV37TDSXX:2:2318:24948:34929 chr13 113859035 N chr13 113859425 N DUP 1
A00297:158:HT275DSXX:3:2660:18747:4492 chr7 216032 N chr7 216117 N DUP 7
A00404:155:HV27LDSXX:2:2533:22236:10723 chr7 215991 N chr7 216076 N DUP 7
A00404:156:HV37TDSXX:2:1151:13675:17033 chr7 216136 N chr7 216267 N DUP 5
A00297:158:HT275DSXX:1:2376:17219:29246 chr7 216026 N chr7 216199 N DUP 9
A00297:158:HT275DSXX:1:2355:25925:2644 chr7 216121 N chr7 216296 N DUP 10
A00404:156:HV37TDSXX:2:1462:19759:14512 chr17 74728983 N chr17 74729061 N DEL 15
A00297:158:HT275DSXX:3:2348:6533:36417 chrX 111668373 N chrX 111668478 N DEL 3
A00404:156:HV37TDSXX:4:2361:28926:17550 chrX 111668393 N chrX 111668456 N DUP 26
A00297:158:HT275DSXX:3:2227:11930:28823 chr21 29147689 N chr21 29148037 N DEL 1
A00404:155:HV27LDSXX:1:1252:30237:6950 chr21 29147755 N chr21 29148161 N DEL 23
A00297:158:HT275DSXX:4:1217:16432:32487 chr21 29147688 N chr21 29147911 N DUP 5
A00404:156:HV37TDSXX:3:2538:30436:17848 chr21 29147666 N chr21 29148085 N DUP 7
A00297:158:HT275DSXX:3:2227:11930:28823 chr21 29147689 N chr21 29148037 N DEL 28
A00297:158:HT275DSXX:1:2613:27444:7404 chr21 29147738 N chr21 29148088 N DEL 7
A00404:155:HV27LDSXX:3:2306:8124:31814 chr21 29147738 N chr21 29148088 N DEL 7
A00404:156:HV37TDSXX:4:2128:10574:12540 chr21 29147738 N chr21 29148088 N DEL 7
A00404:155:HV27LDSXX:2:1521:28230:19288 chr21 29147738 N chr21 29148088 N DEL 7
A00297:158:HT275DSXX:2:1314:22290:10974 chr21 29147738 N chr21 29148088 N DEL 7
A00297:158:HT275DSXX:1:2318:26268:9721 chr21 29147738 N chr21 29148088 N DEL 7
A00297:158:HT275DSXX:4:2128:5367:22341 chr21 29147738 N chr21 29148088 N DEL 7
A00404:155:HV27LDSXX:4:2657:24352:25692 chr21 29148271 N chr21 29148400 N DEL 5
A00297:158:HT275DSXX:4:2173:14823:11851 chr19 3322560 N chr19 3322824 N DEL 7
A00404:156:HV37TDSXX:1:1335:3549:19695 chr19 3322605 N chr19 3322776 N DUP 5
A00404:156:HV37TDSXX:1:1240:19000:2268 chr19 3322803 N chr19 3322972 N DEL 1
A00297:158:HT275DSXX:1:2219:20166:28557 chr19 3322773 N chr19 3323014 N DEL 7
A00404:155:HV27LDSXX:3:1129:26078:13996 chr19 3322535 N chr19 3323277 N DUP 5
A00404:156:HV37TDSXX:4:2452:22290:19335 chr2 44067797 N chr2 44068070 N DEL 4
A00404:155:HV27LDSXX:2:2601:15420:7686 chr2 44067797 N chr2 44068070 N DEL 10
A00404:156:HV37TDSXX:4:1576:23827:14544 chr2 44067514 N chr2 44067727 N DEL 5
A00404:156:HV37TDSXX:4:2414:5791:32158 chr2 44067560 N chr2 44068085 N DEL 1
A00404:156:HV37TDSXX:1:1531:2781:13510 chr10 42088978 N chr10 42089570 N DUP 5
A00297:158:HT275DSXX:1:1470:16984:26146 chr10 42088923 N chr10 42089540 N DEL 5
A00404:155:HV27LDSXX:3:2156:15221:2174 chr10 42089217 N chr10 42089808 N DUP 10
A00404:156:HV37TDSXX:1:2402:7681:24032 chr10 42089424 N chr10 42089570 N DUP 5
A00404:156:HV37TDSXX:2:2414:3495:21042 chr10 42089050 N chr10 42089230 N DEL 2
A00404:156:HV37TDSXX:1:1531:2781:13510 chr10 42088664 N chr10 42089281 N DEL 3
A00404:156:HV37TDSXX:1:2311:10836:21261 chr10 42088663 N chr10 42089228 N DEL 15
A00404:156:HV37TDSXX:2:2435:15926:1924 chr10 42088890 N chr10 42089579 N DEL 5
A00297:158:HT275DSXX:4:1676:27932:2174 chr10 42088617 N chr10 42089283 N DEL 2
A00297:158:HT275DSXX:3:1114:20989:22780 chr10 42088890 N chr10 42089579 N DEL 5
A00297:158:HT275DSXX:1:1202:13123:3959 chr10 42089057 N chr10 42089578 N DUP 2
A00297:158:HT275DSXX:3:1410:10601:11929 chr10 42088576 N chr10 42089580 N DUP 5
A00297:158:HT275DSXX:1:2354:15691:30827 chr10 42088626 N chr10 42089581 N DUP 5
A00404:155:HV27LDSXX:3:1134:18430:24298 chr10 42089050 N chr10 42089230 N DEL 2
A00404:156:HV37TDSXX:3:1209:21558:4883 chr10 42088663 N chr10 42089228 N DEL 15
A00404:155:HV27LDSXX:2:1374:24153:13636 chr10 42088697 N chr10 42089360 N DUP 6
A00297:158:HT275DSXX:1:1222:1145:23610 chr10 42089269 N chr10 42089860 N DUP 5
A00404:155:HV27LDSXX:2:2610:19497:15311 chr10 42088697 N chr10 42089360 N DUP 6
A00297:158:HT275DSXX:4:2124:28989:16752 chr10 42088869 N chr10 42089486 N DEL 3
A00297:158:HT275DSXX:4:2208:26847:7592 chr10 42088610 N chr10 42089276 N DEL 9
A00404:155:HV27LDSXX:1:2543:32470:29105 chr10 42088924 N chr10 42089541 N DEL 5
A00297:158:HT275DSXX:3:1423:15989:36886 chr10 42088765 N chr10 42089601 N DEL 5
A00404:155:HV27LDSXX:4:1276:3405:3568 chr10 42088978 N chr10 42089570 N DUP 5
A00404:155:HV27LDSXX:2:1242:9516:28557 chr10 42088912 N chr10 42089667 N DUP 1
A00404:155:HV27LDSXX:3:1650:6994:18333 chr10 42088630 N chr10 42089296 N DEL 5
A00404:156:HV37TDSXX:1:1156:32624:3223 chr10 42089223 N chr10 42089814 N DUP 9
A00404:156:HV37TDSXX:2:2342:5348:17895 chr10 42088918 N chr10 42089535 N DEL 5
A00404:156:HV37TDSXX:1:1531:3658:12367 chr10 42088978 N chr10 42089570 N DUP 5
A00297:158:HT275DSXX:4:2658:9299:8547 chr10 42089248 N chr10 42089763 N DEL 1
A00404:156:HV37TDSXX:1:2224:27968:8124 chr10 42088694 N chr10 42089233 N DEL 14
A00297:158:HT275DSXX:4:2658:9299:8547 chr10 42088998 N chr10 42089592 N DEL 10
A00404:155:HV27LDSXX:3:1447:7997:28995 chr10 42088705 N chr10 42089541 N DEL 6
A00404:156:HV37TDSXX:2:2125:12933:29716 chr10 42089217 N chr10 42089808 N DUP 10
A00404:155:HV27LDSXX:2:1256:29369:7576 chr10 42088924 N chr10 42089541 N DEL 15
A00404:156:HV37TDSXX:4:2543:2076:33646 chr10 42088590 N chr10 42089596 N DEL 5
A00404:156:HV37TDSXX:4:1644:9878:12085 chr10 42089057 N chr10 42089578 N DUP 2
A00404:155:HV27LDSXX:4:1125:32796:10379 chr10 42089281 N chr10 42089872 N DUP 4
A00404:155:HV27LDSXX:3:1106:24795:4100 chr10 42088918 N chr10 42089535 N DEL 5
A00404:156:HV37TDSXX:4:1429:21856:19867 chr10 42088663 N chr10 42089228 N DEL 14
A00404:155:HV27LDSXX:4:1217:21314:8061 chr10 42088639 N chr10 42089596 N DEL 6
A00404:155:HV27LDSXX:1:1137:11153:12320 chr10 42089120 N chr10 42089712 N DUP 5
A00404:156:HV37TDSXX:4:1462:12328:12258 chr10 42089073 N chr10 42089573 N DEL 3
A00297:158:HT275DSXX:4:2315:21124:29465 chr10 42089217 N chr10 42089808 N DUP 10
A00404:156:HV37TDSXX:3:1346:6741:17331 chr10 42089281 N chr10 42089872 N DUP 5
A00404:155:HV27LDSXX:2:1502:9335:35853 chr10 42088978 N chr10 42089570 N DUP 5
A00297:158:HT275DSXX:2:1342:10239:1501 chr10 42088921 N chr10 42089538 N DEL 5
A00297:158:HT275DSXX:3:2673:3278:13495 chr10 42088924 N chr10 42089541 N DEL 5
A00404:155:HV27LDSXX:4:1433:2329:28072 chr10 42089455 N chr10 42089646 N DUP 4
A00404:156:HV37TDSXX:2:1155:12481:20979 chr10 42089120 N chr10 42089712 N DUP 5
A00404:156:HV37TDSXX:3:1562:19886:26725 chr10 42088978 N chr10 42089570 N DUP 5
A00404:156:HV37TDSXX:3:2510:28565:17769 chr10 42088538 N chr10 42089279 N DEL 5
A00404:156:HV37TDSXX:2:2324:16025:6699 chr10 42089135 N chr10 42089727 N DUP 8
A00404:156:HV37TDSXX:1:1262:8847:13401 chr10 42088626 N chr10 42089581 N DUP 5
A00404:156:HV37TDSXX:2:1123:22318:9455 chr10 42089281 N chr10 42089872 N DUP 5
A00404:155:HV27LDSXX:2:1509:32416:11913 chr10 42088952 N chr10 42089546 N DEL 1
A00404:155:HV27LDSXX:1:2218:4038:34006 chr10 42088663 N chr10 42089228 N DEL 15
A00404:155:HV27LDSXX:1:2525:23086:33646 chr10 42088663 N chr10 42089228 N DEL 15
A00404:156:HV37TDSXX:2:1630:20763:18630 chr10 42089148 N chr10 42089739 N DUP 13
A00297:158:HT275DSXX:3:1659:14443:14168 chr10 42088912 N chr10 42089667 N DUP 1
A00404:155:HV27LDSXX:3:2154:7021:10645 chr10 42089129 N chr10 42089721 N DUP 1
A00297:158:HT275DSXX:1:2163:5584:14732 chr10 42088706 N chr10 42089542 N DEL 5
A00297:158:HT275DSXX:4:2116:18891:31892 chr10 42089217 N chr10 42089808 N DUP 10
A00404:155:HV27LDSXX:2:1654:19108:35744 chr10 42088696 N chr10 42089235 N DEL 11
A00297:158:HT275DSXX:1:1350:22670:24940 chr10 42088951 N chr10 42089545 N DEL 2
A00297:158:HT275DSXX:4:1449:24740:10050 chr10 42088998 N chr10 42089592 N DEL 7
A00404:155:HV27LDSXX:3:2642:28763:21433 chr10 42088978 N chr10 42089570 N DUP 5
A00404:155:HV27LDSXX:3:2138:19009:15154 chr10 42089120 N chr10 42089712 N DUP 5
A00404:156:HV37TDSXX:2:2220:8088:22482 chr10 42088664 N chr10 42089281 N DEL 3
A00404:156:HV37TDSXX:4:2327:27498:14732 chr10 42089071 N chr10 42089594 N DEL 5
A00404:155:HV27LDSXX:4:1110:8359:5791 chr10 42088774 N chr10 42089438 N DUP 8
A00404:156:HV37TDSXX:1:1531:3658:12367 chr10 42088664 N chr10 42089281 N DEL 3
A00404:156:HV37TDSXX:4:1661:20573:18928 chr10 42089269 N chr10 42089860 N DUP 5
A00297:158:HT275DSXX:2:2153:23204:2628 chr10 42089269 N chr10 42089860 N DUP 5
A00404:155:HV27LDSXX:4:2660:7961:13495 chr10 42089148 N chr10 42089739 N DUP 10
A00404:156:HV37TDSXX:4:2327:27425:14544 chr10 42089071 N chr10 42089594 N DEL 5
A00297:158:HT275DSXX:3:1365:14633:36886 chr10 42088616 N chr10 42089282 N DEL 3
A00404:156:HV37TDSXX:3:2423:29387:33473 chr10 42088774 N chr10 42089438 N DUP 6
A00297:158:HT275DSXX:2:1547:14814:7138 chr10 42088590 N chr10 42089596 N DEL 5
A00297:158:HT275DSXX:3:1377:32868:4085 chr10 42089275 N chr10 42089866 N DUP 10
A00404:155:HV27LDSXX:4:1377:4291:15468 chr10 42088891 N chr10 42089580 N DEL 5
A00404:155:HV27LDSXX:2:2343:26494:31313 chr10 42089330 N chr10 42089717 N DUP 4
A00297:158:HT275DSXX:1:2472:16043:19758 chr10 42088949 N chr10 42089566 N DEL 5
A00404:155:HV27LDSXX:2:2340:15917:3474 chr10 42089228 N chr10 42089328 N DUP 16
A00297:158:HT275DSXX:2:1272:5195:11459 chr10 42088695 N chr10 42089234 N DEL 12
A00297:158:HT275DSXX:2:2616:28583:9846 chr10 42089071 N chr10 42089594 N DEL 5
A00404:155:HV27LDSXX:4:2177:24216:35321 chr10 42088615 N chr10 42089281 N DEL 4
A00404:156:HV37TDSXX:4:1464:10230:22842 chr10 42089424 N chr10 42089572 N DEL 1
A00404:155:HV27LDSXX:1:2543:32470:29105 chr10 42089279 N chr10 42089870 N DUP 5
A00297:158:HT275DSXX:3:1531:2528:3959 chr10 42089269 N chr10 42089860 N DUP 5
A00404:156:HV37TDSXX:3:2165:4309:22200 chr10 42088774 N chr10 42089438 N DUP 5
A00404:156:HV37TDSXX:1:1470:5086:28839 chr10 42089072 N chr10 42089595 N DEL 5
A00404:156:HV37TDSXX:3:1223:3341:5212 chr10 42088921 N chr10 42089538 N DEL 5
A00404:155:HV27LDSXX:4:2344:16604:26428 chr10 42088998 N chr10 42089592 N DEL 10
A00297:158:HT275DSXX:3:2276:6903:23657 chr10 42089120 N chr10 42089712 N DUP 5
A00404:156:HV37TDSXX:1:1153:24623:24940 chr10 42088923 N chr10 42089540 N DEL 5
A00404:156:HV37TDSXX:3:2464:25147:18771 chr10 42088951 N chr10 42089545 N DEL 2
A00297:158:HT275DSXX:1:2116:8287:33786 chr10 42088998 N chr10 42089592 N DEL 5
A00404:156:HV37TDSXX:3:1308:9372:22200 chr10 42088543 N chr10 42089454 N DEL 5
A00297:158:HT275DSXX:4:2575:16984:28588 chr10 42089135 N chr10 42089727 N DUP 7
A00297:158:HT275DSXX:2:2367:24171:11193 chr10 42088978 N chr10 42089570 N DUP 5
A00297:158:HT275DSXX:4:2448:27896:12571 chr10 42088774 N chr10 42089438 N DUP 5
A00404:156:HV37TDSXX:1:2170:20609:31516 chr10 42088949 N chr10 42089543 N DEL 4
A00404:156:HV37TDSXX:1:1441:29704:20494 chr10 42089129 N chr10 42089721 N DUP 1
A00404:155:HV27LDSXX:4:1615:26675:24518 chr10 42089217 N chr10 42089808 N DUP 15
A00404:155:HV27LDSXX:1:1546:19280:1626 chr10 42088611 N chr10 42089277 N DEL 8
A00297:158:HT275DSXX:1:2219:2853:12727 chr10 42088646 N chr10 42089263 N DEL 7
A00404:156:HV37TDSXX:2:2143:1054:14027 chr10 42088673 N chr10 42088793 N DUP 1
A00297:158:HT275DSXX:3:1531:23990:23093 chr10 42089217 N chr10 42089808 N DUP 10
A00297:158:HT275DSXX:4:1415:13621:15342 chr10 42088998 N chr10 42089592 N DEL 5
A00404:156:HV37TDSXX:3:2141:8061:24502 chr10 42088708 N chr10 42089636 N DUP 1
A00404:155:HV27LDSXX:2:1466:21386:31328 chr10 42088978 N chr10 42089570 N DUP 5
A00404:156:HV37TDSXX:4:1235:1940:3004 chr10 42088774 N chr10 42089438 N DUP 8
A00404:155:HV27LDSXX:1:2247:1063:33364 chr10 42088923 N chr10 42089540 N DEL 5
A00404:155:HV27LDSXX:3:2417:1913:33646 chr10 42088625 N chr10 42089291 N DEL 10
A00404:156:HV37TDSXX:3:2308:24623:19429 chr10 42088792 N chr10 42089638 N DUP 2
A00404:155:HV27LDSXX:3:2608:30734:31986 chr10 42089424 N chr10 42089570 N DUP 5
A00297:158:HT275DSXX:2:2106:26142:28886 chr10 42088590 N chr10 42089596 N DEL 5
A00297:158:HT275DSXX:2:2202:20754:1548 chr10 42089269 N chr10 42089860 N DUP 5
A00404:156:HV37TDSXX:1:2269:3106:21934 chr10 42088998 N chr10 42089592 N DEL 5
A00404:155:HV27LDSXX:2:1334:6334:7639 chr10 42089228 N chr10 42089328 N DUP 16
A00404:156:HV37TDSXX:1:2639:32750:26177 chr10 42088663 N chr10 42089228 N DEL 15
A00404:156:HV37TDSXX:3:1561:28212:18787 chr10 42089269 N chr10 42089860 N DUP 5
A00404:156:HV37TDSXX:4:1150:23158:3364 chr10 42089269 N chr10 42089860 N DUP 5
A00297:158:HT275DSXX:4:2575:16984:28588 chr10 42088615 N chr10 42089281 N DEL 4
A00404:155:HV27LDSXX:2:2532:26187:7639 chr10 42089425 N chr10 42089571 N DUP 1
A00404:155:HV27LDSXX:4:2137:4029:4961 chr10 42088774 N chr10 42089438 N DUP 10
A00404:156:HV37TDSXX:2:1419:12527:31955 chr10 42089072 N chr10 42089595 N DEL 5
A00404:156:HV37TDSXX:3:1139:7880:35149 chr10 42088674 N chr10 42089580 N DUP 2
A00404:156:HV37TDSXX:2:2178:17056:26835 chr10 42088992 N chr10 42089586 N DEL 1
A00404:156:HV37TDSXX:3:2337:20618:25770 chr10 42088626 N chr10 42089581 N DUP 5
A00404:155:HV27LDSXX:4:2607:18665:2096 chr10 42088950 N chr10 42089544 N DEL 3
A00404:156:HV37TDSXX:3:1568:21197:26428 chr10 42089288 N chr10 42089578 N DUP 5
A00404:155:HV27LDSXX:1:2238:5132:4116 chr10 42089148 N chr10 42089739 N DUP 5
A00404:155:HV27LDSXX:2:1361:19208:13307 chr10 42089135 N chr10 42089727 N DUP 12
A00404:155:HV27LDSXX:4:1265:26512:20541 chr10 42088718 N chr10 42089381 N DUP 6
A00404:156:HV37TDSXX:3:2550:5041:21997 chr10 42089135 N chr10 42089727 N DUP 7
A00404:155:HV27LDSXX:2:2376:8901:12367 chr10 42089027 N chr10 42089619 N DUP 7
A00297:158:HT275DSXX:4:2512:11776:33191 chr10 42088792 N chr10 42089638 N DUP 2
A00404:155:HV27LDSXX:3:1124:8115:24158 chr10 42088543 N chr10 42089454 N DEL 5
A00404:155:HV27LDSXX:4:2137:4020:4946 chr10 42088774 N chr10 42089438 N DUP 10
A00404:155:HV27LDSXX:2:1140:11406:24220 chr10 42088590 N chr10 42089596 N DEL 5
A00297:158:HT275DSXX:3:2409:24939:15311 chr10 42088613 N chr10 42089279 N DEL 6
A00297:158:HT275DSXX:2:2663:4336:15859 chr10 42088588 N chr10 42089594 N DEL 5
A00404:156:HV37TDSXX:3:2510:28565:17769 chr10 42088590 N chr10 42089596 N DEL 5
A00404:156:HV37TDSXX:1:2622:20103:22874 chr10 42088618 N chr10 42089284 N DEL 1
A00404:156:HV37TDSXX:1:2241:21016:7921 chr10 42088543 N chr10 42089454 N DEL 5
A00404:156:HV37TDSXX:2:1143:20383:30655 chr10 42089057 N chr10 42089578 N DUP 2
A00404:156:HV37TDSXX:1:2241:21106:9330 chr10 42088543 N chr10 42089454 N DEL 5
A00297:158:HT275DSXX:2:1354:32434:9940 chr10 42088978 N chr10 42089570 N DUP 5
A00404:155:HV27LDSXX:1:2112:13530:34757 chr10 42089148 N chr10 42089739 N DUP 8
A00404:156:HV37TDSXX:4:2123:1687:33755 chr10 42089057 N chr10 42089578 N DUP 3
A00404:156:HV37TDSXX:2:1467:5611:34851 chr10 42088918 N chr10 42089535 N DEL 5
A00297:158:HT275DSXX:4:2210:19434:2362 chr10 42088814 N chr10 42089431 N DEL 25
A00297:158:HT275DSXX:4:1402:26359:30796 chr10 42088629 N chr10 42089540 N DEL 11
A00297:158:HT275DSXX:3:1449:9408:21104 chr10 42089217 N chr10 42089808 N DUP 14
A00404:156:HV37TDSXX:2:1101:18855:28698 chr10 42089120 N chr10 42089712 N DUP 5
A00404:156:HV37TDSXX:2:2151:27010:17206 chr10 42088945 N chr10 42089539 N DEL 8
A00297:158:HT275DSXX:1:2315:18168:13041 chr10 42088774 N chr10 42089438 N DUP 7
A00404:156:HV37TDSXX:4:2347:6560:12258 chr10 42089071 N chr10 42089594 N DEL 5
A00404:155:HV27LDSXX:1:2548:23411:21277 chr10 42088626 N chr10 42089581 N DUP 5
A00297:158:HT275DSXX:3:1352:1515:33802 chr10 42088992 N chr10 42089586 N DEL 1
A00404:156:HV37TDSXX:2:1324:29722:9126 chr10 42089217 N chr10 42089808 N DUP 15
A00404:156:HV37TDSXX:2:1560:7518:20055 chr10 42088892 N chr10 42089581 N DEL 5
A00404:155:HV27LDSXX:4:1613:10529:16125 chr10 42088897 N chr10 42089586 N DEL 6
A00404:156:HV37TDSXX:2:2105:3351:20478 chr10 42088645 N chr10 42089602 N DEL 5
A00297:158:HT275DSXX:4:2176:24071:9048 chr10 42089269 N chr10 42089860 N DUP 5
A00404:155:HV27LDSXX:1:2112:13521:34710 chr10 42089148 N chr10 42089739 N DUP 8
A00297:158:HT275DSXX:1:1202:12147:1266 chr10 42089057 N chr10 42089578 N DUP 2
A00404:155:HV27LDSXX:2:1174:24975:11334 chr10 42089275 N chr10 42089866 N DUP 5
A00297:158:HT275DSXX:2:1226:16712:26490 chr10 42088923 N chr10 42089540 N DEL 5
A00404:156:HV37TDSXX:4:1564:23628:27164 chr10 42088695 N chr10 42089234 N DEL 13
A00297:158:HT275DSXX:4:2474:6858:16845 chr10 42088626 N chr10 42089581 N DUP 5
A00404:156:HV37TDSXX:4:2519:14082:4022 chr10 42088630 N chr10 42089296 N DEL 5
A00404:156:HV37TDSXX:3:1342:7527:4726 chr10 42088938 N chr10 42089670 N DUP 2
A00404:156:HV37TDSXX:4:2543:1732:33520 chr10 42088590 N chr10 42089596 N DEL 5
A00404:155:HV27LDSXX:3:2460:30246:18803 chr10 42089217 N chr10 42089808 N DUP 10
A00404:156:HV37TDSXX:1:2121:6470:29606 chr10 42088951 N chr10 42089545 N DEL 2
A00404:155:HV27LDSXX:1:1430:26187:4445 chr10 42088938 N chr10 42089670 N DUP 3
A00404:155:HV27LDSXX:1:2152:6289:11099 chr10 42088463 N chr10 42089691 N DUP 1
A00404:156:HV37TDSXX:4:2117:27281:30076 chr10 42088998 N chr10 42089592 N DEL 5
A00297:158:HT275DSXX:3:1216:7979:3881 chr10 42088618 N chr10 42089284 N DEL 1
A00404:156:HV37TDSXX:2:2638:32931:7263 chr10 42088626 N chr10 42089581 N DUP 5
A00404:155:HV27LDSXX:4:1103:1027:28573 chr10 42088950 N chr10 42089544 N DEL 3
A00404:156:HV37TDSXX:2:1350:3803:33818 chr10 42088928 N chr10 42089300 N DEL 5
A00297:158:HT275DSXX:1:1253:2031:12774 chr10 42089217 N chr10 42089808 N DUP 15
A00404:156:HV37TDSXX:3:1112:31837:2613 chr10 42089224 N chr10 42089815 N DUP 8
A00404:155:HV27LDSXX:2:1122:6424:28839 chr10 42088543 N chr10 42089454 N DEL 5
A00404:155:HV27LDSXX:3:2409:27245:17206 chr10 42089051 N chr10 42089231 N DEL 1
A00404:155:HV27LDSXX:4:1341:30020:25363 chr10 42089304 N chr10 42089691 N DUP 5
A00404:156:HV37TDSXX:2:1617:21269:9549 chr10 42088978 N chr10 42089570 N DUP 9
A00404:156:HV37TDSXX:3:2613:8477:33176 chr10 42089207 N chr10 42089286 N DEL 2
A00297:158:HT275DSXX:1:1660:9155:2848 chr10 42088613 N chr10 42089279 N DEL 6
A00297:158:HT275DSXX:4:1319:14669:12743 chr10 42088978 N chr10 42089570 N DUP 5
A00297:158:HT275DSXX:2:1417:19913:4695 chr10 42088694 N chr10 42089233 N DEL 7
A00297:158:HT275DSXX:2:2212:23484:7467 chr10 42088998 N chr10 42089592 N DEL 5
A00404:155:HV27LDSXX:2:2646:23755:31234 chr10 42089281 N chr10 42089872 N DUP 5
A00404:156:HV37TDSXX:4:2356:11207:6057 chr10 42088957 N chr10 42089551 N DEL 1
A00404:155:HV27LDSXX:4:1110:8359:5791 chr10 42088918 N chr10 42089535 N DEL 5
A00404:156:HV37TDSXX:4:1661:20573:18928 chr10 42088992 N chr10 42089586 N DEL 1
A00404:156:HV37TDSXX:2:1526:21124:18474 chr10 42088918 N chr10 42089535 N DEL 5
A00404:156:HV37TDSXX:3:2553:22616:25316 chr10 42088463 N chr10 42089691 N DUP 1
A00404:156:HV37TDSXX:3:2372:11433:24236 chr10 42088918 N chr10 42089535 N DEL 5
A00297:158:HT275DSXX:1:2632:26820:11522 chr10 42088951 N chr10 42089545 N DEL 2
A00404:155:HV27LDSXX:3:1178:24442:9377 chr10 42089049 N chr10 42089229 N DEL 3
A00404:155:HV27LDSXX:4:1341:30210:25723 chr10 42089304 N chr10 42089691 N DUP 5
A00297:158:HT275DSXX:2:2636:20265:8093 chr10 42089269 N chr10 42089860 N DUP 5
A00404:155:HV27LDSXX:1:1539:2483:10019 chr10 42089065 N chr10 42089271 N DEL 6
A00297:158:HT275DSXX:2:2367:24171:11193 chr10 42088612 N chr10 42089278 N DEL 7
A00297:158:HT275DSXX:1:1214:15347:15702 chr10 42088578 N chr10 42089389 N DUP 4
A00404:155:HV27LDSXX:4:2505:4309:23860 chr10 42088912 N chr10 42089667 N DUP 1
A00297:158:HT275DSXX:3:2355:5095:15389 chr10 42089057 N chr10 42089578 N DUP 2
A00404:156:HV37TDSXX:2:2258:25283:17785 chr10 42088576 N chr10 42089580 N DUP 4
A00404:156:HV37TDSXX:4:1636:29441:18223 chr10 42088663 N chr10 42089228 N DEL 15
A00404:155:HV27LDSXX:2:2462:32009:11271 chr10 42088612 N chr10 42089278 N DEL 7
A00404:156:HV37TDSXX:2:1630:20754:18615 chr10 42089155 N chr10 42089746 N DUP 13
A00297:158:HT275DSXX:1:1329:11198:7921 chr10 42088589 N chr10 42089595 N DEL 5
A00404:155:HV27LDSXX:2:2351:10248:25316 chr10 42088952 N chr10 42089546 N DEL 1
A00404:155:HV27LDSXX:4:2463:20998:20165 chr10 42089270 N chr10 42089861 N DUP 5
A00404:155:HV27LDSXX:4:2615:28438:18991 chr10 42089217 N chr10 42089808 N DUP 15
A00404:156:HV37TDSXX:1:1234:6479:24361 chr10 42089438 N chr10 42089631 N DEL 14
A00404:156:HV37TDSXX:1:2318:29749:33786 chr10 42088717 N chr10 42089380 N DUP 6
A00404:155:HV27LDSXX:1:2171:23701:26036 chr10 42089129 N chr10 42089721 N DUP 1
A00404:156:HV37TDSXX:1:2467:26169:28369 chr10 42089424 N chr10 42089570 N DUP 5
A00297:158:HT275DSXX:3:2676:5773:22482 chr10 42088626 N chr10 42089581 N DUP 5
A00404:155:HV27LDSXX:2:2340:17852:2942 chr10 42089228 N chr10 42089328 N DUP 16
A00404:155:HV27LDSXX:1:1477:19515:12555 chr10 42088696 N chr10 42089235 N DEL 11
A00404:155:HV27LDSXX:2:2610:19497:15311 chr10 42088992 N chr10 42089586 N DEL 1
A00404:155:HV27LDSXX:1:1626:23628:2487 chr10 42088706 N chr10 42089542 N DEL 5
A00404:155:HV27LDSXX:2:1178:20907:8891 chr10 42089057 N chr10 42089578 N DUP 3
A00404:155:HV27LDSXX:4:2343:11632:1752 chr10 42089288 N chr10 42089578 N DUP 5
A00404:156:HV37TDSXX:2:2436:30246:32769 chr10 42088618 N chr10 42089284 N DEL 1
A00404:155:HV27LDSXX:3:1444:13259:1971 chr10 42088998 N chr10 42089592 N DEL 5
A00404:156:HV37TDSXX:2:1156:14407:3959 chr10 42088626 N chr10 42089581 N DUP 5
A00404:156:HV37TDSXX:1:2545:2157:22106 chr10 42088795 N chr10 42089580 N DUP 5
A00297:158:HT275DSXX:4:1272:4770:24533 chr10 42089228 N chr10 42089328 N DUP 16
A00404:156:HV37TDSXX:4:1209:18521:15436 chr10 42089027 N chr10 42089619 N DUP 5
A00404:156:HV37TDSXX:3:1209:22092:4147 chr10 42088663 N chr10 42089228 N DEL 15
A00297:158:HT275DSXX:4:2559:31268:16689 chr10 42089075 N chr10 42089693 N DUP 14
A00404:156:HV37TDSXX:4:2176:13196:22373 chr10 42089269 N chr10 42089860 N DUP 5
A00297:158:HT275DSXX:4:2550:20618:3756 chrX 130504630 N chrX 130504682 N DEL 7
A00297:158:HT275DSXX:1:2136:8892:30514 chrX 130504623 N chrX 130504749 N DUP 5
A00297:158:HT275DSXX:4:1402:6225:2566 chrX 130504540 N chrX 130504594 N DUP 15
A00404:155:HV27LDSXX:4:2145:15230:31970 chrX 130504716 N chrX 130504841 N DUP 4
A00404:155:HV27LDSXX:1:2467:5611:33818 chr12 7590008 N chr12 7590182 N DUP 5
A00297:158:HT275DSXX:2:2231:26133:23860 chr12 7589989 N chr12 7590114 N DUP 11
A00297:158:HT275DSXX:4:1233:9796:4523 chr12 7589989 N chr12 7590114 N DUP 11
A00404:155:HV27LDSXX:4:2635:23068:22592 chr12 7589989 N chr12 7590114 N DUP 11
A00404:155:HV27LDSXX:4:1569:20410:26036 chr12 7589941 N chr12 7590039 N DEL 3
A00404:155:HV27LDSXX:4:1569:21052:25958 chr12 7589941 N chr12 7590039 N DEL 3
A00404:155:HV27LDSXX:4:1569:21178:17910 chr12 7589941 N chr12 7590039 N DEL 3
A00404:156:HV37TDSXX:1:1653:2817:31172 chr12 7589889 N chr12 7590063 N DUP 5
A00404:155:HV27LDSXX:3:1210:2736:14058 chr12 7589955 N chr12 7590131 N DEL 10
A00404:155:HV27LDSXX:3:1401:21766:7404 chr12 7589962 N chr12 7590138 N DEL 10
A00297:158:HT275DSXX:4:2528:27281:8970 chr12 7589955 N chr12 7590131 N DEL 10
A00404:156:HV37TDSXX:2:1668:25780:19272 chr12 7589955 N chr12 7590131 N DEL 10
A00297:158:HT275DSXX:4:2153:15320:29684 chr20 62172905 N chr20 62173021 N DUP 5
A00404:155:HV27LDSXX:2:2611:30825:16454 chr20 62172905 N chr20 62173021 N DUP 5
A00404:156:HV37TDSXX:2:2129:15817:34898 chr20 62172905 N chr20 62173021 N DUP 5
A00297:158:HT275DSXX:1:2254:12120:12931 chr4 8792336 N chr4 8792467 N DUP 2
A00404:155:HV27LDSXX:4:2378:7401:16376 chr7 66231173 N chr7 66231334 N DEL 15
A00404:156:HV37TDSXX:1:2512:18819:10097 chr7 5565855 N chr7 5566022 N DEL 3
A00404:156:HV37TDSXX:1:2121:24966:15358 chr19 46436400 N chr19 46436717 N DEL 2
A00404:156:HV37TDSXX:3:2519:12897:24893 chr8 54500563 N chr8 54500808 N DUP 7
A00297:158:HT275DSXX:3:1235:28673:12195 chr8 54500630 N chr8 54500813 N DEL 7
A00297:158:HT275DSXX:2:1161:14082:11318 chr8 54500631 N chr8 54500814 N DEL 6
A00404:155:HV27LDSXX:2:1552:3775:13636 chr15 80152646 N chr15 80152932 N DEL 5
A00404:155:HV27LDSXX:3:2206:3794:34898 chr13 112832014 N chr13 112832064 N DUP 1
A00404:156:HV37TDSXX:3:2455:27688:11428 chr6 33060317 N chr6 33060470 N DUP 12
A00404:156:HV37TDSXX:3:1310:8965:28228 chr10 129930484 N chr10 129930872 N DEL 3
A00297:158:HT275DSXX:1:2662:21712:7560 chr10 129930610 N chr10 129930941 N DEL 13
A00297:158:HT275DSXX:1:2662:21712:7560 chr10 129930610 N chr10 129930941 N DEL 17
A00404:156:HV37TDSXX:1:1425:19795:34491 chr10 129930641 N chr10 129930756 N DEL 5
A00404:156:HV37TDSXX:1:1533:30318:16673 chr10 129930811 N chr10 129931034 N DEL 5
A00404:156:HV37TDSXX:4:2158:19642:19789 chr21 40182692 N chr21 40182920 N DEL 3
A00404:156:HV37TDSXX:1:1244:1759:7200 chr21 40182745 N chr21 40182973 N DEL 5
A00297:158:HT275DSXX:4:1134:5385:36401 chr21 40182745 N chr21 40182973 N DEL 5
A00297:158:HT275DSXX:4:2402:5059:27352 chr21 40182767 N chr21 40182883 N DUP 19
A00404:155:HV27LDSXX:2:2349:4661:9596 chr21 40182880 N chr21 40183021 N DEL 10
A00297:158:HT275DSXX:3:2408:14118:2519 chr21 40182904 N chr21 40183131 N DUP 12
A00404:156:HV37TDSXX:3:1265:3757:2863 chr21 40182820 N chr21 40182877 N DUP 9
A00404:155:HV27LDSXX:4:2270:11162:24518 chr21 40182849 N chr21 40182903 N DUP 15
A00297:158:HT275DSXX:1:2626:11659:19179 chr21 40182777 N chr21 40182947 N DUP 7
A00404:156:HV37TDSXX:3:2267:4481:12414 chr21 40182827 N chr21 40183054 N DEL 12
A00297:158:HT275DSXX:1:1655:7880:23844 chr21 40182947 N chr21 40183033 N DEL 5
A00297:158:HT275DSXX:1:2273:11704:34225 chr21 40182849 N chr21 40183046 N DEL 9
A00404:156:HV37TDSXX:2:1524:20482:27853 chr21 40182708 N chr21 40182964 N DEL 12
A00297:158:HT275DSXX:4:2609:15221:24972 chr21 40182767 N chr21 40183135 N DUP 29
A00404:156:HV37TDSXX:1:1533:2645:26490 chr21 40182750 N chr21 40183146 N DUP 5
A00404:155:HV27LDSXX:4:2541:15374:1157 chr21 40182738 N chr21 40182880 N DUP 28
A00297:158:HT275DSXX:3:2623:22733:31876 chr21 40182877 N chr21 40183047 N DUP 11
A00404:155:HV27LDSXX:2:1549:9769:33004 chr21 40182776 N chr21 40182946 N DUP 14
A00297:158:HT275DSXX:4:1578:26829:19805 chr21 40183022 N chr21 40183279 N DEL 8
A00404:156:HV37TDSXX:3:2459:11939:33692 chr21 40182946 N chr21 40183202 N DEL 5
A00404:156:HV37TDSXX:2:1433:2284:4225 chr21 40182751 N chr21 40183263 N DEL 10
A00404:156:HV37TDSXX:1:2470:28420:1454 chr21 40182849 N chr21 40183246 N DEL 7
A00404:155:HV27LDSXX:3:1245:21621:26005 chr21 40182851 N chr21 40183248 N DEL 7
A00297:158:HT275DSXX:1:1642:26160:14826 chr21 40182795 N chr21 40183279 N DEL 15
A00297:158:HT275DSXX:3:2408:14118:2519 chr21 40182795 N chr21 40183279 N DEL 13
A00404:156:HV37TDSXX:4:2208:17833:17190 chr21 40182795 N chr21 40183279 N DEL 5
A00297:158:HT275DSXX:1:1339:31684:15969 chr21 40182711 N chr21 40183280 N DEL 5
A00404:156:HV37TDSXX:4:2539:17879:10817 chr5 139453702 N chr5 139453884 N DEL 5
A00297:158:HT275DSXX:4:1421:26124:7874 chr5 139453702 N chr5 139453894 N DEL 2
A00404:156:HV37TDSXX:3:2309:11749:17394 chr5 139453712 N chr5 139453980 N DEL 15
A00404:155:HV27LDSXX:1:2430:22345:25097 chr5 139453702 N chr5 139453991 N DEL 5
A00404:156:HV37TDSXX:3:2658:2338:14591 chr5 139453710 N chr5 139454011 N DEL 5
A00404:155:HV27LDSXX:2:1261:5593:10488 chr5 139453702 N chr5 139454087 N DEL 5
A00404:156:HV37TDSXX:2:1337:25735:9768 chr5 139453704 N chr5 139454226 N DEL 5
A00404:156:HV37TDSXX:2:2275:23601:14967 chr5 139453702 N chr5 139454263 N DEL 5
A00297:158:HT275DSXX:1:2102:28185:26537 chr5 139453702 N chr5 139454329 N DEL 5
A00404:156:HV37TDSXX:4:2631:4698:5963 chr5 139453712 N chr5 139454429 N DEL 5
A00404:156:HV37TDSXX:3:2169:28131:17174 chr5 139453703 N chr5 139454580 N DEL 8
A00297:158:HT275DSXX:1:2363:6867:16485 chr5 139453709 N chr5 139454614 N DEL 5
A00404:155:HV27LDSXX:4:1150:32271:1329 chr5 139453702 N chr5 139454613 N DEL 5
A00404:156:HV37TDSXX:1:1474:31792:34601 chr5 139453704 N chr5 139454631 N DEL 5
A00404:156:HV37TDSXX:4:1358:22254:31234 chr5 139453706 N chr5 139454646 N DEL 10
A00404:156:HV37TDSXX:1:1178:2763:34272 chr5 139453707 N chr5 139454661 N DEL 5
A00404:156:HV37TDSXX:3:2234:28863:13150 chr7 16732542 N chr7 16732595 N DEL 4
A00297:158:HT275DSXX:3:2376:10149:31751 chr10 46526238 N chr10 46526458 N DUP 1
A00404:155:HV27LDSXX:2:2168:11776:35008 chr10 46526238 N chr10 46526458 N DUP 1
A00297:158:HT275DSXX:4:1417:18873:8187 chr10 46526237 N chr10 46526536 N DUP 1
A00404:156:HV37TDSXX:4:2331:8675:1548 chr10 46526237 N chr10 46526536 N DUP 1
A00404:156:HV37TDSXX:2:1216:3848:32612 chr10 46526460 N chr10 46526583 N DUP 2
A00404:155:HV27LDSXX:1:2544:2293:6840 chr10 46526460 N chr10 46526583 N DUP 3
A00297:158:HT275DSXX:2:1148:15157:19570 chr5 173203619 N chr5 173203670 N DEL 12
A00297:158:HT275DSXX:2:2642:12156:20635 chr5 173203611 N chr5 173203670 N DEL 5
A00297:158:HT275DSXX:2:2642:12255:20462 chr5 173203611 N chr5 173203670 N DEL 5
A00297:158:HT275DSXX:2:2474:17409:31172 chr5 173203607 N chr5 173203670 N DEL 5
A00297:158:HT275DSXX:4:2615:27444:21559 chr5 173203603 N chr5 173203670 N DEL 5
A00297:158:HT275DSXX:1:1370:22408:35822 chr5 173203601 N chr5 173203672 N DEL 5
A00297:158:HT275DSXX:3:1507:4463:5525 chr9 137739630 N chr9 137739760 N DEL 10
A00297:158:HT275DSXX:4:2143:15998:7874 chr9 137739635 N chr9 137739722 N DEL 5
A00404:156:HV37TDSXX:1:1149:12147:10880 chr9 137739635 N chr9 137739722 N DEL 5
A00404:156:HV37TDSXX:4:1508:19253:13761 chr9 137739606 N chr9 137739736 N DEL 1
A00297:158:HT275DSXX:3:1507:4463:5525 chr9 137739601 N chr9 137739774 N DEL 4
A00297:158:HT275DSXX:1:2427:7374:4617 chr19 56873912 N chr19 56873968 N DEL 11
A00404:155:HV27LDSXX:3:2171:2799:11287 chr19 56873912 N chr19 56873968 N DEL 11
A00404:155:HV27LDSXX:3:2458:26992:21339 chr19 56873912 N chr19 56873968 N DEL 11
A00404:155:HV27LDSXX:3:2114:14841:13322 chr19 56873912 N chr19 56873968 N DEL 11
A00404:156:HV37TDSXX:2:1142:15772:7858 chr19 56873912 N chr19 56873968 N DEL 11
A00404:156:HV37TDSXX:2:1142:16125:8124 chr19 56873912 N chr19 56873968 N DEL 11
A00404:156:HV37TDSXX:3:2577:16080:1658 chr19 56873912 N chr19 56873970 N DEL 13
A00404:156:HV37TDSXX:4:2611:15076:27477 chr19 56873912 N chr19 56873968 N DEL 11
A00404:155:HV27LDSXX:4:2312:11153:17738 chr19 56873962 N chr19 56874075 N DUP 18
A00297:158:HT275DSXX:4:2547:27480:17237 chr19 56873966 N chr19 56874079 N DUP 13
A00404:156:HV37TDSXX:1:1250:9778:20650 chr19 56874019 N chr19 56874091 N DUP 18
A00404:155:HV27LDSXX:2:2167:22670:33771 chr19 56873965 N chr19 56874060 N DEL 13
A00404:156:HV37TDSXX:1:1114:18665:14465 chr19 56873965 N chr19 56874060 N DEL 13
A00404:155:HV27LDSXX:4:2661:5629:32878 chr19 56873977 N chr19 56874074 N DEL 1
A00297:158:HT275DSXX:2:1637:14931:12665 chr19 56873981 N chr19 56874102 N DEL 5
A00404:155:HV27LDSXX:2:1126:1777:36135 chr19 56873981 N chr19 56874102 N DEL 5
A00404:155:HV27LDSXX:2:2123:30825:32393 chr19 56873977 N chr19 56874102 N DEL 5
A00404:155:HV27LDSXX:3:2140:12852:19366 chr19 56873981 N chr19 56874155 N DEL 14
A00404:156:HV37TDSXX:4:2338:25789:20228 chr16 24115336 N chr16 24115407 N DUP 5
A00404:156:HV37TDSXX:4:2409:21594:11490 chr6 31045224 N chr6 31045314 N DEL 4
A00404:155:HV27LDSXX:2:1628:5593:28808 chr6 31045224 N chr6 31045314 N DEL 8
A00404:155:HV27LDSXX:2:1628:7600:25426 chr6 31045224 N chr6 31045314 N DEL 8
A00404:155:HV27LDSXX:2:1628:4237:29465 chr6 31045224 N chr6 31045314 N DEL 10
A00297:158:HT275DSXX:3:2537:32145:31704 chr6 31045224 N chr6 31045314 N DEL 20
A00404:156:HV37TDSXX:3:1449:13286:24345 chr6 31045224 N chr6 31045314 N DEL 19
A00297:158:HT275DSXX:4:2117:11966:36714 chr6 31045224 N chr6 31045314 N DEL 10
A00404:156:HV37TDSXX:3:2118:4915:1172 chr6 31045224 N chr6 31045314 N DEL 10
A00297:158:HT275DSXX:1:1621:18502:1125 chr6 31045227 N chr6 31045317 N DEL 10
A00404:155:HV27LDSXX:2:1417:15980:5713 chr9 135177623 N chr9 135177747 N DEL 5
A00404:156:HV37TDSXX:1:2456:12870:3051 chr9 135177623 N chr9 135177747 N DEL 8
A00404:156:HV37TDSXX:1:1553:27977:1689 chr9 135177623 N chr9 135177747 N DEL 10
A00404:156:HV37TDSXX:1:1168:27371:9596 chr9 135177623 N chr9 135177747 N DEL 10
A00404:156:HV37TDSXX:1:2561:13078:5353 chr9 135177580 N chr9 135177662 N DUP 10
A00297:158:HT275DSXX:4:2201:21866:4726 chr9 135177580 N chr9 135177662 N DUP 10
A00404:156:HV37TDSXX:3:1236:30110:36573 chr9 135177580 N chr9 135177662 N DUP 10
A00404:156:HV37TDSXX:3:2273:16423:1783 chr9 135177653 N chr9 135178106 N DEL 5
A00404:155:HV27LDSXX:1:1531:29921:8093 chr9 135177653 N chr9 135178106 N DEL 5
A00404:156:HV37TDSXX:4:2557:23149:15875 chr9 135177653 N chr9 135178106 N DEL 5
A00297:158:HT275DSXX:1:1113:22978:31829 chr9 135177736 N chr9 135177817 N DUP 5
A00404:156:HV37TDSXX:2:1240:14163:19570 chr9 135177951 N chr9 135178075 N DEL 14
A00404:156:HV37TDSXX:2:2569:7093:18818 chr9 135177664 N chr9 135177951 N DUP 5
A00297:158:HT275DSXX:3:2434:7265:22153 chr9 135177664 N chr9 135177951 N DUP 5
A00297:158:HT275DSXX:1:1652:26756:18145 chr9 135177664 N chr9 135177951 N DUP 5
A00404:156:HV37TDSXX:2:1202:10990:34397 chr9 135177664 N chr9 135177951 N DUP 5
A00404:156:HV37TDSXX:3:2302:6334:30405 chr9 135177664 N chr9 135177951 N DUP 5
A00404:155:HV27LDSXX:3:2472:18801:1078 chr9 135177664 N chr9 135177951 N DUP 5
A00404:156:HV37TDSXX:1:1458:13810:31735 chr9 135177664 N chr9 135177951 N DUP 5
A00404:155:HV27LDSXX:1:2212:14082:9251 chr9 135177664 N chr9 135177951 N DUP 5
A00297:158:HT275DSXX:2:2416:20573:31923 chr9 135177664 N chr9 135177951 N DUP 5
A00404:155:HV27LDSXX:1:1164:22923:4679 chr9 135177624 N chr9 135177952 N DUP 5
A00404:155:HV27LDSXX:3:2444:26901:27445 chr9 135177626 N chr9 135177954 N DUP 5
A00297:158:HT275DSXX:1:1220:11984:6496 chr9 135177608 N chr9 135177980 N DEL 5
A00297:158:HT275DSXX:4:2201:21866:4726 chr9 135177619 N chr9 135177991 N DEL 4
A00404:156:HV37TDSXX:1:2561:13078:5353 chr9 135177792 N chr9 135177999 N DEL 7
A00297:158:HT275DSXX:4:2522:20347:26459 chr3 101551638 N chr3 101552017 N DEL 2
A00404:155:HV27LDSXX:2:2136:6081:24580 chr22 31336673 N chr22 31336979 N DEL 16
A00404:155:HV27LDSXX:2:1228:20491:7420 chr22 31336809 N chr22 31336979 N DEL 42
A00297:158:HT275DSXX:1:2353:7365:34788 chr1 232262701 N chr1 232262779 N DEL 4
A00297:158:HT275DSXX:2:1626:14271:6104 chr17 65971640 N chr17 65971742 N DUP 4
A00404:156:HV37TDSXX:3:2140:4056:6825 chr15 71670450 N chr15 71670866 N DEL 20
A00404:155:HV27LDSXX:3:1239:6253:5243 chr15 71670616 N chr15 71671031 N DUP 5
A00404:156:HV37TDSXX:3:1411:1714:18709 chr15 71670337 N chr15 71670754 N DEL 15
A00297:158:HT275DSXX:4:2443:24216:4225 chr15 71670518 N chr15 71670932 N DUP 1
A00404:155:HV27LDSXX:1:1530:23276:9549 chr15 71670450 N chr15 71670866 N DEL 13
A00404:155:HV27LDSXX:1:1530:23276:9549 chr15 71670518 N chr15 71670932 N DUP 6
A00404:156:HV37TDSXX:4:2225:32380:14387 chr15 71670564 N chr15 71670981 N DEL 11
A00404:156:HV37TDSXX:4:2225:32380:14387 chr15 71670564 N chr15 71670981 N DEL 11
A00404:155:HV27LDSXX:3:1640:21802:24471 chr15 71670564 N chr15 71670981 N DEL 6
A00404:156:HV37TDSXX:1:1306:9670:16078 chr15 71670564 N chr15 71670981 N DEL 6
A00404:156:HV37TDSXX:3:2659:26585:7639 chr15 71670564 N chr15 71670981 N DEL 6
A00404:156:HV37TDSXX:3:2659:26729:6981 chr15 71670564 N chr15 71670981 N DEL 6
A00404:156:HV37TDSXX:2:2151:12463:10958 chr15 71670590 N chr15 71671007 N DEL 4
A00297:158:HT275DSXX:1:1564:31340:11866 chr15 71670564 N chr15 71670981 N DEL 6
A00297:158:HT275DSXX:1:1129:21477:17957 chr15 71670566 N chr15 71670983 N DEL 6
A00404:156:HV37TDSXX:4:1530:30056:4194 chr15 71670578 N chr15 71670995 N DEL 1
A00404:155:HV27LDSXX:3:2235:11957:27211 chr8 10672488 N chr8 10672551 N DEL 2
A00404:155:HV27LDSXX:2:1305:19199:26381 chr3 175670557 N chr3 175670630 N DUP 11
A00404:156:HV37TDSXX:4:2621:25807:4038 chr3 175670557 N chr3 175670630 N DUP 11
A00297:158:HT275DSXX:2:1427:3450:9001 chr3 175670557 N chr3 175670630 N DUP 11
A00404:155:HV27LDSXX:4:1168:3125:6120 chr3 175670557 N chr3 175670630 N DUP 11
A00404:155:HV27LDSXX:4:1168:3152:5979 chr3 175670557 N chr3 175670630 N DUP 11
A00404:156:HV37TDSXX:4:1239:26802:8609 chr3 175670557 N chr3 175670630 N DUP 12
A00404:155:HV27LDSXX:2:1442:4869:32910 chr3 175670557 N chr3 175670630 N DUP 15
A00404:155:HV27LDSXX:1:1675:13494:17221 chr3 175670557 N chr3 175670630 N DUP 18
A00404:155:HV27LDSXX:4:2538:8386:24721 chr3 175670557 N chr3 175670630 N DUP 18
A00404:155:HV27LDSXX:2:1346:4282:14293 chr3 175670588 N chr3 175670674 N DEL 3
A00404:155:HV27LDSXX:3:1543:13349:24111 chr5 166683336 N chr5 166683401 N DUP 12
A00297:158:HT275DSXX:1:1606:2121:29027 chr5 166683327 N chr5 166683456 N DUP 22
A00404:155:HV27LDSXX:1:2375:18837:21621 chr5 166683335 N chr5 166683434 N DUP 14
A00404:156:HV37TDSXX:1:1569:18964:25692 chr5 166683335 N chr5 166683434 N DUP 17
A00404:155:HV27LDSXX:3:2471:25545:33458 chr5 166683327 N chr5 166683456 N DUP 28
A00404:155:HV27LDSXX:1:1518:26223:7263 chr5 166683378 N chr5 166683456 N DUP 19
A00297:158:HT275DSXX:2:1208:25672:12383 chr5 166683378 N chr5 166683456 N DUP 18
A00404:156:HV37TDSXX:4:2541:17418:26616 chr2 12627737 N chr2 12627800 N DEL 5
A00297:158:HT275DSXX:4:2616:32172:18380 chr7 55402587 N chr7 55402713 N DUP 5
A00404:156:HV37TDSXX:2:1304:1741:5948 chr7 55402582 N chr7 55402852 N DEL 13
A00297:158:HT275DSXX:3:2418:24677:32800 chr19 32746933 N chr19 32747212 N DEL 1
A00297:158:HT275DSXX:2:1278:26286:8281 chr19 32746843 N chr19 32747128 N DUP 4
A00404:155:HV27LDSXX:4:2338:19542:14168 chr19 32746954 N chr19 32747185 N DEL 5
A00404:156:HV37TDSXX:1:2130:8495:25848 chr19 32746858 N chr19 32747047 N DUP 5
A00297:158:HT275DSXX:2:1278:26286:8281 chr19 32746852 N chr19 32747263 N DUP 4
A00404:155:HV27LDSXX:3:1137:7473:34632 chr6 1544420 N chr6 1544501 N DEL 7
A00404:156:HV37TDSXX:2:1622:8467:32189 chr12 132619261 N chr12 132619380 N DEL 11
A00297:158:HT275DSXX:3:1618:15646:31970 chr12 132619335 N chr12 132619434 N DEL 18
A00404:155:HV27LDSXX:1:1201:2139:29872 chr12 132619237 N chr12 132619452 N DEL 3
A00404:156:HV37TDSXX:2:2677:6442:21950 chr12 12413824 N chr12 12414225 N DEL 5
A00404:156:HV37TDSXX:1:1427:18466:25989 chr12 12413835 N chr12 12414061 N DEL 5
A00297:158:HT275DSXX:4:2474:22941:9251 chr12 12413872 N chr12 12413951 N DEL 11
A00404:156:HV37TDSXX:4:2275:30951:32706 chr12 12413876 N chr12 12414275 N DUP 5
A00297:158:HT275DSXX:4:2520:17173:16016 chr12 12414047 N chr12 12414223 N DEL 5
A00404:155:HV27LDSXX:3:2526:21775:16845 chr12 12413976 N chr12 12414073 N DUP 5
A00297:158:HT275DSXX:4:1620:3079:24392 chr12 12413843 N chr12 12414195 N DEL 1
A00404:156:HV37TDSXX:2:1578:15537:2879 chr12 12414014 N chr12 12414239 N DEL 2
A00404:155:HV27LDSXX:3:1139:15754:2002 chr12 12413898 N chr12 12414396 N DUP 5
A00297:158:HT275DSXX:2:1205:7636:2973 chr12 12414304 N chr12 12414403 N DEL 22
A00404:156:HV37TDSXX:4:2569:29378:13855 chr12 12413994 N chr12 12414367 N DEL 5
A00404:155:HV27LDSXX:3:1139:15754:2002 chr12 12413997 N chr12 12414269 N DUP 5
A00297:158:HT275DSXX:2:2328:5520:20760 chr12 12413856 N chr12 12414532 N DEL 2
A00404:155:HV27LDSXX:4:2319:16857:33442 chr12 12414011 N chr12 12414560 N DEL 5
A00404:156:HV37TDSXX:2:1655:5493:10128 chr12 12414011 N chr12 12414560 N DEL 5
A00404:156:HV37TDSXX:4:1162:8052:6386 chr12 12414232 N chr12 12414682 N DUP 5
A00404:156:HV37TDSXX:4:1678:8919:27430 chr12 12414232 N chr12 12414682 N DUP 5
A00404:156:HV37TDSXX:4:2678:9652:34679 chr12 12414232 N chr12 12414682 N DUP 5
A00404:155:HV27LDSXX:1:2442:32904:16172 chr9 60526789 N chr9 60526933 N DUP 5
A00404:155:HV27LDSXX:2:2347:1642:12696 chr9 60526940 N chr9 60527035 N DUP 5
A00404:156:HV37TDSXX:3:2649:26169:30812 chr9 60526915 N chr9 60527058 N DUP 4
A00297:158:HT275DSXX:3:2129:17526:5384 chr9 60526915 N chr9 60527058 N DUP 4
A00404:155:HV27LDSXX:1:2212:19642:2159 chr9 60526940 N chr9 60527035 N DUP 5
A00404:156:HV37TDSXX:2:2255:25726:14262 chr9 60526917 N chr9 60527060 N DUP 2
A00404:155:HV27LDSXX:2:2578:9471:3333 chr19 6429233 N chr19 6429295 N DEL 3
A00404:156:HV37TDSXX:1:2156:10664:30044 chr19 6429180 N chr19 6429247 N DUP 7
A00297:158:HT275DSXX:2:1653:28185:10066 chr19 6429180 N chr19 6429247 N DUP 14
A00404:156:HV37TDSXX:3:1325:28167:12884 chr19 6429180 N chr19 6429247 N DUP 15
A00404:156:HV37TDSXX:3:1325:28691:12477 chr19 6429180 N chr19 6429247 N DUP 15
A00404:155:HV27LDSXX:4:1308:32615:18803 chr19 6429217 N chr19 6429299 N DEL 10
A00404:155:HV27LDSXX:1:1437:26485:5744 chr19 6429222 N chr19 6429326 N DEL 19
A00404:155:HV27LDSXX:1:2628:20862:21277 chr12 10027783 N chr12 10027844 N DUP 2
A00297:158:HT275DSXX:2:1637:9408:27618 chr9 121090159 N chr9 121090221 N DUP 4
A00404:156:HV37TDSXX:4:1113:18331:7028 chr10 108548642 N chr10 108548728 N DEL 5
A00297:158:HT275DSXX:2:2162:19587:33254 chr12 110144513 N chr12 110144645 N DUP 5
A00297:158:HT275DSXX:3:2676:25916:4445 chr12 110144513 N chr12 110144645 N DUP 5
A00297:158:HT275DSXX:4:1534:26386:8766 chr22 31265094 N chr22 31265402 N DEL 9
A00297:158:HT275DSXX:4:1162:20835:26303 chr22 31265519 N chr22 31265691 N DEL 7
A00297:158:HT275DSXX:2:1631:5385:18584 chr3 83105122 N chr3 83105229 N DUP 5
A00404:155:HV27LDSXX:2:1120:4806:5963 chr10 71432436 N chr10 71432514 N DEL 2
A00404:155:HV27LDSXX:3:1438:3712:7044 chr10 71432436 N chr10 71432514 N DEL 2
A00297:158:HT275DSXX:4:1316:18087:22232 chr10 71432363 N chr10 71432571 N DEL 2
A00297:158:HT275DSXX:4:1120:20853:15092 chr5 44440423 N chr5 44440531 N DEL 4
A00404:156:HV37TDSXX:4:1248:24288:3505 chr1 153668900 N chr1 153668955 N DUP 5
A00404:156:HV37TDSXX:1:2224:12572:19570 chr12 34211799 N chr12 34212005 N DEL 9
A00404:156:HV37TDSXX:1:1377:26738:2394 chr12 34211728 N chr12 34211934 N DEL 2
A00297:158:HT275DSXX:1:2355:13105:26976 chr12 34211857 N chr12 34212063 N DEL 8
A00297:158:HT275DSXX:2:2414:24623:26318 chr5 31766881 N chr5 31767180 N DEL 6
A00404:155:HV27LDSXX:1:2313:28103:4194 chr22 10571950 N chr22 10572199 N DUP 11
A00404:155:HV27LDSXX:2:2308:12002:32456 chr22 10571953 N chr22 10572058 N DUP 6
A00297:158:HT275DSXX:4:2276:7030:10473 chr5 94533379 N chr5 94533677 N DEL 5
A00404:156:HV37TDSXX:4:1507:11360:23234 chr5 94533154 N chr5 94533453 N DEL 10
A00297:158:HT275DSXX:4:2525:14262:25410 chr2 241052687 N chr2 241052738 N DUP 2
A00404:156:HV37TDSXX:1:1260:14271:31093 chr2 241052687 N chr2 241052738 N DUP 5
A00297:158:HT275DSXX:2:2601:14886:18317 chr2 241052626 N chr2 241052680 N DEL 5
A00404:155:HV27LDSXX:1:1368:4010:18552 chr2 241052793 N chr2 241053012 N DEL 13
A00404:156:HV37TDSXX:1:2664:5303:5916 chr2 241052693 N chr2 241052964 N DEL 4
A00404:156:HV37TDSXX:1:1167:23746:13182 chr11 59632741 N chr11 59632812 N DUP 6
A00404:155:HV27LDSXX:4:2250:23845:27853 chr11 59632765 N chr11 59632822 N DUP 9
A00404:155:HV27LDSXX:1:1145:2175:28119 chr11 59632751 N chr11 59632816 N DEL 8
A00297:158:HT275DSXX:4:1513:27462:13009 chr11 59632778 N chr11 59632847 N DEL 3
A00404:155:HV27LDSXX:3:2455:17445:18239 chr11 59632748 N chr11 59632904 N DEL 8
A00404:155:HV27LDSXX:3:2213:1416:14873 chr12 132313247 N chr12 132313729 N DEL 5
A00297:158:HT275DSXX:2:1374:28076:18552 chr12 132313326 N chr12 132313415 N DEL 5
A00404:155:HV27LDSXX:3:2239:15971:11177 chr12 132313275 N chr12 132313813 N DEL 13
A00297:158:HT275DSXX:4:2434:17535:2895 chr12 132314150 N chr12 132314211 N DEL 40
A00297:158:HT275DSXX:4:2449:30472:30029 chr12 132313406 N chr12 132314239 N DEL 5
A00404:155:HV27LDSXX:4:2345:23493:25300 chr20 46507299 N chr20 46507411 N DUP 5
A00404:155:HV27LDSXX:4:1521:26775:3803 chr20 24957250 N chr20 24957318 N DUP 5
A00404:156:HV37TDSXX:2:2265:29577:12289 chr20 24957254 N chr20 24957322 N DUP 1
A00297:158:HT275DSXX:4:2135:9706:3333 chr11 22316688 N chr11 22316815 N DEL 42
A00297:158:HT275DSXX:1:2576:5981:33364 chr7 6742210 N chr7 6742342 N DUP 5
A00297:158:HT275DSXX:4:1513:8748:12665 chr21 38622584 N chr21 38623092 N DUP 3
A00404:155:HV27LDSXX:2:1469:32560:31140 chr21 38622582 N chr21 38622668 N DUP 5
A00404:155:HV27LDSXX:1:2155:29903:17018 chr21 10801044 N chr21 10801387 N DUP 6
A00404:155:HV27LDSXX:1:1643:11080:1548 chr21 10801119 N chr21 10801636 N DEL 5
A00404:156:HV37TDSXX:2:1120:14742:8797 chr21 10800812 N chr21 10801499 N DUP 1
A00297:158:HT275DSXX:1:1209:3784:13213 chr21 10800659 N chr21 10801348 N DEL 3
A00404:155:HV27LDSXX:3:1421:12038:27633 chr21 10801045 N chr21 10801388 N DUP 5
A00297:158:HT275DSXX:1:1267:19931:20353 chr21 10800773 N chr21 10801637 N DEL 8
A00404:155:HV27LDSXX:4:1149:10917:3396 chr21 10801102 N chr21 10801617 N DUP 3
A00404:155:HV27LDSXX:1:1610:25925:27038 chr21 10800773 N chr21 10801637 N DEL 8
A00404:155:HV27LDSXX:3:1515:27498:26537 chr21 10801023 N chr21 10801366 N DEL 13
A00404:156:HV37TDSXX:1:1371:25274:26663 chr21 10801046 N chr21 10801389 N DUP 5
A00404:156:HV37TDSXX:2:2224:30201:35884 chr21 10801038 N chr21 10801381 N DUP 10
A00297:158:HT275DSXX:1:1267:19877:20917 chr21 10800773 N chr21 10801637 N DEL 8
A00404:155:HV27LDSXX:1:1243:32289:4899 chr21 10801102 N chr21 10801617 N DUP 1
A00297:158:HT275DSXX:3:2138:19009:27649 chr21 10801211 N chr21 10801556 N DEL 2
A00297:158:HT275DSXX:2:1470:7410:8124 chr21 10800499 N chr21 10800842 N DEL 5
A00404:156:HV37TDSXX:4:1143:24279:30170 chr21 10801119 N chr21 10801636 N DEL 5
A00404:156:HV37TDSXX:3:2235:1651:15749 chr21 10800487 N chr21 10801347 N DEL 5
A00404:156:HV37TDSXX:3:2118:27959:35822 chr21 10801125 N chr21 10801298 N DEL 5
A00297:158:HT275DSXX:3:2603:25274:21057 chr21 10801102 N chr21 10801617 N DUP 3
A00297:158:HT275DSXX:2:1518:30960:19852 chr21 10801119 N chr21 10801636 N DEL 5
A00404:156:HV37TDSXX:2:1243:3531:13808 chr1 23767145 N chr1 23767450 N DEL 4
A00404:156:HV37TDSXX:4:1620:2663:31187 chr1 163628599 N chr1 163628655 N DEL 5
A00404:155:HV27LDSXX:2:2506:5195:22764 chr21 44948291 N chr21 44948514 N DEL 27
A00297:158:HT275DSXX:4:2364:10321:32487 chr21 44948329 N chr21 44948514 N DEL 33
A00404:156:HV37TDSXX:4:1453:7518:34209 chr21 44948335 N chr21 44948490 N DEL 6
A00297:158:HT275DSXX:1:1544:22272:13510 chr21 44948339 N chr21 44948524 N DEL 12
A00297:158:HT275DSXX:3:1602:30553:21496 chr16 30223204 N chr16 30223379 N DEL 9
A00404:155:HV27LDSXX:4:1126:9299:14434 chr16 30223189 N chr16 30223451 N DEL 12
A00404:155:HV27LDSXX:1:1544:2003:32518 chr6 40623320 N chr6 40623466 N DEL 5
A00404:155:HV27LDSXX:1:2445:30083:6715 chr6 40623320 N chr6 40623466 N DEL 5
A00404:155:HV27LDSXX:4:1560:1018:18223 chr6 40623320 N chr6 40623466 N DEL 5
A00404:156:HV37TDSXX:3:1409:30002:25864 chr6 40623516 N chr6 40623664 N DEL 11
A00297:158:HT275DSXX:1:2441:15103:7639 chr8 128118811 N chr8 128118937 N DUP 15
A00404:155:HV27LDSXX:3:2141:19470:26913 chr8 128118811 N chr8 128118888 N DUP 15
A00404:156:HV37TDSXX:1:1570:31720:27618 chr8 128118812 N chr8 128118889 N DUP 11
A00404:156:HV37TDSXX:4:2133:5339:21543 chr8 128118802 N chr8 128118928 N DUP 10
A00404:156:HV37TDSXX:1:1647:20057:8985 chr8 128118815 N chr8 128118941 N DUP 4
A00404:156:HV37TDSXX:2:2263:17616:2691 chr8 128118811 N chr8 128118937 N DUP 9
A00404:155:HV27LDSXX:2:2163:20582:16877 chr8 128118811 N chr8 128118937 N DUP 10
A00297:158:HT275DSXX:1:1517:14498:32049 chr8 128118887 N chr8 128119013 N DUP 5
A00297:158:HT275DSXX:2:2274:22128:15358 chr8 128118811 N chr8 128118937 N DUP 10
A00297:158:HT275DSXX:1:2341:22625:29810 chr8 116678652 N chr8 116678847 N DUP 3
A00297:158:HT275DSXX:3:1409:15447:6324 chr8 116678656 N chr8 116678851 N DUP 5
A00297:158:HT275DSXX:3:1618:25626:15468 chr18 3576744 N chr18 3577043 N DEL 35
A00404:156:HV37TDSXX:2:1514:26458:4664 chr20 46626441 N chr20 46626491 N DUP 4
A00404:155:HV27LDSXX:2:2508:14208:34334 chr6 158169491 N chr6 158169546 N DUP 27
A00404:156:HV37TDSXX:4:2304:17833:19006 chr6 158169510 N chr6 158169894 N DUP 17
A00404:156:HV37TDSXX:3:1147:29396:19022 chr6 158169625 N chr6 158169706 N DEL 18
A00404:155:HV27LDSXX:3:2615:15393:23829 chr6 158169665 N chr6 158169817 N DEL 22
A00404:156:HV37TDSXX:3:1545:23701:33708 chr6 158169875 N chr6 158169935 N DUP 30
A00297:158:HT275DSXX:3:1672:4182:13432 chr6 158169836 N chr6 158169887 N DUP 28
A00297:158:HT275DSXX:4:1204:6027:16595 chr6 158169804 N chr6 158169942 N DUP 25
A00404:155:HV27LDSXX:3:2442:28004:33959 chr6 158169843 N chr6 158169957 N DUP 31
A00404:156:HV37TDSXX:4:2329:24975:15342 chr6 158169836 N chr6 158169887 N DUP 29
A00404:155:HV27LDSXX:4:1568:16559:17049 chr6 158169586 N chr6 158169836 N DEL 16
A00297:158:HT275DSXX:2:2231:1805:27602 chr6 158169651 N chr6 158169935 N DUP 15
A00404:155:HV27LDSXX:1:2155:31810:33818 chr6 158169836 N chr6 158169887 N DUP 40
A00297:158:HT275DSXX:3:1141:27299:13260 chr6 158169875 N chr6 158169935 N DUP 25
A00404:156:HV37TDSXX:1:1466:12346:6872 chr6 158169748 N chr6 158169922 N DEL 23
A00297:158:HT275DSXX:2:1634:9552:13589 chr6 158169827 N chr6 158169962 N DEL 2
A00404:156:HV37TDSXX:2:1336:32895:7388 chr6 158169587 N chr6 158169922 N DEL 15
A00404:156:HV37TDSXX:4:2152:24614:22639 chr6 158169587 N chr6 158169922 N DEL 12
A00404:155:HV27LDSXX:4:2518:7120:9095 chr6 158169588 N chr6 158169923 N DEL 11
A00404:155:HV27LDSXX:3:2615:15393:23829 chr6 158169563 N chr6 158169926 N DEL 10
A00404:156:HV37TDSXX:3:1237:25789:6950 chr5 78363270 N chr5 78363588 N DEL 3
A00404:155:HV27LDSXX:1:1477:31828:11772 chr1 53096719 N chr1 53097128 N DEL 2
A00404:155:HV27LDSXX:2:2506:4381:8359 chr1 53097555 N chr1 53097646 N DEL 3
A00404:156:HV37TDSXX:3:2329:3875:34601 chr1 53097525 N chr1 53097593 N DUP 5
A00297:158:HT275DSXX:3:1324:10710:16532 chr1 53097600 N chr1 53097666 N DUP 5
A00297:158:HT275DSXX:1:1637:24749:12070 chr1 53097624 N chr1 53097826 N DUP 4
A00404:155:HV27LDSXX:1:1414:4562:32816 chr1 53097132 N chr1 53097828 N DUP 5
A00404:155:HV27LDSXX:1:1414:5520:33004 chr1 53097132 N chr1 53097828 N DUP 5
A00404:156:HV37TDSXX:1:1114:4463:9690 chr1 53097132 N chr1 53097828 N DUP 5
A00404:156:HV37TDSXX:2:2561:20781:24455 chr1 53096716 N chr1 53097845 N DEL 5
A00404:156:HV37TDSXX:2:1435:1452:5822 chr1 53096716 N chr1 53097845 N DEL 5
A00404:156:HV37TDSXX:4:1218:24551:25066 chr1 53096716 N chr1 53097845 N DEL 5
A00297:158:HT275DSXX:2:2417:1985:29011 chr1 53097154 N chr1 53097852 N DEL 5
A00404:155:HV27LDSXX:2:1470:32334:26647 chr1 53097042 N chr1 53098127 N DUP 1
A00404:155:HV27LDSXX:2:2470:30834:20102 chr1 53097042 N chr1 53098127 N DUP 1
A00404:156:HV37TDSXX:2:1528:14398:28588 chr7 89959262 N chr7 89959318 N DUP 12
A00404:155:HV27LDSXX:4:2575:27706:10050 chr7 89959262 N chr7 89959318 N DUP 16
A00404:156:HV37TDSXX:2:1131:19117:2127 chr7 89959262 N chr7 89959318 N DUP 24
A00404:155:HV27LDSXX:2:1107:28574:32377 chr7 89959311 N chr7 89959363 N DUP 28
A00404:155:HV27LDSXX:1:2214:21866:33974 chr7 89959311 N chr7 89959363 N DUP 26
A00404:156:HV37TDSXX:1:1509:23014:8500 chr7 89959311 N chr7 89959363 N DUP 26
A00404:156:HV37TDSXX:4:1637:2094:6183 chr7 89959311 N chr7 89959363 N DUP 16
A00297:158:HT275DSXX:2:2345:1768:35368 chr1 99112050 N chr1 99112183 N DUP 7
A00297:158:HT275DSXX:1:1110:22941:11068 chr16 20622114 N chr16 20622240 N DEL 12
A00297:158:HT275DSXX:3:2508:20528:25864 chr1 8501187 N chr1 8501648 N DUP 12
A00297:158:HT275DSXX:1:2467:28176:25708 chr1 8501294 N chr1 8501635 N DUP 12
A00404:156:HV37TDSXX:3:2656:32922:32925 chr1 8501294 N chr1 8501635 N DUP 14
A00297:158:HT275DSXX:1:2155:5412:8641 chr1 8501294 N chr1 8501635 N DUP 10
A00404:155:HV27LDSXX:3:1577:14977:9768 chr1 8501232 N chr1 8501904 N DUP 5
A00297:158:HT275DSXX:3:2153:31412:24612 chr1 8501294 N chr1 8501635 N DUP 10
A00297:158:HT275DSXX:1:1678:8486:31751 chr1 8501294 N chr1 8501635 N DUP 10
A00297:158:HT275DSXX:1:2127:10104:32957 chr1 8501294 N chr1 8501635 N DUP 10
A00404:155:HV27LDSXX:4:2658:17653:18881 chr1 8501321 N chr1 8501622 N DEL 6
A00404:155:HV27LDSXX:2:2420:12057:5932 chr1 8501294 N chr1 8501635 N DUP 5
A00404:155:HV27LDSXX:4:2233:11143:18630 chr1 8501321 N chr1 8501622 N DEL 27
A00404:156:HV37TDSXX:3:1556:1624:6308 chr1 8501294 N chr1 8501635 N DUP 5
A00404:155:HV27LDSXX:3:2248:21106:15154 chr1 8501294 N chr1 8501635 N DUP 5
A00297:158:HT275DSXX:4:1264:5222:33395 chr1 8501381 N chr1 8501555 N DEL 1
A00404:155:HV27LDSXX:2:1153:7265:21183 chr1 8501381 N chr1 8501555 N DEL 2
A00404:155:HV27LDSXX:1:1171:10493:2221 chr1 8501381 N chr1 8501555 N DEL 2
A00404:155:HV27LDSXX:4:1163:4209:27571 chr1 8501306 N chr1 8501473 N DUP 5
A00404:155:HV27LDSXX:4:1222:12816:7999 chr1 8501321 N chr1 8501622 N DEL 27
A00297:158:HT275DSXX:3:2648:24795:28213 chr1 8501385 N chr1 8501669 N DEL 1
A00404:155:HV27LDSXX:3:1342:13367:23610 chr1 8501385 N chr1 8501669 N DEL 1
A00404:156:HV37TDSXX:3:1119:15447:7138 chr1 8501493 N chr1 8501825 N DEL 5
A00404:155:HV27LDSXX:3:1468:2537:23234 chr1 8501294 N chr1 8501635 N DUP 8
A00404:156:HV37TDSXX:4:2118:29903:22122 chr1 8501331 N chr1 8501632 N DEL 5
A00404:155:HV27LDSXX:2:1506:30807:24095 chr1 8501202 N chr1 8501623 N DEL 14
A00404:156:HV37TDSXX:1:1246:20971:1172 chr1 8501717 N chr1 8501988 N DEL 14
A00404:156:HV37TDSXX:3:2137:23231:21245 chr1 8501641 N chr1 8501797 N DUP 7
A00404:155:HV27LDSXX:4:2511:17282:29888 chr1 8501641 N chr1 8501845 N DUP 2
A00404:156:HV37TDSXX:3:2653:30626:5995 chr1 8501641 N chr1 8501845 N DUP 5
A00297:158:HT275DSXX:4:1355:27001:8891 chr1 8501733 N chr1 8501828 N DUP 5
A00297:158:HT275DSXX:4:1240:16568:20572 chr1 8501177 N chr1 8501755 N DEL 5
A00404:156:HV37TDSXX:1:1456:8684:33724 chr1 8501733 N chr1 8501828 N DUP 10
A00297:158:HT275DSXX:1:2545:10176:26788 chr1 8501733 N chr1 8501828 N DUP 10
A00297:158:HT275DSXX:2:2652:7075:31407 chr1 8501798 N chr1 8501893 N DUP 5
A00297:158:HT275DSXX:4:2411:18521:9737 chr1 8501733 N chr1 8501828 N DUP 10
A00404:155:HV27LDSXX:1:2274:24071:4225 chr1 8501734 N chr1 8501829 N DUP 10
A00404:155:HV27LDSXX:4:1370:2338:4789 chr1 8501798 N chr1 8501893 N DUP 5
A00404:155:HV27LDSXX:1:1401:4707:6167 chr1 8501220 N chr1 8501798 N DEL 5
A00404:155:HV27LDSXX:2:2237:31458:14700 chr1 8501733 N chr1 8501828 N DUP 10
A00404:156:HV37TDSXX:3:2137:23231:21245 chr1 8501797 N chr1 8501894 N DEL 10
A00404:156:HV37TDSXX:1:2667:23384:26146 chr1 8501320 N chr1 8501874 N DEL 2
A00404:156:HV37TDSXX:2:1258:31458:2237 chr1 8501808 N chr1 8501905 N DEL 4
A00404:155:HV27LDSXX:3:2152:31141:35665 chr1 8501182 N chr1 8502030 N DUP 10
A00404:156:HV37TDSXX:1:2119:2799:29387 chr1 8501176 N chr1 8502076 N DUP 11
A00404:156:HV37TDSXX:4:2620:19714:36824 chr1 8501324 N chr1 8502052 N DUP 1
A00404:155:HV27LDSXX:1:2402:15890:19210 chr1 8501324 N chr1 8502052 N DUP 2
A00404:156:HV37TDSXX:3:2653:30626:5995 chr1 8501324 N chr1 8502052 N DUP 6
A00297:158:HT275DSXX:1:1143:5159:3537 chr2 238317204 N chr2 238317523 N DEL 14
A00404:156:HV37TDSXX:2:1238:18801:21652 chr21 44183901 N chr21 44183953 N DEL 1
A00404:155:HV27LDSXX:2:1334:28266:31219 chr21 44183863 N chr21 44184017 N DEL 3
A00404:156:HV37TDSXX:2:1533:21549:7279 chr6 124892640 N chr6 124892799 N DUP 1
A00404:155:HV27LDSXX:3:1641:18349:14575 chr6 124892640 N chr6 124892799 N DUP 3
A00297:158:HT275DSXX:4:1452:10122:25504 chr6 124892640 N chr6 124892799 N DUP 5
A00297:158:HT275DSXX:4:1452:10140:25504 chr6 124892640 N chr6 124892799 N DUP 5
A00404:155:HV27LDSXX:2:2204:28058:15170 chr6 124892640 N chr6 124892799 N DUP 5
A00404:155:HV27LDSXX:2:2257:15736:23672 chr6 124892640 N chr6 124892799 N DUP 5
A00404:155:HV27LDSXX:4:2474:19859:13839 chr6 124892640 N chr6 124892799 N DUP 5
A00404:155:HV27LDSXX:1:1443:31684:24612 chr6 124892675 N chr6 124892836 N DEL 5
A00404:156:HV37TDSXX:1:2608:30110:19946 chr6 124892679 N chr6 124892840 N DEL 5
A00404:156:HV37TDSXX:3:1547:31557:33004 chr6 124892681 N chr6 124892842 N DEL 4
A00404:156:HV37TDSXX:2:1533:21549:7279 chr6 124892703 N chr6 124892864 N DEL 5
A00404:155:HV27LDSXX:3:1303:17146:17848 chr10 133020968 N chr10 133021038 N DEL 31
A00297:158:HT275DSXX:3:1260:18249:31156 chr14 21427583 N chr14 21427766 N DUP 5
A00404:156:HV37TDSXX:1:1250:20627:14888 chr14 21427609 N chr14 21427745 N DUP 2
A00404:155:HV27LDSXX:4:1511:26747:8046 chr14 21427574 N chr14 21427712 N DEL 5
A00404:155:HV27LDSXX:2:1534:23204:20071 chr14 21427740 N chr14 21427875 N DEL 5
A00404:156:HV37TDSXX:1:1506:28131:2018 chr14 21427558 N chr14 21427964 N DEL 2
A00404:155:HV27LDSXX:2:2277:32615:5431 chr8 129702552 N chr8 129702669 N DUP 3
A00404:155:HV27LDSXX:2:1178:22733:2190 chr8 129702552 N chr8 129702669 N DUP 3
A00297:158:HT275DSXX:1:1533:1904:29966 chr8 129702583 N chr8 129702706 N DUP 17
A00404:156:HV37TDSXX:3:1572:10059:32690 chr8 129702552 N chr8 129702669 N DUP 8
A00404:155:HV27LDSXX:1:1231:24171:13166 chr8 129702583 N chr8 129702706 N DUP 17
A00404:156:HV37TDSXX:1:1604:30228:31704 chr8 129702524 N chr8 129702611 N DEL 15
A00404:155:HV27LDSXX:2:2277:32615:5431 chr8 129702583 N chr8 129702706 N DUP 26
A00297:158:HT275DSXX:2:2430:29026:28557 chr5 85946420 N chr5 85946471 N DEL 11
A00404:155:HV27LDSXX:2:1408:19235:33238 chr5 85946420 N chr5 85946471 N DEL 11
A00404:155:HV27LDSXX:2:1408:19795:33489 chr5 85946420 N chr5 85946471 N DEL 11
A00404:156:HV37TDSXX:1:2329:17029:27007 chr17 80492350 N chr17 80492617 N DEL 5
A00404:156:HV37TDSXX:4:1418:25229:32315 chr17 80492378 N chr17 80492586 N DUP 3
A00404:156:HV37TDSXX:2:2540:2808:32847 chr17 80492359 N chr17 80492602 N DEL 6
A00297:158:HT275DSXX:1:1666:10981:20008 chr1 52185876 N chr1 52186196 N DEL 4
A00404:155:HV27LDSXX:2:1215:2645:1251 chr2 94208548 N chr2 94208663 N DEL 7
A00297:158:HT275DSXX:1:1657:20871:30906 chr2 94208582 N chr2 94208661 N DEL 6
A00404:156:HV37TDSXX:1:1360:30770:35180 chr2 94208582 N chr2 94208661 N DEL 10
A00297:158:HT275DSXX:1:2570:26657:2816 chr2 94208582 N chr2 94208661 N DEL 14
A00404:156:HV37TDSXX:1:2551:14226:1172 chr2 94208548 N chr2 94208663 N DEL 28
A00404:156:HV37TDSXX:3:1527:3604:24330 chr2 94208582 N chr2 94208809 N DEL 28
A00404:155:HV27LDSXX:4:1311:19054:29011 chr2 94208582 N chr2 94208661 N DEL 38
A00404:155:HV27LDSXX:4:2543:24153:30170 chr2 94208661 N chr2 94208880 N DEL 3
A00404:156:HV37TDSXX:3:1527:3604:24330 chr2 94208583 N chr2 94208880 N DEL 47
A00404:155:HV27LDSXX:1:2528:31774:19382 chr2 94208648 N chr2 94208963 N DEL 23
A00404:155:HV27LDSXX:1:1532:6397:4742 chr2 94208679 N chr2 94208880 N DEL 12
A00404:155:HV27LDSXX:3:1570:5882:11209 chr2 94208580 N chr2 94208675 N DUP 2
A00297:158:HT275DSXX:2:1524:12183:12007 chr2 94208678 N chr2 94208809 N DEL 10
A00404:156:HV37TDSXX:1:2529:8097:12665 chr2 94208678 N chr2 94208809 N DEL 17
A00404:155:HV27LDSXX:1:2157:2528:11130 chr2 94208678 N chr2 94208809 N DEL 18
A00404:156:HV37TDSXX:1:1420:20428:13698 chr2 94208678 N chr2 94208809 N DEL 27
A00404:155:HV27LDSXX:1:2172:18945:27226 chr2 94208678 N chr2 94208809 N DEL 33
A00404:155:HV27LDSXX:4:2345:17210:33458 chr2 94208678 N chr2 94208809 N DEL 33
A00404:155:HV27LDSXX:4:1371:16975:32800 chr2 94208691 N chr2 94208742 N DUP 5
A00404:155:HV27LDSXX:3:1672:29369:12680 chr2 94208763 N chr2 94208904 N DEL 10
A00404:156:HV37TDSXX:2:2409:3170:22576 chr2 94208591 N chr2 94208696 N DEL 13
A00404:155:HV27LDSXX:1:2537:4508:32252 chr2 94208591 N chr2 94208696 N DEL 13
A00297:158:HT275DSXX:3:2107:20645:15201 chr2 94208670 N chr2 94208773 N DUP 5
A00404:156:HV37TDSXX:2:1519:5195:23234 chr2 94208661 N chr2 94208826 N DUP 6
A00404:156:HV37TDSXX:2:2266:15347:29637 chr2 94208661 N chr2 94208826 N DUP 6
A00404:156:HV37TDSXX:3:1170:6207:31626 chr2 94208678 N chr2 94208809 N DEL 16
A00404:156:HV37TDSXX:4:1548:16215:15233 chr2 94208678 N chr2 94208809 N DEL 22
A00297:158:HT275DSXX:2:2326:12906:35931 chr2 94208678 N chr2 94208809 N DEL 26
A00404:155:HV27LDSXX:1:2164:20754:23062 chr2 94208615 N chr2 94208790 N DEL 15
A00404:155:HV27LDSXX:4:2106:8567:11819 chr2 94208678 N chr2 94208809 N DEL 41
A00404:156:HV37TDSXX:2:2277:13593:33332 chr2 94208678 N chr2 94208809 N DEL 41
A00404:156:HV37TDSXX:1:2261:30192:20494 chr2 94208678 N chr2 94208809 N DEL 41
A00297:158:HT275DSXX:1:1310:12364:3176 chr2 94208680 N chr2 94208879 N DUP 6
A00404:155:HV27LDSXX:3:1123:30572:17926 chr2 94208678 N chr2 94208809 N DEL 41
A00297:158:HT275DSXX:2:1462:29008:18129 chr2 94208678 N chr2 94208809 N DEL 41
A00404:156:HV37TDSXX:3:1567:14588:17300 chr2 94208705 N chr2 94208854 N DEL 5
A00404:156:HV37TDSXX:3:1547:2401:11130 chr2 94208678 N chr2 94208809 N DEL 41
A00404:155:HV27LDSXX:3:2243:15067:35039 chr2 94208678 N chr2 94208809 N DEL 41
A00404:156:HV37TDSXX:2:1258:2691:28447 chr2 94208678 N chr2 94208809 N DEL 41
A00404:156:HV37TDSXX:3:1358:26160:22498 chr2 94208678 N chr2 94208809 N DEL 35
A00404:156:HV37TDSXX:1:2166:32461:36323 chr2 94208586 N chr2 94208813 N DEL 7
A00404:156:HV37TDSXX:2:1549:16215:7936 chr2 94208678 N chr2 94208809 N DEL 16
A00297:158:HT275DSXX:4:2515:7111:16532 chr2 94208573 N chr2 94208844 N DEL 26
A00404:155:HV27LDSXX:4:1371:16975:32800 chr2 94208830 N chr2 94208899 N DUP 10
A00404:156:HV37TDSXX:2:2465:28230:28432 chr2 94208705 N chr2 94208854 N DEL 5
A00404:156:HV37TDSXX:4:1318:7636:19413 chr2 94208847 N chr2 94208968 N DUP 5
A00404:155:HV27LDSXX:2:2272:21341:23296 chr2 94208588 N chr2 94208859 N DEL 5
A00404:156:HV37TDSXX:3:1547:2428:11146 chr2 94208687 N chr2 94208914 N DEL 41
A00404:155:HV27LDSXX:3:2175:27453:35321 chr2 94208891 N chr2 94208970 N DEL 18
A00404:155:HV27LDSXX:1:2604:29107:33708 chr2 94208897 N chr2 94208994 N DEL 23
A00404:156:HV37TDSXX:3:1247:11523:24111 chr2 94208863 N chr2 94208916 N DEL 13
A00404:155:HV27LDSXX:2:2571:20320:14450 chr2 94208564 N chr2 94208923 N DEL 6
A00404:156:HV37TDSXX:4:1569:7789:14888 chr2 94208679 N chr2 94208976 N DEL 43
A00404:156:HV37TDSXX:2:2237:21151:9752 chr2 94208891 N chr2 94208988 N DEL 3
A00297:158:HT275DSXX:1:2566:11324:29747 chr2 94208661 N chr2 94208976 N DEL 35
A00297:158:HT275DSXX:1:1508:4463:2644 chr2 94208921 N chr2 94208974 N DEL 5
A00404:155:HV27LDSXX:2:1527:6234:3239 chr2 94208618 N chr2 94208985 N DEL 8
A00404:155:HV27LDSXX:4:1643:19298:23703 chr2 94208674 N chr2 94208989 N DEL 2
A00404:155:HV27LDSXX:2:2324:29631:20776 chr10 93693630 N chr10 93693823 N DEL 8
A00404:156:HV37TDSXX:2:2269:32723:29230 chr10 93693636 N chr10 93693825 N DEL 4
A00297:158:HT275DSXX:3:2236:29505:34366 chr10 93693630 N chr10 93693823 N DEL 16
A00404:156:HV37TDSXX:2:1273:16947:9737 chr10 93693687 N chr10 93693817 N DUP 9
A00297:158:HT275DSXX:1:2519:6207:1564 chr10 93693659 N chr10 93693832 N DUP 13
A00404:156:HV37TDSXX:4:2609:7600:10676 chr10 93693673 N chr10 93693823 N DEL 18
A00297:158:HT275DSXX:3:2239:15745:35994 chr10 93693673 N chr10 93693823 N DEL 16
A00297:158:HT275DSXX:2:2220:22064:20353 chr10 3399597 N chr10 3399750 N DUP 5
A00404:156:HV37TDSXX:1:2172:19687:9502 chr10 3399612 N chr10 3399767 N DEL 5
A00404:156:HV37TDSXX:3:2150:29188:16376 chr18 53206222 N chr18 53206339 N DEL 5
A00297:158:HT275DSXX:3:1506:3992:31078 chr7 66865719 N chr7 66865787 N DEL 5
A00404:156:HV37TDSXX:3:1128:25735:8766 chr7 66865706 N chr7 66865772 N DUP 5
A00404:155:HV27LDSXX:3:1113:17029:13855 chr7 66865706 N chr7 66865772 N DUP 5
A00404:155:HV27LDSXX:4:2625:28429:17096 chr7 66865706 N chr7 66865772 N DUP 5
A00404:155:HV27LDSXX:4:2625:28709:18427 chr7 66865706 N chr7 66865772 N DUP 5
A00297:158:HT275DSXX:2:1247:18231:1908 chr7 66865721 N chr7 66865789 N DEL 5
A00297:158:HT275DSXX:2:2521:8024:37027 chr22 34578954 N chr22 34579079 N DEL 25
A00404:155:HV27LDSXX:3:1165:1054:28181 chr22 34578946 N chr22 34579013 N DEL 20
A00404:156:HV37TDSXX:3:2304:14488:2942 chr22 34578936 N chr22 34579054 N DEL 5
A00404:156:HV37TDSXX:1:1444:27697:12414 chr22 34578931 N chr22 34579049 N DEL 10
A00297:158:HT275DSXX:3:1211:20347:5572 chr1 46241361 N chr1 46241586 N DUP 5
A00404:155:HV27LDSXX:4:1302:26775:22028 chr1 46241588 N chr1 46241893 N DEL 10
A00297:158:HT275DSXX:3:2676:26313:3724 chr1 46241587 N chr1 46241713 N DUP 5
A00404:156:HV37TDSXX:1:2567:15203:19116 chr1 46241347 N chr1 46241698 N DUP 5
A00297:158:HT275DSXX:1:1658:1307:18912 chr1 46241634 N chr1 46241811 N DEL 7
A00297:158:HT275DSXX:2:2466:6090:23093 chr1 46241609 N chr1 46241914 N DEL 5
A00404:155:HV27LDSXX:2:1165:31358:36793 chr1 46241492 N chr1 46241716 N DUP 2
A00404:155:HV27LDSXX:1:2616:8431:11710 chr1 46241383 N chr1 46241610 N DEL 5
A00404:155:HV27LDSXX:2:1620:30147:29246 chr1 46241708 N chr1 46242241 N DEL 5
A00297:158:HT275DSXX:2:1672:26512:13432 chr1 46241708 N chr1 46242192 N DEL 2
A00297:158:HT275DSXX:4:2507:22941:23625 chr1 46241408 N chr1 46241635 N DEL 5
A00297:158:HT275DSXX:3:1623:29803:31407 chr1 46241347 N chr1 46241747 N DUP 11
A00404:156:HV37TDSXX:2:2415:29595:13072 chr1 46241347 N chr1 46241747 N DUP 6
A00404:155:HV27LDSXX:4:1347:31675:19680 chr1 46241583 N chr1 46241710 N DEL 7
A00297:158:HT275DSXX:4:1539:29116:18474 chr1 46241753 N chr1 46242284 N DUP 5
A00297:158:HT275DSXX:2:2229:20220:8171 chr1 46241753 N chr1 46242284 N DUP 5
A00404:155:HV27LDSXX:2:2202:12906:3458 chr1 46241753 N chr1 46242284 N DUP 5
A00297:158:HT275DSXX:1:2260:7853:9173 chr1 46241755 N chr1 46242060 N DUP 3
A00404:156:HV37TDSXX:4:1676:32407:9424 chr1 46241756 N chr1 46242238 N DUP 5
A00297:158:HT275DSXX:4:2608:15266:11115 chr1 46241368 N chr1 46241771 N DEL 5
A00404:156:HV37TDSXX:2:1540:27190:17362 chr1 46241383 N chr1 46241786 N DEL 9
A00404:155:HV27LDSXX:3:1539:28474:20964 chr1 46241892 N chr1 46242072 N DEL 10
A00297:158:HT275DSXX:1:2677:1669:10770 chr1 46241397 N chr1 46241800 N DEL 5
A00297:158:HT275DSXX:2:1375:31964:19523 chr1 46241851 N chr1 46241978 N DUP 5
A00404:155:HV27LDSXX:1:2129:21649:33567 chr1 46241795 N chr1 46242583 N DUP 5
A00297:158:HT275DSXX:3:1158:27706:29403 chr1 46241710 N chr1 46241886 N DUP 4
A00297:158:HT275DSXX:4:2652:32895:30311 chr1 46241634 N chr1 46241811 N DEL 5
A00404:155:HV27LDSXX:2:1219:13819:32722 chr1 46241804 N chr1 46242337 N DUP 3
A00404:156:HV37TDSXX:2:2204:9254:26381 chr1 46241637 N chr1 46241814 N DEL 5
A00297:158:HT275DSXX:3:2217:3260:36198 chr1 46241647 N chr1 46241824 N DEL 2
A00297:158:HT275DSXX:2:1672:26512:13432 chr1 46241572 N chr1 46241875 N DEL 7
A00404:155:HV27LDSXX:3:1502:2383:2644 chr1 46241574 N chr1 46241875 N DEL 11
A00404:155:HV27LDSXX:2:1601:18611:13714 chr1 46241909 N chr1 46242089 N DEL 2
A00404:155:HV27LDSXX:4:1334:19307:23813 chr1 46241575 N chr1 46241875 N DEL 13
A00297:158:HT275DSXX:4:1312:11351:30295 chr1 46241909 N chr1 46242089 N DEL 3
A00404:155:HV27LDSXX:4:1461:24659:36276 chr1 46241889 N chr1 46242294 N DUP 1
A00297:158:HT275DSXX:3:2413:7066:27946 chr1 46242003 N chr1 46242182 N DEL 12
A00404:155:HV27LDSXX:2:1250:22607:27806 chr1 46242013 N chr1 46242066 N DEL 5
A00297:158:HT275DSXX:2:1218:14507:33974 chr1 46241485 N chr1 46242013 N DUP 5
A00404:155:HV27LDSXX:1:2616:8431:11710 chr1 46241694 N chr1 46241921 N DEL 5
A00404:155:HV27LDSXX:4:1428:29957:1579 chr1 46241887 N chr1 46242016 N DEL 5
A00297:158:HT275DSXX:2:2229:20220:8171 chr1 46241899 N chr1 46241978 N DEL 3
A00297:158:HT275DSXX:4:2652:32895:30311 chr1 46241746 N chr1 46242052 N DEL 6
A00404:155:HV27LDSXX:3:1577:19397:35556 chr1 46241598 N chr1 46242117 N DUP 1
A00297:158:HT275DSXX:2:1278:3739:34084 chr1 46242149 N chr1 46242248 N DEL 1
A00297:158:HT275DSXX:1:1447:15564:12821 chr1 46241609 N chr1 46242041 N DEL 5
A00404:155:HV27LDSXX:4:1622:29559:16454 chr1 46241609 N chr1 46242041 N DEL 5
A00404:155:HV27LDSXX:3:1565:15347:24690 chr1 46241697 N chr1 46242052 N DEL 6
A00404:155:HV27LDSXX:3:2468:23005:5165 chr1 46241615 N chr1 46242047 N DEL 5
A00404:156:HV37TDSXX:2:2209:18231:14779 chr1 46241910 N chr1 46242088 N DUP 2
A00297:158:HT275DSXX:1:1447:15564:12821 chr1 46241910 N chr1 46242088 N DUP 5
A00404:155:HV27LDSXX:4:1517:14271:14465 chr1 46241385 N chr1 46242095 N DEL 5
A00297:158:HT275DSXX:2:2664:31901:20228 chr1 46242098 N chr1 46242326 N DEL 4
A00404:155:HV27LDSXX:2:1565:15013:32440 chr1 46241623 N chr1 46242107 N DEL 1
A00297:158:HT275DSXX:2:2333:28348:7623 chr1 46241644 N chr1 46242128 N DEL 5
A00404:156:HV37TDSXX:1:2277:28899:8265 chr1 46241572 N chr1 46242182 N DEL 7
A00404:156:HV37TDSXX:2:1357:26847:19805 chr1 46242182 N chr1 46242281 N DUP 10
A00404:156:HV37TDSXX:4:2337:29722:33458 chr1 46241875 N chr1 46242281 N DUP 12
A00404:155:HV27LDSXX:1:1261:5421:17550 chr1 46241875 N chr1 46242233 N DUP 14
A00404:156:HV37TDSXX:4:2275:14543:9204 chr1 46241875 N chr1 46242282 N DUP 14
A00297:158:HT275DSXX:3:2273:13657:36104 chr1 46241875 N chr1 46242280 N DUP 5
A00404:156:HV37TDSXX:3:2677:30897:35681 chr1 46241389 N chr1 46242326 N DEL 5
A00297:158:HT275DSXX:2:1309:26051:11788 chr1 46241443 N chr1 46242380 N DEL 10
A00404:155:HV27LDSXX:4:1517:14271:14465 chr1 46241402 N chr1 46242339 N DEL 5
A00404:156:HV37TDSXX:2:1215:26811:22467 chr1 46241403 N chr1 46242340 N DEL 1
A00404:156:HV37TDSXX:4:1277:15953:27430 chr1 46242041 N chr1 46242448 N DEL 5
A00297:158:HT275DSXX:3:2237:19732:24392 chr1 46241887 N chr1 46242422 N DEL 5
A00404:155:HV27LDSXX:2:1307:11333:5368 chr1 46241746 N chr1 46242457 N DEL 5
A00404:155:HV27LDSXX:2:2661:1787:4742 chr1 46242052 N chr1 46242410 N DEL 5
A00297:158:HT275DSXX:2:1522:23674:10488 chr1 46242325 N chr1 46242504 N DEL 14
A00297:158:HT275DSXX:3:2328:31485:3129 chr1 46241557 N chr1 46242495 N DEL 1
A00404:155:HV27LDSXX:1:2223:24894:9189 chr1 46241553 N chr1 46242491 N DEL 5
A00404:156:HV37TDSXX:1:2277:28899:8265 chr1 46241407 N chr1 46242522 N DEL 5
A00404:155:HV27LDSXX:2:1657:12861:34851 chr1 46241421 N chr1 46242536 N DEL 1
A00404:155:HV27LDSXX:2:2173:12129:29919 chr1 46241421 N chr1 46242536 N DEL 1
A00404:155:HV27LDSXX:2:1574:26069:6965 chr5 102050836 N chr5 102050943 N DUP 14
A00404:156:HV37TDSXX:1:1607:14235:27211 chr5 102050937 N chr5 102051000 N DEL 12
A00297:158:HT275DSXX:4:1313:19660:19351 chr5 102050937 N chr5 102051000 N DEL 14
A00404:155:HV27LDSXX:4:2436:5855:9940 chr5 102050857 N chr5 102051000 N DEL 7
A00404:155:HV27LDSXX:4:2436:7536:23844 chr5 102050884 N chr5 102051029 N DEL 8
A00297:158:HT275DSXX:3:1360:30743:33536 chr5 102050857 N chr5 102051000 N DEL 7
A00297:158:HT275DSXX:1:1658:20808:11851 chr5 102051092 N chr5 102051227 N DEL 5
A00404:156:HV37TDSXX:2:1666:23737:14168 chr5 102050863 N chr5 102051006 N DEL 7
A00404:155:HV27LDSXX:3:1313:31729:8563 chr5 102050967 N chr5 102051060 N DEL 12
A00404:155:HV27LDSXX:3:1313:32371:8171 chr5 102050967 N chr5 102051060 N DEL 12
A00404:156:HV37TDSXX:4:2427:1814:23766 chr5 102050858 N chr5 102051061 N DEL 7
A00404:156:HV37TDSXX:1:1677:10267:2394 chr5 102050880 N chr5 102051083 N DEL 1
A00297:158:HT275DSXX:1:2556:27615:22263 chr5 102051125 N chr5 102051258 N DEL 10
A00404:155:HV27LDSXX:4:2435:12310:5963 chr5 102051125 N chr5 102051258 N DEL 14
A00297:158:HT275DSXX:2:2607:1976:32534 chr5 102051125 N chr5 102051258 N DEL 14
A00404:155:HV27LDSXX:4:2435:11577:5353 chr5 102051125 N chr5 102051258 N DEL 14
A00404:155:HV27LDSXX:4:1424:25120:22921 chr5 102050834 N chr5 102051259 N DEL 9
A00404:155:HV27LDSXX:4:1424:25328:23312 chr5 102050834 N chr5 102051259 N DEL 9
A00297:158:HT275DSXX:2:2556:29071:27226 chr5 102051105 N chr5 102051430 N DUP 5
A00297:158:HT275DSXX:4:2560:16920:27696 chr5 102051105 N chr5 102051430 N DUP 5
A00404:156:HV37TDSXX:2:1666:23737:14168 chr5 102051105 N chr5 102051430 N DUP 5
A00404:155:HV27LDSXX:1:2124:27679:21715 chr5 102051089 N chr5 102051352 N DEL 5
A00404:155:HV27LDSXX:1:2145:9570:34914 chr5 102050856 N chr5 102051347 N DEL 6
A00404:155:HV27LDSXX:2:1635:1958:33160 chr5 102051089 N chr5 102051352 N DEL 5
A00297:158:HT275DSXX:1:1658:20808:11851 chr5 102051119 N chr5 102051412 N DEL 5
A00404:156:HV37TDSXX:2:2267:24089:22326 chr5 102050830 N chr5 102051417 N DEL 2
A00404:156:HV37TDSXX:2:2267:24424:21089 chr5 102050830 N chr5 102051417 N DEL 2
A00297:158:HT275DSXX:1:2630:7030:11412 chr5 102051245 N chr5 102051472 N DEL 5
A00297:158:HT275DSXX:2:2607:1976:32534 chr5 102051245 N chr5 102051472 N DEL 5
A00404:156:HV37TDSXX:2:1271:31684:3568 chr5 102051245 N chr5 102051472 N DEL 5
A00297:158:HT275DSXX:3:2662:26042:19225 chr5 102051245 N chr5 102051472 N DEL 5
A00297:158:HT275DSXX:1:2556:27615:22263 chr5 102050856 N chr5 102051481 N DEL 5
A00404:156:HV37TDSXX:4:1353:10140:9314 chr1 88579064 N chr1 88579337 N DEL 13
A00297:158:HT275DSXX:1:2102:14253:12962 chr1 88579056 N chr1 88579329 N DEL 8
A00297:158:HT275DSXX:3:2673:7690:14184 chr2 20834753 N chr2 20834820 N DEL 8
A00404:155:HV27LDSXX:1:2126:7319:25379 chrX 66559931 N chrX 66560008 N DEL 5
A00404:155:HV27LDSXX:1:2522:25690:24283 chr7 158327405 N chr7 158327466 N DUP 4
A00297:158:HT275DSXX:4:2623:15266:17002 chr7 158327312 N chr7 158327524 N DUP 8
A00404:156:HV37TDSXX:3:1432:19732:16908 chr7 158327524 N chr7 158327586 N DEL 13
A00404:155:HV27LDSXX:3:1165:18258:34648 chr7 158327451 N chr7 158327514 N DEL 5
A00404:155:HV27LDSXX:2:2460:30563:27962 chr7 158327451 N chr7 158327514 N DEL 5
A00404:156:HV37TDSXX:4:1151:7609:9909 chr7 158327303 N chr7 158327622 N DUP 9
A00404:156:HV37TDSXX:1:1260:31566:19805 chr7 158327303 N chr7 158327622 N DUP 9
A00404:156:HV37TDSXX:1:1260:32009:18787 chr7 158327303 N chr7 158327622 N DUP 9
A00404:155:HV27LDSXX:2:1278:21432:7983 chr7 158327303 N chr7 158327622 N DUP 9
A00404:156:HV37TDSXX:4:2366:24343:32847 chr7 158327577 N chr7 158327630 N DEL 9
A00297:158:HT275DSXX:1:2142:21884:7639 chr7 158327577 N chr7 158327630 N DEL 9
A00404:155:HV27LDSXX:4:2206:20853:4820 chr7 158327577 N chr7 158327630 N DEL 9
A00404:156:HV37TDSXX:3:2453:28492:7936 chr7 158327577 N chr7 158327630 N DEL 9
A00297:158:HT275DSXX:2:1304:29649:10410 chrY 16324624 N chrY 16324691 N DEL 10
A00297:158:HT275DSXX:1:2625:30138:28635 chr7 152740304 N chr7 152740385 N DEL 2
A00404:155:HV27LDSXX:2:2576:6732:35164 chr7 152740365 N chr7 152740424 N DUP 5
A00297:158:HT275DSXX:4:2403:22878:3004 chr7 152740340 N chr7 152740408 N DUP 12
A00297:158:HT275DSXX:1:2519:10565:32753 chr7 152740314 N chr7 152740404 N DEL 9
A00297:158:HT275DSXX:1:1356:11695:10629 chr2 231264393 N chr2 231264713 N DEL 24
A00404:155:HV27LDSXX:2:1167:28809:17315 chr2 231264588 N chr2 231264907 N DEL 5
A00297:158:HT275DSXX:1:2408:3477:3881 chr2 231264413 N chr2 231264733 N DEL 42
A00404:155:HV27LDSXX:2:1167:28809:17315 chr2 231264535 N chr2 231264854 N DEL 20
A00404:156:HV37TDSXX:1:1644:11008:1892 chr1 240868205 N chr1 240868277 N DEL 5
A00404:155:HV27LDSXX:1:2678:31819:34741 chr1 240868206 N chr1 240868278 N DEL 4
A00297:158:HT275DSXX:3:2557:20012:1861 chr19 50538873 N chr19 50539034 N DUP 5
A00404:156:HV37TDSXX:3:1174:13539:3521 chr7 29749000 N chr7 29749070 N DUP 4
A00404:155:HV27LDSXX:1:2502:2600:6872 chr5 147765119 N chr5 147765196 N DUP 16
A00404:155:HV27LDSXX:4:1334:1814:4225 chr5 147765119 N chr5 147765196 N DUP 16
A00297:158:HT275DSXX:4:2230:4996:27054 chr1 2788509 N chr1 2788590 N DUP 5
A00404:156:HV37TDSXX:2:2429:19443:35947 chr17 30679553 N chr17 30679700 N DEL 23
A00404:155:HV27LDSXX:4:2262:21052:6386 chr17 30679563 N chr17 30679881 N DEL 3
A00404:156:HV37TDSXX:1:2629:31521:33285 chr19 1963511 N chr19 1963808 N DEL 10
A00404:156:HV37TDSXX:2:2662:21811:20979 chr19 20823109 N chr19 20823201 N DEL 5
A00404:156:HV37TDSXX:4:1523:30698:11569 chr19 20823109 N chr19 20823201 N DEL 10
A00404:155:HV27LDSXX:3:2424:12174:12461 chr19 20823096 N chr19 20823281 N DEL 6
A00404:155:HV27LDSXX:2:2260:13150:21198 chr19 20823096 N chr19 20823281 N DEL 9
A00404:155:HV27LDSXX:4:1469:6352:9204 chr19 20823096 N chr19 20823281 N DEL 10
A00404:156:HV37TDSXX:2:2503:23466:22185 chr19 20823096 N chr19 20823281 N DEL 13
A00404:156:HV37TDSXX:2:2577:6361:21778 chr19 20823096 N chr19 20823281 N DEL 20
A00404:156:HV37TDSXX:2:2577:7708:21668 chr19 20823096 N chr19 20823281 N DEL 20
A00404:156:HV37TDSXX:3:1447:9661:22420 chr19 20823096 N chr19 20823281 N DEL 22
A00404:156:HV37TDSXX:1:1104:3685:36464 chr19 20823096 N chr19 20823281 N DEL 31
A00404:156:HV37TDSXX:1:2622:10990:4961 chr19 20823097 N chr19 20823282 N DEL 14
A00297:158:HT275DSXX:3:1219:27245:27665 chr19 20823098 N chr19 20823283 N DEL 13
A00297:158:HT275DSXX:3:1309:10321:10191 chr19 20823104 N chr19 20823289 N DEL 7
A00297:158:HT275DSXX:3:1309:10917:10222 chr19 20823104 N chr19 20823289 N DEL 7
A00297:158:HT275DSXX:4:2201:8440:33051 chr19 20823104 N chr19 20823289 N DEL 7
A00404:156:HV37TDSXX:3:1577:19497:12994 chr19 20823100 N chr19 20823285 N DEL 11
A00404:156:HV37TDSXX:4:1248:4915:31892 chr19 20823097 N chr19 20823282 N DEL 14
A00404:156:HV37TDSXX:3:1220:32515:31031 chr19 20823096 N chr19 20823281 N DEL 16
A00404:155:HV27LDSXX:4:1177:13250:12101 chr19 20823096 N chr19 20823281 N DEL 18
A00297:158:HT275DSXX:1:2260:7374:28855 chr19 20823217 N chr19 20823280 N DEL 5
A00297:158:HT275DSXX:3:2668:1524:11459 chr19 20823223 N chr19 20823286 N DEL 5
A00297:158:HT275DSXX:4:1307:24334:29825 chr19 20823222 N chr19 20823285 N DEL 5
A00404:155:HV27LDSXX:4:1659:18765:10128 chr19 20823100 N chr19 20823285 N DEL 11
A00404:156:HV37TDSXX:1:1409:3902:16517 chr19 20823096 N chr19 20823281 N DEL 22
A00404:155:HV27LDSXX:1:1104:10881:25254 chr19 20823096 N chr19 20823281 N DEL 15
A00297:158:HT275DSXX:1:1663:18412:20322 chr19 20823096 N chr19 20823281 N DEL 15
A00404:155:HV27LDSXX:2:1509:8458:12038 chr19 20823385 N chr19 20823449 N DEL 5
A00404:155:HV27LDSXX:4:1162:14850:7607 chr19 20823385 N chr19 20823449 N DEL 5
A00404:155:HV27LDSXX:4:1162:16251:6402 chr19 20823140 N chr19 20823507 N DUP 10
A00404:155:HV27LDSXX:4:1120:2636:16454 chr19 20823385 N chr19 20823449 N DEL 5
A00297:158:HT275DSXX:3:1309:10321:10191 chr19 20823232 N chr19 20823508 N DUP 5
A00297:158:HT275DSXX:3:1309:10917:10222 chr19 20823232 N chr19 20823508 N DUP 5
A00297:158:HT275DSXX:4:2201:8440:33051 chr19 20823232 N chr19 20823508 N DUP 5
A00404:156:HV37TDSXX:3:2520:17318:29105 chr19 20823232 N chr19 20823508 N DUP 5
A00404:156:HV37TDSXX:4:2108:26657:16250 chr19 20823294 N chr19 20823508 N DUP 5
A00404:156:HV37TDSXX:3:1626:13566:12305 chr19 20823257 N chr19 20823535 N DEL 5
A00404:156:HV37TDSXX:1:2260:16288:34366 chr19 20823258 N chr19 20823536 N DEL 5
A00297:158:HT275DSXX:4:2513:27362:10269 chr19 20823198 N chr19 20823538 N DEL 4
A00297:158:HT275DSXX:4:2513:30445:16642 chr19 20823198 N chr19 20823538 N DEL 4
A00404:155:HV27LDSXX:4:2256:29134:2534 chr5 101088069 N chr5 101088134 N DEL 5
A00404:156:HV37TDSXX:1:2133:13883:18302 chr5 101088069 N chr5 101088134 N DEL 7
A00404:155:HV27LDSXX:2:1119:30255:30499 chr5 101088069 N chr5 101088134 N DEL 18
A00404:156:HV37TDSXX:2:2375:16450:22498 chr5 101088069 N chr5 101088134 N DEL 21
A00404:155:HV27LDSXX:2:2337:21513:16391 chr5 101088069 N chr5 101088134 N DEL 26
A00404:155:HV27LDSXX:2:2337:21522:16376 chr5 101088069 N chr5 101088134 N DEL 24
A00404:156:HV37TDSXX:4:1473:20374:30483 chr5 101088073 N chr5 101088238 N DUP 29
A00297:158:HT275DSXX:3:1509:28610:6668 chr5 101088106 N chr5 101088239 N DUP 6
A00404:156:HV37TDSXX:1:1617:12111:31829 chr5 101088106 N chr5 101088239 N DUP 6
A00404:156:HV37TDSXX:1:2569:12762:9784 chr5 101088073 N chr5 101088238 N DUP 27
A00404:155:HV27LDSXX:3:1213:28971:35227 chr5 101088105 N chr5 101088202 N DUP 14
A00404:155:HV27LDSXX:3:1120:6515:4664 chr5 101088137 N chr5 101088238 N DUP 20
A00404:156:HV37TDSXX:2:1672:10257:12743 chr5 101088137 N chr5 101088238 N DUP 21
A00297:158:HT275DSXX:1:1622:11333:9690 chr5 101088169 N chr5 101088238 N DUP 20
A00297:158:HT275DSXX:4:2159:19262:34569 chr5 101088169 N chr5 101088238 N DUP 21
A00404:156:HV37TDSXX:4:1578:25735:25175 chr5 101088137 N chr5 101088238 N DUP 21
A00297:158:HT275DSXX:4:2667:7808:5556 chr5 101088137 N chr5 101088238 N DUP 21
A00404:155:HV27LDSXX:3:2556:27118:11005 chr5 101088137 N chr5 101088238 N DUP 21
A00297:158:HT275DSXX:1:2340:19488:36119 chr5 101088169 N chr5 101088238 N DUP 20
A00404:155:HV27LDSXX:3:1566:22905:3082 chr5 101088137 N chr5 101088238 N DUP 21
A00404:155:HV27LDSXX:3:2566:21477:12132 chr5 101088137 N chr5 101088238 N DUP 21
A00404:155:HV27LDSXX:4:1375:21206:12164 chr5 101088105 N chr5 101088202 N DUP 14
A00404:155:HV27LDSXX:4:2375:20464:20494 chr5 101088105 N chr5 101088202 N DUP 14
A00404:155:HV27LDSXX:4:2375:20672:20635 chr5 101088105 N chr5 101088202 N DUP 14
A00404:156:HV37TDSXX:1:2615:9435:15828 chr5 101088105 N chr5 101088202 N DUP 14
A00297:158:HT275DSXX:3:2139:23854:22795 chr5 101088137 N chr5 101088238 N DUP 21
A00404:155:HV27LDSXX:4:2237:10004:21198 chr5 101088137 N chr5 101088238 N DUP 21
A00404:155:HV27LDSXX:4:2254:27208:28166 chr5 101088169 N chr5 101088238 N DUP 20
A00297:158:HT275DSXX:4:1568:11605:35837 chr5 101088137 N chr5 101088238 N DUP 20
A00404:156:HV37TDSXX:2:1439:28483:3537 chr5 101088169 N chr5 101088238 N DUP 20
A00297:158:HT275DSXX:2:1303:3441:15562 chr5 101088137 N chr5 101088238 N DUP 19
A00297:158:HT275DSXX:3:2571:28167:30201 chr5 101088137 N chr5 101088238 N DUP 19
A00297:158:HT275DSXX:1:1632:9001:13197 chr5 101088105 N chr5 101088202 N DUP 13
A00404:155:HV27LDSXX:4:1135:13612:36276 chr5 101088105 N chr5 101088202 N DUP 13
A00297:158:HT275DSXX:1:1113:27697:32706 chr5 101088137 N chr5 101088238 N DUP 16
A00297:158:HT275DSXX:2:1436:18602:22467 chr5 101088137 N chr5 101088238 N DUP 16
A00297:158:HT275DSXX:3:1174:12491:8719 chr5 101088137 N chr5 101088238 N DUP 16
A00297:158:HT275DSXX:3:2170:8449:26678 chr5 101088137 N chr5 101088238 N DUP 15
A00297:158:HT275DSXX:1:2660:4535:3208 chr5 101088169 N chr5 101088238 N DUP 15
A00404:155:HV27LDSXX:3:2556:27118:11005 chr5 101088137 N chr5 101088238 N DUP 18
A00404:155:HV27LDSXX:3:1120:6515:4664 chr5 101088169 N chr5 101088238 N DUP 20
A00404:156:HV37TDSXX:4:1521:27416:24612 chr5 101088137 N chr5 101088238 N DUP 18
A00404:155:HV27LDSXX:1:1173:29125:20149 chr5 101088169 N chr5 101088238 N DUP 16
A00297:158:HT275DSXX:1:2660:4535:3208 chr5 101088098 N chr5 101088231 N DUP 2
A00404:155:HV27LDSXX:2:2235:25870:36526 chr5 101088098 N chr5 101088231 N DUP 2
A00404:155:HV27LDSXX:3:1675:31566:20369 chr5 101088098 N chr5 101088231 N DUP 2
A00297:158:HT275DSXX:1:1654:27181:2534 chr5 101088069 N chr5 101088134 N DEL 26
A00404:155:HV27LDSXX:3:2148:21793:27367 chr5 101088069 N chr5 101088134 N DEL 24
A00297:158:HT275DSXX:4:2415:24786:34147 chr5 101088069 N chr5 101088134 N DEL 24
A00404:156:HV37TDSXX:4:2646:20473:12555 chr5 101088069 N chr5 101088134 N DEL 26
A00404:155:HV27LDSXX:1:1133:22950:5134 chr5 101088069 N chr5 101088134 N DEL 25
A00404:156:HV37TDSXX:4:1411:18231:26929 chr5 101088079 N chr5 101088144 N DEL 5
A00404:155:HV27LDSXX:2:1501:18557:13182 chr8 2080935 N chr8 2080987 N DEL 1
A00404:156:HV37TDSXX:4:1602:6153:26929 chr8 2081098 N chr8 2081306 N DEL 1
A00404:155:HV27LDSXX:1:2207:17011:25003 chr8 2081098 N chr8 2081409 N DEL 5
A00297:158:HT275DSXX:1:2456:26313:24549 chr8 2081016 N chr8 2081430 N DEL 7
A00404:155:HV27LDSXX:2:1469:27199:11960 chr8 2081264 N chr8 2081315 N DUP 12
A00404:155:HV27LDSXX:2:1123:22860:20509 chr8 2081268 N chr8 2081474 N DUP 5
A00404:155:HV27LDSXX:2:2539:4797:21543 chr8 2081272 N chr8 2081478 N DUP 5
A00404:155:HV27LDSXX:2:1628:29460:28401 chr8 2081371 N chr8 2081474 N DUP 5
A00404:156:HV37TDSXX:1:1510:30101:15640 chr8 2081371 N chr8 2081474 N DUP 5
A00404:155:HV27LDSXX:4:2349:31394:4946 chr8 2081371 N chr8 2081474 N DUP 5
A00297:158:HT275DSXX:3:2358:23258:1971 chr8 2081199 N chr8 2081510 N DEL 5
A00297:158:HT275DSXX:1:2456:26313:24549 chr8 2081199 N chr8 2081510 N DEL 5
A00404:156:HV37TDSXX:3:2213:5565:14669 chr8 2080992 N chr8 2081510 N DEL 5
A00404:156:HV37TDSXX:4:1226:16034:8813 chr8 2080992 N chr8 2081510 N DEL 5
A00404:155:HV27LDSXX:3:2401:32741:35587 chr8 2080992 N chr8 2081510 N DEL 5
A00404:156:HV37TDSXX:2:1116:2636:16172 chr8 2080998 N chr8 2081516 N DEL 5
A00297:158:HT275DSXX:3:2229:1470:21167 chr8 2080953 N chr8 2081522 N DEL 3
A00297:158:HT275DSXX:3:2229:1723:21104 chr8 2080953 N chr8 2081522 N DEL 3
A00404:156:HV37TDSXX:2:2320:23366:17973 chr8 2080953 N chr8 2081522 N DEL 3
A00404:156:HV37TDSXX:2:2320:23981:17848 chr8 2080953 N chr8 2081522 N DEL 3
A00404:155:HV27LDSXX:4:2144:25880:9706 chr13 95690766 N chr13 95691071 N DEL 5
A00297:158:HT275DSXX:3:1364:15935:11553 chr13 95690825 N chr13 95691078 N DUP 5
A00297:158:HT275DSXX:2:1205:27751:19116 chr13 95690858 N chr13 95690986 N DEL 7
A00404:156:HV37TDSXX:3:1218:24975:35102 chr13 95690851 N chr13 95690979 N DEL 10
A00404:155:HV27LDSXX:2:2340:17824:18646 chr13 95690768 N chr13 95691071 N DUP 1
A00404:156:HV37TDSXX:2:1436:8341:5729 chr13 95690770 N chr13 95691122 N DUP 3
A00404:155:HV27LDSXX:3:2433:31665:34319 chr13 95690768 N chr13 95691071 N DUP 9
A00404:155:HV27LDSXX:2:2153:30210:20619 chr13 95690819 N chr13 95691124 N DEL 3
A00404:156:HV37TDSXX:4:2627:24406:24596 chr13 95690770 N chr13 95691074 N DEL 2
A00297:158:HT275DSXX:2:1433:8974:23735 chr5 123750303 N chr5 123750502 N DUP 5
A00297:158:HT275DSXX:1:1174:6976:32174 chr5 123750303 N chr5 123750502 N DUP 8
A00297:158:HT275DSXX:2:2654:8043:25723 chr5 123750303 N chr5 123750502 N DUP 3
A00404:155:HV27LDSXX:4:2530:28772:21355 chr11 131266346 N chr11 131266407 N DUP 5
A00404:155:HV27LDSXX:2:1354:14886:24486 chr11 131266346 N chr11 131266407 N DUP 5
A00404:156:HV37TDSXX:3:2519:21477:5776 chr11 131266346 N chr11 131266407 N DUP 5
A00404:155:HV27LDSXX:2:1468:13765:27023 chr11 131266346 N chr11 131266407 N DUP 5
A00297:158:HT275DSXX:3:1542:6298:1752 chr11 131266346 N chr11 131266407 N DUP 5
A00404:155:HV27LDSXX:3:2155:32579:19304 chr8 69626268 N chr8 69626386 N DEL 5
A00404:155:HV27LDSXX:2:2312:9200:31892 chr8 69626268 N chr8 69626386 N DEL 15
A00404:156:HV37TDSXX:2:1521:10493:31093 chr8 69626268 N chr8 69626386 N DEL 15
A00297:158:HT275DSXX:4:1237:14642:4241 chr8 69626268 N chr8 69626386 N DEL 33
A00297:158:HT275DSXX:2:1139:26802:27743 chr8 69626268 N chr8 69626386 N DEL 34
A00297:158:HT275DSXX:2:1465:29875:4946 chr8 69626268 N chr8 69626386 N DEL 39
A00404:156:HV37TDSXX:3:2343:27489:7733 chr8 69626140 N chr8 69626299 N DEL 7
A00404:156:HV37TDSXX:4:1641:14262:23688 chr8 69626277 N chr8 69626395 N DEL 6
A00404:156:HV37TDSXX:1:1437:6614:27821 chr8 69626278 N chr8 69626396 N DEL 5
A00404:156:HV37TDSXX:4:1327:29179:24659 chr8 69626278 N chr8 69626396 N DEL 5
A00404:156:HV37TDSXX:4:2327:30653:19601 chr8 69626278 N chr8 69626396 N DEL 5
A00404:155:HV27LDSXX:4:2374:27905:19163 chr4 53237672 N chr4 53237798 N DUP 10
A00404:156:HV37TDSXX:4:2269:24813:35352 chr4 53237703 N chr4 53237780 N DUP 7
A00297:158:HT275DSXX:2:2158:4924:30405 chr4 53237692 N chr4 53237818 N DUP 5
A00404:156:HV37TDSXX:1:1209:29731:18098 chr4 53237774 N chr4 53238184 N DEL 10
A00297:158:HT275DSXX:3:1325:1172:10629 chr4 53237690 N chr4 53237816 N DUP 10
A00404:156:HV37TDSXX:1:1317:4318:36213 chr4 53237936 N chr4 53238013 N DUP 10
A00404:156:HV37TDSXX:4:2269:24813:35352 chr4 53237819 N chr4 53238227 N DUP 5
A00404:155:HV27LDSXX:2:1552:3739:13604 chr4 53237627 N chr4 53237801 N DEL 1
A00297:158:HT275DSXX:4:1605:29215:22592 chr4 53237744 N chr4 53237870 N DUP 5
A00404:155:HV27LDSXX:2:1635:15185:34554 chr4 53237743 N chr4 53237869 N DUP 5
A00404:155:HV27LDSXX:4:1477:1705:36573 chr4 53237646 N chr4 53238130 N DUP 1
A00297:158:HT275DSXX:2:1663:16550:5040 chr4 53237816 N chr4 53238079 N DEL 14
A00404:155:HV27LDSXX:4:2533:21007:9251 chr4 53237706 N chr4 53238047 N DEL 5
A00297:158:HT275DSXX:2:1535:18249:34569 chr4 53237816 N chr4 53238079 N DEL 8
A00297:158:HT275DSXX:2:2410:5430:33317 chr4 53237774 N chr4 53238086 N DEL 4
A00404:156:HV37TDSXX:3:1605:31412:29215 chr4 53238019 N chr4 53238214 N DUP 12
A00404:155:HV27LDSXX:3:1535:11460:9846 chr4 53237738 N chr4 53238273 N DUP 5
A00404:155:HV27LDSXX:4:2574:30535:4210 chr4 53237738 N chr4 53238273 N DUP 8
A00404:155:HV27LDSXX:3:2257:24279:3239 chr4 53238152 N chr4 53238327 N DUP 5
A00297:158:HT275DSXX:1:2557:17354:28635 chr10 31969116 N chr10 31969212 N DEL 6
A00404:155:HV27LDSXX:2:2438:24433:22576 chr10 31969133 N chr10 31969202 N DUP 5
A00297:158:HT275DSXX:3:1236:24849:19633 chr10 31969125 N chr10 31969276 N DUP 5
A00297:158:HT275DSXX:1:2171:20500:10848 chr10 31969183 N chr10 31969247 N DEL 11
A00404:156:HV37TDSXX:2:1224:3938:31767 chr10 31969145 N chr10 31969247 N DEL 11
A00297:158:HT275DSXX:4:1149:3929:15029 chr10 31969132 N chr10 31969253 N DEL 9
A00404:155:HV27LDSXX:4:1646:2202:21903 chr10 31969132 N chr10 31969253 N DEL 9
A00404:155:HV27LDSXX:1:1172:28574:10614 chr10 31969162 N chr10 31969277 N DEL 5
A00404:155:HV27LDSXX:2:2648:17770:17926 chr5 4843864 N chr5 4843976 N DUP 7
A00404:156:HV37TDSXX:1:2563:7473:21230 chr5 4843864 N chr5 4843976 N DUP 10
A00404:155:HV27LDSXX:1:2220:19795:13072 chr5 4843984 N chr5 4844039 N DEL 8
A00404:156:HV37TDSXX:1:1257:28700:22764 chr5 4843984 N chr5 4844039 N DEL 16
A00404:156:HV37TDSXX:2:2514:31367:29387 chr5 4843984 N chr5 4844039 N DEL 28
A00404:155:HV27LDSXX:3:2108:29668:6872 chr5 4843984 N chr5 4844039 N DEL 31
A00404:156:HV37TDSXX:2:1353:19660:13620 chr6 114560614 N chr6 114560695 N DEL 1
A00404:156:HV37TDSXX:4:1308:30843:22216 chr6 114560598 N chr6 114560726 N DUP 1
A00404:156:HV37TDSXX:4:2101:24948:29262 chr7 61056204 N chr7 61056441 N DUP 5
A00404:155:HV27LDSXX:3:2265:23475:24205 chr7 61056168 N chr7 61056267 N DEL 10
A00404:156:HV37TDSXX:1:2521:11586:25880 chr7 61056299 N chr7 61056435 N DUP 3
A00404:155:HV27LDSXX:3:2473:28962:19335 chr7 61056164 N chr7 61056364 N DEL 20
A00404:155:HV27LDSXX:4:1205:22146:16579 chr19 15972421 N chr19 15972504 N DEL 12
A00297:158:HT275DSXX:1:1341:16450:14982 chr17 21843747 N chr17 21843816 N DEL 16
A00404:156:HV37TDSXX:4:2169:6822:34287 chrX 627035 N chrX 627148 N DUP 10
A00297:158:HT275DSXX:1:2107:13675:34569 chrX 627060 N chrX 627138 N DEL 2
A00404:155:HV27LDSXX:3:1370:16360:24565 chr1 210976351 N chr1 210976705 N DEL 5
A00404:156:HV37TDSXX:1:1204:10511:20165 chr1 210976351 N chr1 210976705 N DEL 5
A00297:158:HT275DSXX:4:1502:17861:30389 chr1 210976351 N chr1 210976705 N DEL 5
A00297:158:HT275DSXX:2:2218:19904:10880 chr1 210976351 N chr1 210976705 N DEL 5
A00297:158:HT275DSXX:2:1425:4472:28714 chr1 210976351 N chr1 210976705 N DEL 5
A00297:158:HT275DSXX:2:1425:4481:28729 chr1 210976351 N chr1 210976705 N DEL 5
A00297:158:HT275DSXX:1:1535:15528:20682 chr1 210976351 N chr1 210976705 N DEL 5
A00404:156:HV37TDSXX:2:2259:30210:30044 chr1 210976351 N chr1 210976705 N DEL 5
A00297:158:HT275DSXX:2:2218:19904:10880 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:4:1149:11623:10097 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:4:1565:19461:11209 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:1:2630:28067:31000 chr1 210976351 N chr1 210976705 N DEL 5
A00404:156:HV37TDSXX:4:2645:2781:10128 chr1 210976351 N chr1 210976705 N DEL 5
A00404:156:HV37TDSXX:3:1234:24903:30624 chr1 210976578 N chr1 210976932 N DEL 5
A00404:155:HV27LDSXX:4:1376:28890:21903 chr1 210976680 N chr1 210977032 N DUP 1
A00297:158:HT275DSXX:1:1426:29568:26584 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:1:2275:3414:19523 chr1 210976680 N chr1 210977032 N DUP 5
A00404:155:HV27LDSXX:1:2211:5150:30577 chr1 210976680 N chr1 210977032 N DUP 5
A00404:155:HV27LDSXX:1:2675:9182:7623 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:1:1473:3495:25050 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:3:2527:14217:22169 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:1:1620:24605:28573 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:4:2331:7997:33411 chr1 210976680 N chr1 210977032 N DUP 5
A00404:155:HV27LDSXX:1:2151:11198:24893 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:1:2571:9986:15749 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:1:1632:9263:22388 chr1 210976680 N chr1 210977032 N DUP 5
A00297:158:HT275DSXX:4:1565:6931:17816 chr1 210976680 N chr1 210977032 N DUP 5
A00404:156:HV37TDSXX:1:1609:20455:23422 chr1 210976697 N chr1 210977051 N DEL 5
A00404:155:HV27LDSXX:2:1204:4562:4194 chr1 210976698 N chr1 210977052 N DEL 5
A00404:155:HV27LDSXX:2:1204:8287:1532 chr1 210976698 N chr1 210977052 N DEL 5
A00404:155:HV27LDSXX:1:1237:30129:22138 chr1 210976701 N chr1 210977055 N DEL 5
A00404:156:HV37TDSXX:2:2634:11442:22592 chr1 210976703 N chr1 210977057 N DEL 5
A00404:155:HV27LDSXX:2:1110:12608:26303 chr5 344553 N chr5 344646 N DEL 20
A00404:155:HV27LDSXX:4:1572:9516:32252 chr5 344615 N chr5 344875 N DUP 5
A00404:156:HV37TDSXX:1:1167:31141:15969 chr2 119444274 N chr2 119444431 N DUP 5
A00404:156:HV37TDSXX:4:2236:4101:32863 chr2 119444459 N chr2 119444536 N DUP 31
A00297:158:HT275DSXX:2:2265:32298:30248 chr2 119444459 N chr2 119444536 N DUP 31
A00404:156:HV37TDSXX:4:2205:20934:14262 chr2 119444459 N chr2 119444510 N DUP 16
A00297:158:HT275DSXX:1:1665:2031:4820 chr2 119444459 N chr2 119444510 N DUP 22
A00297:158:HT275DSXX:3:1457:6488:6590 chr2 119444459 N chr2 119444536 N DUP 29
A00404:155:HV27LDSXX:1:2640:8919:21856 chr2 119444459 N chr2 119444536 N DUP 29
A00404:156:HV37TDSXX:3:1467:32868:15358 chr2 119444459 N chr2 119444536 N DUP 29
A00297:158:HT275DSXX:4:2432:32072:31046 chr2 119444459 N chr2 119444536 N DUP 28
A00297:158:HT275DSXX:4:2552:21884:29089 chr2 119444459 N chr2 119444536 N DUP 27
A00297:158:HT275DSXX:1:1371:31485:26428 chr2 119444459 N chr2 119444536 N DUP 29
A00297:158:HT275DSXX:3:2339:24822:27195 chr2 119444440 N chr2 119444563 N DUP 21
A00404:156:HV37TDSXX:1:1167:31141:15969 chr2 119444459 N chr2 119444536 N DUP 30
A00404:156:HV37TDSXX:2:2137:14208:13416 chr2 119444459 N chr2 119444536 N DUP 31
A00297:158:HT275DSXX:1:1171:15501:1532 chr13 36317549 N chr13 36317631 N DUP 5
A00297:158:HT275DSXX:1:1171:15709:1611 chr13 36317549 N chr13 36317631 N DUP 5
A00297:158:HT275DSXX:1:2608:27019:2566 chr13 36317564 N chr13 36317648 N DEL 5
A00404:155:HV27LDSXX:3:1447:23466:27289 chr13 36317565 N chr13 36317649 N DEL 5
A00404:155:HV27LDSXX:2:2536:28456:31422 chr13 36317568 N chr13 36317652 N DEL 5
A00404:155:HV27LDSXX:4:1424:16839:24956 chr11 1159666 N chr11 1159821 N DEL 3
A00297:158:HT275DSXX:2:1328:13512:31782 chr11 1159666 N chr11 1159821 N DEL 4
A00297:158:HT275DSXX:4:2334:6931:6167 chr11 1159691 N chr11 1159836 N DEL 10
A00297:158:HT275DSXX:1:2668:1497:18584 chr11 1159691 N chr11 1159836 N DEL 13
A00297:158:HT275DSXX:2:2264:27805:10504 chr11 1159691 N chr11 1159836 N DEL 16
A00404:155:HV27LDSXX:3:2374:12771:11365 chr11 1159738 N chr11 1159861 N DUP 10
A00297:158:HT275DSXX:3:1546:1280:3458 chr11 1159688 N chr11 1159796 N DEL 30
A00297:158:HT275DSXX:2:1613:7952:16329 chr11 1159752 N chr11 1159865 N DUP 6
A00404:155:HV27LDSXX:2:2347:8693:2895 chr11 1159748 N chr11 1159861 N DUP 5
A00297:158:HT275DSXX:2:1226:16297:28244 chr3 17119887 N chr3 17120158 N DEL 8
A00404:155:HV27LDSXX:1:1407:10908:13056 chr3 17119979 N chr3 17120143 N DEL 5
A00297:158:HT275DSXX:1:1436:17146:36104 chr22 36728233 N chr22 36728335 N DUP 1
A00297:158:HT275DSXX:1:1618:7401:34914 chr22 36728233 N chr22 36728335 N DUP 6
A00404:156:HV37TDSXX:2:1278:30291:35070 chr22 36728233 N chr22 36728335 N DUP 2
A00404:155:HV27LDSXX:2:1456:6325:24972 chr22 36728264 N chr22 36728366 N DEL 4
A00404:156:HV37TDSXX:2:2271:11107:31219 chr22 36728264 N chr22 36728366 N DEL 4
A00404:156:HV37TDSXX:2:1673:2022:31360 chr22 36728261 N chr22 36728363 N DEL 9
A00404:155:HV27LDSXX:2:1237:29351:30279 chr22 36728267 N chr22 36728369 N DEL 9
A00404:155:HV27LDSXX:2:1206:27263:20149 chr5 1871123 N chr5 1871324 N DUP 9
A00297:158:HT275DSXX:3:1152:10402:7012 chr5 1871255 N chr5 1871320 N DUP 5
A00297:158:HT275DSXX:1:1420:8784:22936 chr5 1871222 N chr5 1871289 N DEL 35
A00404:156:HV37TDSXX:3:1263:23493:13213 chr2 104519712 N chr2 104519838 N DEL 5
A00404:156:HV37TDSXX:3:1533:16848:13479 chr17 543959 N chr17 544140 N DUP 1
A00404:155:HV27LDSXX:4:2233:6451:4617 chr16 28666312 N chr16 28666363 N DEL 15
A00404:155:HV27LDSXX:4:1431:17987:4272 chr4 24773641 N chr4 24773714 N DEL 5
A00404:155:HV27LDSXX:4:1431:18159:4445 chr4 24773641 N chr4 24773714 N DEL 5
A00404:156:HV37TDSXX:1:2378:7419:30029 chr4 24773641 N chr4 24773714 N DEL 5
A00404:156:HV37TDSXX:4:2645:24903:7858 chr4 24773645 N chr4 24773718 N DEL 5
A00404:156:HV37TDSXX:4:2170:6198:24220 chr4 24773647 N chr4 24773720 N DEL 5
A00404:155:HV27LDSXX:4:2253:19687:5368 chr8 29321092 N chr8 29321156 N DEL 15
A00404:155:HV27LDSXX:4:1361:12138:30248 chr1 143206632 N chr1 143206702 N DEL 10
A00404:155:HV27LDSXX:1:1378:14027:14669 chr1 143206529 N chr1 143206603 N DUP 5
A00404:156:HV37TDSXX:3:1544:31819:1329 chr1 143206335 N chr1 143206796 N DEL 2
A00404:155:HV27LDSXX:2:2618:11731:21934 chr1 143206543 N chr1 143206619 N DEL 3
A00404:155:HV27LDSXX:1:2103:12554:20134 chr1 143206334 N chr1 143206675 N DEL 5
A00297:158:HT275DSXX:1:2177:29930:27273 chr1 143206320 N chr1 143206707 N DEL 5
A00404:156:HV37TDSXX:1:1508:30698:1642 chr1 143206682 N chr1 143206754 N DEL 11
A00404:156:HV37TDSXX:4:2633:1063:25755 chr1 143206547 N chr1 143206690 N DUP 5
A00404:156:HV37TDSXX:4:2652:30969:8093 chr1 143206334 N chr1 143206387 N DEL 2
A00404:155:HV27LDSXX:2:1263:5828:32784 chr1 143206422 N chr1 143206686 N DUP 4
A00404:155:HV27LDSXX:3:1174:12246:21449 chr1 143206351 N chr1 143206810 N DUP 2
A00404:155:HV27LDSXX:4:2509:7048:32424 chr1 143206289 N chr1 143206702 N DEL 5
A00404:155:HV27LDSXX:2:1631:12852:6684 chr1 143206349 N chr1 143206713 N DEL 1
A00404:155:HV27LDSXX:2:2465:14145:11083 chr1 143206682 N chr1 143206754 N DEL 5
A00297:158:HT275DSXX:1:2570:3821:19820 chr1 143206288 N chr1 143206701 N DEL 5
A00404:156:HV37TDSXX:1:1260:5692:25535 chr1 143206438 N chr1 143206704 N DEL 5
A00404:156:HV37TDSXX:3:1568:26901:12352 chr1 143206273 N chr1 143206491 N DUP 2
A00404:155:HV27LDSXX:4:2443:27326:21324 chr1 143206529 N chr1 143206603 N DUP 5
A00404:155:HV27LDSXX:4:2331:11550:12007 chr1 143206347 N chr1 143206688 N DEL 7
A00404:155:HV27LDSXX:1:1433:16776:18082 chr1 143206334 N chr1 143206387 N DEL 57
A00404:155:HV27LDSXX:4:1113:13386:15154 chr1 143206529 N chr1 143206603 N DUP 5
A00297:158:HT275DSXX:2:2177:27597:3724 chr1 143206334 N chr1 143206606 N DEL 5
A00404:156:HV37TDSXX:4:1207:31810:16219 chr1 143206438 N chr1 143206704 N DEL 5
A00404:155:HV27LDSXX:3:1147:20817:11929 chr1 143206438 N chr1 143206704 N DEL 5
A00404:155:HV27LDSXX:4:1440:24451:16438 chr1 143206438 N chr1 143206704 N DEL 5
A00297:158:HT275DSXX:4:2332:1362:26741 chr1 143206320 N chr1 143206707 N DEL 5
A00404:155:HV27LDSXX:1:1144:12698:6856 chr1 143206311 N chr1 143206387 N DEL 26
A00404:156:HV37TDSXX:4:2520:28637:3396 chr1 143206335 N chr1 143206674 N DUP 5
A00297:158:HT275DSXX:3:2121:21224:4178 chr2 112889388 N chr2 112889523 N DEL 55
A00404:155:HV27LDSXX:4:1537:28185:21746 chr4 52464677 N chr4 52465027 N DEL 12
A00297:158:HT275DSXX:2:1524:12789:24424 chr4 52465169 N chr4 52465258 N DUP 7
A00404:156:HV37TDSXX:3:2527:19289:27195 chr9 134977402 N chr9 134977531 N DEL 5
A00404:156:HV37TDSXX:3:1107:5990:15342 chr9 134977402 N chr9 134977531 N DEL 5
A00404:156:HV37TDSXX:1:2538:2266:13839 chr9 134977402 N chr9 134977531 N DEL 5
A00297:158:HT275DSXX:4:1668:25771:22388 chr9 134977404 N chr9 134977461 N DEL 7
A00404:156:HV37TDSXX:3:1224:8657:8312 chr9 134977404 N chr9 134977461 N DEL 14
A00297:158:HT275DSXX:4:2620:25473:23750 chr9 134977404 N chr9 134977461 N DEL 10
A00297:158:HT275DSXX:4:1157:11605:33520 chr9 134977411 N chr9 134977506 N DUP 22
A00404:155:HV27LDSXX:1:2364:29324:7936 chr9 134977428 N chr9 134977485 N DUP 15
A00297:158:HT275DSXX:4:2620:25473:23750 chr9 134977367 N chr9 134977438 N DEL 2
A00404:156:HV37TDSXX:3:2347:25925:10441 chr9 134977365 N chr9 134977436 N DEL 4
A00404:156:HV37TDSXX:2:1242:29577:5556 chr9 134977417 N chr9 134977478 N DEL 5
A00404:155:HV27LDSXX:4:2243:3549:32628 chr9 134977540 N chr9 134977657 N DEL 5
A00404:156:HV37TDSXX:3:1643:30300:10097 chr17 82176327 N chr17 82176412 N DEL 4
A00404:155:HV27LDSXX:3:2149:15763:13135 chr20 61562135 N chr20 61562324 N DEL 5
A00404:155:HV27LDSXX:4:1173:1108:7357 chr20 61562136 N chr20 61562419 N DEL 10
A00404:155:HV27LDSXX:1:2218:5430:23202 chr20 61562187 N chr20 61562470 N DEL 10
A00404:155:HV27LDSXX:4:2255:7075:15060 chr20 61562323 N chr20 61562514 N DEL 10
A00404:155:HV27LDSXX:1:2303:25997:35336 chr20 61562177 N chr20 61562318 N DEL 6
A00404:156:HV37TDSXX:4:2307:26124:6402 chr20 61562370 N chr20 61562465 N DEL 9
A00404:156:HV37TDSXX:4:2271:5032:10645 chr20 61562370 N chr20 61562465 N DEL 9
A00404:156:HV37TDSXX:2:1637:14479:33739 chr20 61562370 N chr20 61562465 N DEL 9
A00404:155:HV27LDSXX:2:2411:32289:28322 chr20 61562370 N chr20 61562465 N DEL 9
A00404:155:HV27LDSXX:4:1557:16966:33254 chr20 61562133 N chr20 61562416 N DEL 9
A00404:155:HV27LDSXX:3:2149:15763:13135 chr20 61562133 N chr20 61562416 N DEL 9
A00404:155:HV27LDSXX:1:2516:23086:35430 chr20 61562165 N chr20 61562400 N DEL 9
A00297:158:HT275DSXX:3:1376:3974:5932 chr20 61562165 N chr20 61562400 N DEL 9
A00297:158:HT275DSXX:4:1421:30671:35571 chr20 61562173 N chr20 61562408 N DEL 7
A00404:156:HV37TDSXX:2:1534:10104:5869 chr20 61562322 N chr20 61562465 N DEL 5
A00404:156:HV37TDSXX:2:1534:9661:6511 chr20 61562322 N chr20 61562465 N DEL 5
A00404:156:HV37TDSXX:4:2474:10691:16720 chr20 61562322 N chr20 61562465 N DEL 5
A00404:156:HV37TDSXX:4:2474:12680:16783 chr20 61562322 N chr20 61562465 N DEL 5
A00404:156:HV37TDSXX:4:2631:18973:28338 chr20 61562322 N chr20 61562465 N DEL 5
A00297:158:HT275DSXX:1:2536:4336:5243 chr20 61562322 N chr20 61562465 N DEL 5
A00404:156:HV37TDSXX:4:1108:19913:1908 chr20 61562322 N chr20 61562465 N DEL 5
A00297:158:HT275DSXX:4:2152:31394:36292 chr20 61562243 N chr20 61562478 N DEL 2
A00297:158:HT275DSXX:1:2309:23194:36338 chr8 1022407 N chr8 1022463 N DEL 11
A00297:158:HT275DSXX:1:2512:21323:1031 chr8 1022336 N chr8 1022445 N DUP 5
A00404:155:HV27LDSXX:2:2475:18909:24283 chr8 1022377 N chr8 1022486 N DUP 12
A00404:156:HV37TDSXX:3:2576:23818:2033 chr8 1022456 N chr8 1022510 N DUP 5
A00297:158:HT275DSXX:1:2309:23194:36338 chr8 1022317 N chr8 1022483 N DEL 5
A00404:155:HV27LDSXX:3:1514:29848:22341 chr8 1022594 N chr8 1022705 N DEL 5
A00404:156:HV37TDSXX:4:2523:11984:27665 chr8 1022590 N chr8 1022866 N DEL 15
A00404:155:HV27LDSXX:2:1660:19108:2425 chr8 1022345 N chr8 1022566 N DEL 25
A00404:155:HV27LDSXX:1:2348:1814:10019 chr8 1022345 N chr8 1022566 N DEL 8
A00404:156:HV37TDSXX:4:2228:11605:4304 chr8 1022497 N chr8 1022608 N DEL 5
A00404:155:HV27LDSXX:3:1514:29848:22341 chr8 1022528 N chr8 1022859 N DEL 5
A00404:155:HV27LDSXX:3:1657:5222:19210 chr8 1022428 N chr8 1022869 N DEL 14
A00297:158:HT275DSXX:3:1223:19280:32158 chr8 1022458 N chr8 1022899 N DEL 20
A00297:158:HT275DSXX:1:1403:5810:34131 chr8 1022601 N chr8 1022932 N DEL 37
A00404:155:HV27LDSXX:3:2644:32669:19366 chr8 1022632 N chr8 1022908 N DEL 9
A00297:158:HT275DSXX:4:2424:10890:10989 chr10 45033075 N chr10 45033263 N DEL 45
A00297:158:HT275DSXX:4:2320:16089:17926 chr19 56444588 N chr19 56445004 N DEL 5
A00404:156:HV37TDSXX:2:1568:23204:3975 chr19 56444588 N chr19 56444755 N DEL 2
A00404:156:HV37TDSXX:1:1157:12590:36980 chr19 56444749 N chr19 56444999 N DEL 5
A00404:155:HV27LDSXX:3:1520:4372:24502 chr19 56444721 N chr19 56444804 N DEL 1
A00404:155:HV27LDSXX:1:1241:19678:24799 chr19 56444945 N chr19 56445359 N DUP 2
A00404:156:HV37TDSXX:2:1241:10511:26146 chr19 56445373 N chr19 56445455 N DUP 5
A00404:156:HV37TDSXX:1:1575:15863:21167 chr19 56444708 N chr19 56444875 N DEL 5
A00297:158:HT275DSXX:4:1601:7961:5040 chr19 56444928 N chr19 56445261 N DEL 5
A00404:155:HV27LDSXX:4:2450:4625:21465 chr19 56444752 N chr19 56445251 N DEL 3
A00297:158:HT275DSXX:2:2249:3676:21731 chr19 56444928 N chr19 56445261 N DEL 5
A00297:158:HT275DSXX:3:1569:3233:23312 chr19 56445373 N chr19 56445455 N DUP 5
A00297:158:HT275DSXX:3:1126:4092:11177 chr19 56444877 N chr19 56445458 N DUP 5
A00297:158:HT275DSXX:1:1220:9227:11898 chr12 127696670 N chr12 127696799 N DEL 35
A00404:155:HV27LDSXX:1:2461:22824:33599 chr12 127696640 N chr12 127696768 N DEL 29
A00404:155:HV27LDSXX:2:1661:28212:33285 chr12 127696670 N chr12 127696799 N DEL 35
A00404:156:HV37TDSXX:1:2235:6352:3505 chr12 127696670 N chr12 127696799 N DEL 35
A00404:155:HV27LDSXX:4:1625:31792:27211 chr12 127696670 N chr12 127696799 N DEL 35
A00404:156:HV37TDSXX:2:1163:10619:2910 chr12 127696670 N chr12 127696799 N DEL 29
A00404:156:HV37TDSXX:4:2105:31250:23234 chr12 127696670 N chr12 127696799 N DEL 17
A00404:155:HV27LDSXX:2:2277:13883:25535 chr12 127696670 N chr12 127696799 N DEL 16
A00297:158:HT275DSXX:2:1161:7383:35383 chr12 127696670 N chr12 127696799 N DEL 12
A00404:155:HV27LDSXX:1:2673:30626:20369 chr12 127696670 N chr12 127696799 N DEL 19
A00404:156:HV37TDSXX:4:2105:30761:22326 chr12 127696670 N chr12 127696799 N DEL 14
A00404:155:HV27LDSXX:4:2503:1551:8844 chr12 127696670 N chr12 127696799 N DEL 7
A00404:155:HV27LDSXX:4:1226:6225:2002 chr12 127696670 N chr12 127696799 N DEL 6
A00404:156:HV37TDSXX:3:1264:20799:1376 chr12 127696670 N chr12 127696799 N DEL 6
A00297:158:HT275DSXX:1:1624:26015:8155 chr12 127696671 N chr12 127696800 N DEL 6
A00297:158:HT275DSXX:1:1625:26657:6480 chr12 127696671 N chr12 127696800 N DEL 6
A00297:158:HT275DSXX:1:2626:22860:2910 chr12 127696671 N chr12 127696800 N DEL 6
A00404:156:HV37TDSXX:2:2353:32597:25473 chr12 127696675 N chr12 127696804 N DEL 6
A00404:155:HV27LDSXX:1:2223:17743:33786 chr12 127696682 N chr12 127696811 N DEL 1
A00297:158:HT275DSXX:1:1307:22345:31109 chr4 186509612 N chr4 186509675 N DUP 5
A00297:158:HT275DSXX:1:1307:22571:31250 chr4 186509612 N chr4 186509675 N DUP 5
A00404:155:HV27LDSXX:1:1633:29270:27445 chr4 186509612 N chr4 186509675 N DUP 13
A00404:156:HV37TDSXX:2:2558:22770:18599 chr14 71544084 N chr14 71544155 N DEL 5
A00404:156:HV37TDSXX:4:1501:16984:7200 chr14 71544084 N chr14 71544155 N DEL 5
A00404:156:HV37TDSXX:4:1501:17815:7451 chr14 71544084 N chr14 71544155 N DEL 5
A00404:156:HV37TDSXX:2:1159:10700:15608 chr14 71543993 N chr14 71544052 N DEL 18
A00297:158:HT275DSXX:2:2456:32687:4492 chr14 71543993 N chr14 71544052 N DEL 14
A00297:158:HT275DSXX:4:1117:9173:1125 chr14 71543993 N chr14 71544052 N DEL 14
A00404:155:HV27LDSXX:3:1228:13621:19038 chr14 71543996 N chr14 71544055 N DEL 12
A00297:158:HT275DSXX:2:2556:25102:23202 chr14 71543980 N chr14 71544066 N DEL 1
A00404:156:HV37TDSXX:2:1643:27037:9173 chr14 71543999 N chr14 71544058 N DEL 9
A00404:155:HV27LDSXX:3:2575:12635:17832 chr14 71543999 N chr14 71544058 N DEL 9
A00297:158:HT275DSXX:4:1347:30644:6308 chr14 71544102 N chr14 71544171 N DUP 5
A00404:155:HV27LDSXX:2:1242:28791:13369 chr14 71544102 N chr14 71544171 N DUP 5
A00404:155:HV27LDSXX:2:1242:28791:13463 chr14 71544102 N chr14 71544171 N DUP 5
A00404:155:HV27LDSXX:4:2468:20980:15374 chr14 71544104 N chr14 71544173 N DUP 5
A00404:155:HV27LDSXX:3:1229:5882:9142 chr14 71544107 N chr14 71544176 N DUP 5
A00297:158:HT275DSXX:1:1662:13973:13197 chr1 192115174 N chr1 192115242 N DEL 2
A00297:158:HT275DSXX:1:1671:2564:2769 chr1 192115174 N chr1 192115242 N DEL 2
A00404:155:HV27LDSXX:3:1444:10800:28056 chr15 84889788 N chr15 84889939 N DEL 5
A00404:155:HV27LDSXX:1:1230:23809:10160 chr15 84889788 N chr15 84889939 N DEL 5
A00297:158:HT275DSXX:3:2424:26720:27602 chr15 84889823 N chr15 84889956 N DUP 17
A00404:155:HV27LDSXX:3:1273:26865:10285 chr15 84889823 N chr15 84889956 N DUP 17
A00404:156:HV37TDSXX:3:1131:20320:6370 chr15 84889823 N chr15 84889956 N DUP 16
A00404:156:HV37TDSXX:2:2209:27353:34053 chr15 84889823 N chr15 84889956 N DUP 16
A00297:158:HT275DSXX:2:2269:15203:20243 chr15 84889823 N chr15 84889956 N DUP 15
A00404:156:HV37TDSXX:2:2572:30716:12352 chr15 84889824 N chr15 84889957 N DUP 14
A00404:155:HV27LDSXX:2:2451:13657:28808 chrX 102412643 N chrX 102412747 N DEL 10
A00404:155:HV27LDSXX:2:1437:15058:11757 chrX 102412642 N chrX 102412758 N DEL 1
A00297:158:HT275DSXX:2:2226:13376:23657 chrX 102412678 N chrX 102412797 N DEL 5
A00404:155:HV27LDSXX:3:2524:25690:9408 chrX 102412660 N chrX 102412797 N DEL 5
A00404:156:HV37TDSXX:4:2248:30951:23187 chr2 1099739 N chr2 1099818 N DUP 12
A00404:156:HV37TDSXX:4:2248:31204:22968 chr2 1099739 N chr2 1099818 N DUP 12
A00404:155:HV27LDSXX:3:1370:3983:16595 chr6 170453167 N chr6 170453303 N DEL 4
A00404:155:HV27LDSXX:4:1675:29803:21699 chr6 170453217 N chr6 170453343 N DUP 5
A00404:155:HV27LDSXX:1:1155:22263:18161 chr16 36175570 N chr16 36175953 N DUP 11
A00297:158:HT275DSXX:1:2228:3224:5196 chr16 36175727 N chr16 36175897 N DEL 5
A00404:155:HV27LDSXX:2:1222:31620:3834 chr4 713379 N chr4 713505 N DEL 26
A00297:158:HT275DSXX:4:1512:12138:23202 chr4 713371 N chr4 713497 N DEL 5
A00404:155:HV27LDSXX:4:1478:11460:23563 chr4 713370 N chr4 713496 N DEL 5
A00404:156:HV37TDSXX:4:1652:1253:6136 chr4 713370 N chr4 713496 N DEL 5
A00297:158:HT275DSXX:4:2340:4110:7795 chr4 713341 N chr4 713503 N DEL 5
A00404:156:HV37TDSXX:1:2324:18683:20134 chr4 713355 N chr4 713552 N DEL 5
A00404:155:HV27LDSXX:3:1372:7681:3740 chr4 713330 N chr4 713580 N DEL 5
A00297:158:HT275DSXX:4:1355:13865:18865 chr4 713347 N chr4 713702 N DUP 10
A00404:155:HV27LDSXX:1:1416:21567:6809 chr4 713361 N chr4 713701 N DEL 13
A00404:155:HV27LDSXX:1:1557:3378:17832 chr4 713361 N chr4 713701 N DEL 13
A00297:158:HT275DSXX:3:1544:7491:20791 chr4 713367 N chr4 713707 N DEL 7
A00404:156:HV37TDSXX:4:1543:5484:2660 chr4 713366 N chr4 713706 N DEL 8
A00297:158:HT275DSXX:3:1116:3269:4586 chr2 3416623 N chr2 3416976 N DEL 26
A00404:156:HV37TDSXX:4:1423:30309:17816 chr2 3416623 N chr2 3416765 N DEL 27
A00297:158:HT275DSXX:2:1557:24243:19617 chr2 3416697 N chr2 3417000 N DUP 5
A00297:158:HT275DSXX:2:2151:31268:10144 chr2 3416698 N chr2 3416931 N DUP 5
A00404:155:HV27LDSXX:4:2525:3179:32205 chr2 3416781 N chr2 3416852 N DEL 3
A00404:155:HV27LDSXX:3:1649:26747:31908 chr2 3416850 N chr2 3416919 N DUP 5
A00404:155:HV27LDSXX:4:2632:30101:15201 chr2 3416676 N chr2 3416911 N DEL 5
A00404:155:HV27LDSXX:1:1228:28619:17926 chr2 3416783 N chr2 3417088 N DUP 8
A00297:158:HT275DSXX:1:2223:19316:5071 chr19 40396829 N chr19 40396986 N DEL 13
A00404:155:HV27LDSXX:2:1250:14290:31469 chr19 40396934 N chr19 40397013 N DEL 5
A00404:155:HV27LDSXX:3:1222:26910:19006 chr21 8404001 N chr21 8404086 N DUP 12
A00404:156:HV37TDSXX:2:1121:20112:10300 chr21 8403932 N chr21 8403997 N DEL 13
A00297:158:HT275DSXX:4:2272:19126:3991 chr21 8403932 N chr21 8403997 N DEL 12
A00297:158:HT275DSXX:4:1642:10664:26193 chr21 8403983 N chr21 8404038 N DEL 12
A00404:155:HV27LDSXX:3:2339:3161:10191 chr21 8404020 N chr21 8404089 N DUP 16
A00297:158:HT275DSXX:3:1249:14913:19022 chr21 8403989 N chr21 8404056 N DEL 5
A00297:158:HT275DSXX:4:2553:15130:23531 chr21 8403993 N chr21 8404054 N DEL 5
A00404:155:HV27LDSXX:3:2251:6171:12555 chr21 8403976 N chr21 8404093 N DEL 5
A00404:155:HV27LDSXX:1:2231:6045:27305 chr21 8403975 N chr21 8404038 N DEL 13
A00404:156:HV37TDSXX:1:1328:21956:1783 chr21 8403974 N chr21 8404051 N DUP 1
A00297:158:HT275DSXX:3:1174:7997:3161 chr21 8404038 N chr21 8404091 N DUP 18
A00404:155:HV27LDSXX:1:1342:1054:6230 chr21 8403975 N chr21 8404044 N DEL 5
A00404:155:HV27LDSXX:3:2575:31955:27430 chr21 8403975 N chr21 8404042 N DEL 6
A00404:156:HV37TDSXX:1:1338:15474:3333 chr21 8403976 N chr21 8404037 N DUP 4
A00404:155:HV27LDSXX:4:2230:13566:24048 chr21 8403911 N chr21 8404044 N DUP 9
A00404:156:HV37TDSXX:1:2136:10393:22592 chr21 8403975 N chr21 8404048 N DEL 5
A00297:158:HT275DSXX:1:2443:8901:1470 chr21 8403980 N chr21 8404093 N DEL 5
A00297:158:HT275DSXX:2:2468:18204:25066 chr21 8403987 N chr21 8404048 N DEL 10
A00297:158:HT275DSXX:1:2538:25427:16877 chr21 8403953 N chr21 8404038 N DEL 21
A00404:156:HV37TDSXX:1:2105:29550:6793 chr21 8403963 N chr21 8404018 N DUP 15
A00404:156:HV37TDSXX:2:1618:5737:18693 chr21 8403911 N chr21 8404028 N DUP 11
A00297:158:HT275DSXX:1:2540:32172:16438 chr21 8403975 N chr21 8404046 N DEL 5
A00297:158:HT275DSXX:4:1123:12237:8500 chr21 8403857 N chr21 8403906 N DUP 15
A00404:155:HV27LDSXX:2:2276:23484:16297 chr21 8403975 N chr21 8404042 N DEL 6
A00404:156:HV37TDSXX:1:2163:27724:33786 chr21 8403976 N chr21 8404037 N DUP 5
A00404:156:HV37TDSXX:3:2132:14751:8563 chr21 8403978 N chr21 8404027 N DUP 5
A00404:155:HV27LDSXX:1:2627:1723:16626 chr21 8403975 N chr21 8404030 N DEL 10
A00297:158:HT275DSXX:3:2319:26169:5697 chr8 141998184 N chr8 141998332 N DUP 5
A00404:156:HV37TDSXX:1:2644:9607:2785 chr8 141998258 N chr8 141998460 N DEL 29
A00404:156:HV37TDSXX:4:2509:26756:22122 chr22 21913093 N chr22 21913147 N DEL 2
A00404:155:HV27LDSXX:4:1467:27335:2268 chr5 9162544 N chr5 9162605 N DUP 8
A00404:156:HV37TDSXX:1:2523:23023:4476 chr5 9162620 N chr5 9162729 N DEL 31
A00404:156:HV37TDSXX:4:1473:12979:32424 chr16 49002317 N chr16 49002453 N DEL 8
A00297:158:HT275DSXX:3:2260:11143:26522 chr16 49002318 N chr16 49002454 N DEL 7
A00404:155:HV27LDSXX:4:1117:25970:25895 chr11 50229005 N chr11 50229061 N DEL 5
A00404:156:HV37TDSXX:3:2276:26521:33332 chr2 41748075 N chr2 41748249 N DUP 1
A00297:158:HT275DSXX:2:1118:10330:23985 chr22 49999787 N chr22 49999869 N DEL 6
A00297:158:HT275DSXX:2:1118:10610:22748 chr22 49999787 N chr22 49999869 N DEL 6
A00297:158:HT275DSXX:2:1118:10610:22780 chr22 49999787 N chr22 49999869 N DEL 6
A00297:158:HT275DSXX:1:1434:19271:26537 chr22 49999787 N chr22 49999869 N DEL 6
A00404:155:HV27LDSXX:3:1375:30355:15170 chr22 49999787 N chr22 49999869 N DEL 6
A00404:156:HV37TDSXX:4:1669:31801:18239 chr22 49999787 N chr22 49999869 N DEL 6
A00404:156:HV37TDSXX:2:1437:11044:10003 chr22 49999796 N chr22 49999894 N DEL 7
A00404:155:HV27LDSXX:3:1254:3513:12461 chr6 135363733 N chr6 135364126 N DEL 5
A00404:155:HV27LDSXX:4:1572:10872:20196 chr6 135363806 N chr6 135363895 N DUP 12
A00297:158:HT275DSXX:3:2430:2239:28635 chr6 135363984 N chr6 135364162 N DEL 21
A00404:155:HV27LDSXX:2:1309:13711:34100 chr6 135363769 N chr6 135363985 N DEL 5
A00404:156:HV37TDSXX:3:1357:26377:21308 chr6 135363811 N chr6 135364027 N DEL 5
A00404:156:HV37TDSXX:1:1170:14226:33771 chr6 135363817 N chr6 135364210 N DEL 2
A00297:158:HT275DSXX:4:1643:24894:29011 chr6 135364057 N chr6 135364234 N DEL 4
A00404:156:HV37TDSXX:2:2145:19949:18035 chr10 129992477 N chr10 129992538 N DEL 17
A00404:155:HV27LDSXX:2:1361:3667:12853 chr4 11565906 N chr4 11566034 N DEL 5
A00404:156:HV37TDSXX:2:2323:19831:18677 chr4 176723501 N chr4 176723710 N DEL 10
A00404:156:HV37TDSXX:2:2323:19831:18677 chr4 176723545 N chr4 176723615 N DEL 5
A00297:158:HT275DSXX:3:1422:25635:2769 chr4 176723577 N chr4 176723665 N DUP 5
A00404:155:HV27LDSXX:4:1348:29161:10160 chr4 176723568 N chr4 176723656 N DUP 5
A00404:155:HV27LDSXX:1:2175:8314:3583 chr4 176723568 N chr4 176723656 N DUP 5
A00404:156:HV37TDSXX:4:2518:26377:27539 chr4 176723568 N chr4 176723656 N DUP 5
A00297:158:HT275DSXX:1:1450:10194:35556 chr4 176723568 N chr4 176723656 N DUP 5
A00404:155:HV27LDSXX:2:2670:32786:29684 chr2 129654469 N chr2 129654659 N DEL 10
A00404:156:HV37TDSXX:1:1336:8015:22106 chr2 129654853 N chr2 129655291 N DEL 16
A00404:155:HV27LDSXX:2:2202:27633:2566 chr2 129654847 N chr2 129655222 N DEL 11
A00404:156:HV37TDSXX:3:2465:10981:12023 chr2 129654581 N chr2 129654873 N DEL 5
A00404:156:HV37TDSXX:3:2465:11035:11866 chr2 129654572 N chr2 129654864 N DEL 5
A00404:155:HV27LDSXX:1:1425:2103:13808 chr2 129654968 N chr2 129655217 N DEL 10
A00404:155:HV27LDSXX:1:2321:26323:31485 chr2 129654991 N chr2 129655240 N DEL 4
A00404:156:HV37TDSXX:2:2137:24758:32753 chr2 129654991 N chr2 129655240 N DEL 5
A00404:155:HV27LDSXX:1:2336:9227:6950 chr2 129654902 N chr2 129655090 N DUP 5
A00404:156:HV37TDSXX:2:2476:22661:28808 chr2 129654675 N chr2 129655091 N DUP 5
A00404:155:HV27LDSXX:4:2377:26892:3349 chr2 129654675 N chr2 129655091 N DUP 5
A00297:158:HT275DSXX:2:1503:13376:25598 chr2 129655102 N chr2 129655350 N DEL 5
A00297:158:HT275DSXX:2:2433:7274:28839 chr2 129654695 N chr2 129655113 N DEL 5
A00404:156:HV37TDSXX:2:2516:19379:24972 chr2 129654571 N chr2 129655115 N DEL 5
A00404:156:HV37TDSXX:1:1421:4273:34601 chr2 129655167 N chr2 129655229 N DUP 1
A00404:155:HV27LDSXX:2:1605:7175:26475 chr2 129654438 N chr2 129655167 N DEL 7
A00404:155:HV27LDSXX:2:1659:20383:19852 chr2 129654960 N chr2 129655209 N DEL 14
A00404:156:HV37TDSXX:3:2527:25102:24142 chr2 129655090 N chr2 129655339 N DEL 5
A00404:156:HV37TDSXX:2:2511:29559:27445 chr2 129654948 N chr2 129655385 N DEL 20
A00404:156:HV37TDSXX:4:1606:16134:21981 chr2 129654958 N chr2 129655395 N DEL 5
A00404:155:HV27LDSXX:2:1603:4435:36542 chr7 157433346 N chr7 157433467 N DUP 5
A00404:155:HV27LDSXX:1:2416:22101:22106 chr7 157433333 N chr7 157433490 N DUP 2
A00297:158:HT275DSXX:2:2302:30264:33144 chr7 157433333 N chr7 157433490 N DUP 5
A00404:155:HV27LDSXX:4:2229:23448:8406 chr3 133416977 N chr3 133417118 N DEL 5
A00404:155:HV27LDSXX:2:1602:19434:20494 chr3 133417266 N chr3 133417324 N DUP 5
A00404:155:HV27LDSXX:3:1420:32362:21652 chr3 133417642 N chr3 133418304 N DUP 5
A00404:156:HV37TDSXX:1:2108:8377:33974 chr3 133417482 N chr3 133417859 N DUP 5
A00404:155:HV27LDSXX:3:1425:14335:7122 chr3 133417047 N chr3 133417860 N DUP 5
A00404:156:HV37TDSXX:3:2305:18873:18082 chr3 133417095 N chr3 133418254 N DEL 6
A00404:156:HV37TDSXX:1:2159:16776:11757 chr3 133417809 N chr3 133418272 N DEL 4
A00404:156:HV37TDSXX:3:2245:7898:32643 chr4 172606760 N chr4 172606829 N DEL 27
A00404:155:HV27LDSXX:3:2434:31313:17300 chr4 172606760 N chr4 172606829 N DEL 37
A00404:155:HV27LDSXX:3:2142:1533:16861 chr4 172606760 N chr4 172606829 N DEL 25
A00404:155:HV27LDSXX:3:1653:24316:16203 chr10 148360 N chr10 148501 N DEL 3
A00297:158:HT275DSXX:3:2467:24668:35978 chr10 148360 N chr10 148501 N DEL 4
A00297:158:HT275DSXX:3:1212:11785:14606 chr10 148360 N chr10 148501 N DEL 5
A00404:156:HV37TDSXX:1:2270:18159:9768 chr10 148360 N chr10 148501 N DEL 5
A00297:158:HT275DSXX:3:2375:6524:29387 chr10 148360 N chr10 148501 N DEL 5
A00297:158:HT275DSXX:1:1548:31991:4006 chr10 148360 N chr10 148501 N DEL 5
A00297:158:HT275DSXX:4:1139:17662:23594 chr10 148360 N chr10 148501 N DEL 5
A00297:158:HT275DSXX:4:2204:2302:12054 chr10 148360 N chr10 148501 N DEL 5
A00297:158:HT275DSXX:3:1463:7844:13636 chr10 148360 N chr10 148501 N DEL 5
A00404:156:HV37TDSXX:1:2673:29405:17566 chr10 148365 N chr10 148560 N DUP 5
A00297:158:HT275DSXX:2:2311:28718:20102 chr10 148365 N chr10 148560 N DUP 5
A00404:155:HV27LDSXX:3:1676:24406:24283 chr10 148365 N chr10 148560 N DUP 5
A00404:155:HV27LDSXX:1:1624:24198:25801 chr10 148365 N chr10 148560 N DUP 5
A00404:155:HV27LDSXX:4:2159:14055:25081 chr10 148365 N chr10 148560 N DUP 5
A00297:158:HT275DSXX:3:1525:6759:33301 chr10 148365 N chr10 148560 N DUP 5
A00297:158:HT275DSXX:3:1525:6768:33317 chr10 148365 N chr10 148560 N DUP 5
A00297:158:HT275DSXX:2:1229:24216:5697 chr10 148365 N chr10 148560 N DUP 5
A00404:156:HV37TDSXX:4:1425:23547:30906 chr10 148428 N chr10 148567 N DUP 5
A00297:158:HT275DSXX:1:1407:12328:14794 chr10 148435 N chr10 148574 N DUP 1
A00404:155:HV27LDSXX:2:2167:9453:5118 chr2 3304756 N chr2 3304870 N DUP 35
A00404:155:HV27LDSXX:3:1366:26124:20619 chr2 3304756 N chr2 3304870 N DUP 30
A00404:155:HV27LDSXX:3:1366:27959:20791 chr2 3304756 N chr2 3304870 N DUP 30
A00404:156:HV37TDSXX:3:2143:21748:29074 chr2 3304756 N chr2 3304870 N DUP 21
A00297:158:HT275DSXX:2:2638:4661:31140 chr2 3304769 N chr2 3304883 N DUP 2
A00297:158:HT275DSXX:3:1339:29993:32236 chr2 3304763 N chr2 3304877 N DUP 8
A00404:156:HV37TDSXX:1:2410:31575:16344 chr2 3304764 N chr2 3304878 N DUP 4
A00297:158:HT275DSXX:4:1662:18059:1736 chr2 3304767 N chr2 3304881 N DUP 5
A00404:155:HV27LDSXX:2:2235:13132:3975 chr8 141347693 N chr8 141347760 N DEL 9
A00404:155:HV27LDSXX:2:1371:1163:18067 chr8 141347701 N chr8 141347760 N DEL 10
A00404:156:HV37TDSXX:4:2520:8612:4288 chr8 141347701 N chr8 141347760 N DEL 10
A00404:155:HV27LDSXX:1:1349:12264:9111 chr8 141347693 N chr8 141347760 N DEL 44
A00297:158:HT275DSXX:3:2633:22652:13009 chr8 141347693 N chr8 141347760 N DEL 44
A00297:158:HT275DSXX:1:1504:31096:14669 chr8 141347701 N chr8 141347760 N DEL 41
A00404:156:HV37TDSXX:4:2203:29586:14998 chr8 141347701 N chr8 141347760 N DEL 41
A00404:155:HV27LDSXX:2:1617:10728:22106 chr5 181444915 N chr5 181444989 N DEL 17
A00404:155:HV27LDSXX:3:1575:15510:5274 chr7 69850433 N chr7 69850538 N DEL 2
A00404:156:HV37TDSXX:1:2344:25672:25285 chr7 69850433 N chr7 69850538 N DEL 5
A00404:156:HV37TDSXX:2:1565:18394:21887 chr20 55967536 N chr20 55967723 N DUP 10
A00404:155:HV27LDSXX:1:1673:1163:25708 chr20 55967572 N chr20 55967637 N DUP 20
A00404:156:HV37TDSXX:3:2520:28619:1204 chr20 55967572 N chr20 55967637 N DUP 24
A00297:158:HT275DSXX:1:1554:20139:12978 chr20 55967583 N chr20 55967660 N DUP 3
A00297:158:HT275DSXX:4:1251:25563:21120 chr20 55967572 N chr20 55967703 N DUP 7
A00404:155:HV27LDSXX:1:1511:7500:23938 chr20 55967572 N chr20 55967703 N DUP 7
A00404:156:HV37TDSXX:1:1667:22996:14262 chr20 55967572 N chr20 55967637 N DUP 15
A00404:155:HV27LDSXX:1:2535:14045:5838 chr20 55967572 N chr20 55967637 N DUP 25
A00404:155:HV27LDSXX:2:2149:10068:7936 chr20 55967572 N chr20 55967637 N DUP 16
A00404:155:HV27LDSXX:4:1148:2817:19617 chr20 55967572 N chr20 55967637 N DUP 25
A00404:155:HV27LDSXX:4:1447:24514:17206 chr20 55967578 N chr20 55967643 N DUP 20
A00404:155:HV27LDSXX:4:2130:31250:24862 chr20 55967572 N chr20 55967637 N DUP 22
A00404:156:HV37TDSXX:1:2309:22978:28322 chr20 55967572 N chr20 55967637 N DUP 15
A00404:156:HV37TDSXX:2:1638:29125:15734 chr20 55967573 N chr20 55967672 N DUP 10
A00404:156:HV37TDSXX:4:2241:27805:25285 chr20 55967572 N chr20 55967637 N DUP 27
A00404:155:HV27LDSXX:2:2411:13702:29512 chr20 55967573 N chr20 55967672 N DUP 10
A00404:156:HV37TDSXX:2:1303:18050:29183 chr20 55967578 N chr20 55967677 N DUP 10
A00404:156:HV37TDSXX:1:2155:30273:32972 chr20 55967573 N chr20 55967672 N DUP 11
A00404:156:HV37TDSXX:4:2127:23809:5838 chr20 55967573 N chr20 55967672 N DUP 13
A00404:156:HV37TDSXX:3:1442:16676:16250 chr20 55967572 N chr20 55967637 N DUP 16
A00404:155:HV27LDSXX:4:2529:11812:34100 chr20 55967572 N chr20 55967637 N DUP 16
A00404:155:HV27LDSXX:2:2441:2917:12900 chr20 55967572 N chr20 55967637 N DUP 18
A00404:156:HV37TDSXX:4:1452:20582:1188 chr20 55967619 N chr20 55967688 N DEL 22
A00297:158:HT275DSXX:2:1360:21649:20384 chr20 55967619 N chr20 55967688 N DEL 16
A00404:155:HV27LDSXX:2:1535:10601:8077 chr20 55967619 N chr20 55967688 N DEL 17
A00404:156:HV37TDSXX:1:2229:30734:9126 chr20 55967619 N chr20 55967688 N DEL 12
A00404:156:HV37TDSXX:2:1315:14751:15170 chr20 55967619 N chr20 55967688 N DEL 12
A00297:158:HT275DSXX:1:1644:6099:17722 chr20 55967619 N chr20 55967688 N DEL 11
A00297:158:HT275DSXX:3:2632:15176:22795 chr20 55967586 N chr20 55967699 N DEL 4
A00297:158:HT275DSXX:4:1274:28167:14105 chr20 55967554 N chr20 55967701 N DEL 2
A00404:156:HV37TDSXX:1:2351:19443:9580 chr11 21342816 N chr11 21342873 N DEL 14
A00404:156:HV37TDSXX:1:1350:1759:18881 chrX 828107 N chrX 828414 N DUP 5
A00297:158:HT275DSXX:3:2110:20871:2065 chrX 25905925 N chrX 25906122 N DEL 6
A00404:156:HV37TDSXX:1:1678:23348:24862 chrX 25906000 N chrX 25906362 N DEL 3
A00404:155:HV27LDSXX:4:2111:32217:16203 chrX 25906023 N chrX 25906383 N DUP 10
A00404:156:HV37TDSXX:2:1205:5972:11146 chrX 25906027 N chrX 25906108 N DEL 5
A00404:156:HV37TDSXX:3:2411:15248:24486 chrX 25906237 N chrX 25906323 N DUP 2
A00297:158:HT275DSXX:3:2652:3848:32111 chr8 6073099 N chr8 6073297 N DEL 11
A00297:158:HT275DSXX:1:2552:26006:19132 chr8 6073262 N chr8 6073369 N DUP 2
A00404:156:HV37TDSXX:3:2270:7518:32424 chr21 46364249 N chr21 46364443 N DEL 40
A00297:158:HT275DSXX:4:2505:19289:25379 chr21 46364291 N chr21 46364485 N DEL 10
A00297:158:HT275DSXX:1:2504:30138:8218 chr21 46364373 N chr21 46364503 N DEL 21
A00297:158:HT275DSXX:4:1246:17933:28228 chr21 46364423 N chr21 46364553 N DEL 49
A00297:158:HT275DSXX:1:1401:1904:1501 chr19 9443090 N chr19 9443407 N DEL 10
A00404:156:HV37TDSXX:3:1438:2410:3380 chr19 9443090 N chr19 9443407 N DEL 12
A00297:158:HT275DSXX:1:1460:8323:7576 chr19 9443228 N chr19 9443549 N DEL 13
A00297:158:HT275DSXX:4:1626:15402:2300 chr19 9443263 N chr19 9443584 N DEL 8
A00404:155:HV27LDSXX:3:1429:10899:10817 chr19 9443158 N chr19 9443475 N DEL 5
A00297:158:HT275DSXX:2:2250:19199:36746 chr19 9443317 N chr19 9443640 N DEL 2
A00297:158:HT275DSXX:1:1661:5150:22498 chrX 1278075 N chrX 1278432 N DEL 5
A00404:156:HV37TDSXX:3:1503:29306:2300 chrX 1278075 N chrX 1278432 N DEL 5
A00404:156:HV37TDSXX:3:1503:29342:2237 chrX 1278075 N chrX 1278432 N DEL 5
A00297:158:HT275DSXX:3:2336:1217:10363 chrX 1278075 N chrX 1278432 N DEL 5
A00404:156:HV37TDSXX:3:2370:6072:16705 chrX 1278075 N chrX 1278432 N DEL 5
A00404:156:HV37TDSXX:4:2550:28393:33912 chrX 1278075 N chrX 1278432 N DEL 5
A00404:156:HV37TDSXX:1:2631:24144:23422 chrX 1278075 N chrX 1278432 N DEL 5
A00297:158:HT275DSXX:1:2144:30689:4820 chrX 1278126 N chrX 1278834 N DUP 5
A00404:156:HV37TDSXX:3:2552:29161:9126 chrX 1278126 N chrX 1278834 N DUP 5
A00297:158:HT275DSXX:3:1121:2691:15828 chrX 1278106 N chrX 1278461 N DUP 5
A00404:155:HV27LDSXX:4:2545:29776:3646 chrX 1278192 N chrX 1278544 N DUP 10
A00404:156:HV37TDSXX:1:1638:12472:31266 chrX 1278192 N chrX 1278544 N DUP 10
A00404:156:HV37TDSXX:1:1638:12563:31140 chrX 1278192 N chrX 1278544 N DUP 10
A00404:156:HV37TDSXX:3:2139:4444:34147 chrX 1278192 N chrX 1278544 N DUP 10
A00404:156:HV37TDSXX:1:2654:27688:22357 chrX 1278192 N chrX 1278544 N DUP 10
A00404:155:HV27LDSXX:2:1440:16721:21746 chrX 1278192 N chrX 1278544 N DUP 10
A00297:158:HT275DSXX:3:1341:10619:11428 chrX 1278197 N chrX 1278549 N DUP 6
A00404:156:HV37TDSXX:4:2677:24876:5087 chrX 1278200 N chrX 1278552 N DUP 5
A00404:156:HV37TDSXX:1:2227:26160:12195 chrX 1278255 N chrX 1278960 N DEL 2
A00404:155:HV27LDSXX:3:1402:9679:2534 chrX 1278344 N chrX 1278698 N DEL 5
A00404:155:HV27LDSXX:1:1324:31277:15608 chrX 1278347 N chrX 1278701 N DEL 9
A00297:158:HT275DSXX:3:2653:24370:34460 chrX 1278019 N chrX 1278376 N DEL 12
A00404:156:HV37TDSXX:1:2424:27887:20885 chrX 1278192 N chrX 1278544 N DUP 5
A00404:156:HV37TDSXX:1:2424:28230:22858 chrX 1278192 N chrX 1278544 N DUP 5
A00297:158:HT275DSXX:3:2219:14588:12696 chrX 1278192 N chrX 1278544 N DUP 5
A00297:158:HT275DSXX:2:1217:1398:14465 chrX 1278192 N chrX 1278544 N DUP 5
A00404:155:HV27LDSXX:2:1368:30743:33818 chrX 1278192 N chrX 1278544 N DUP 5
A00404:155:HV27LDSXX:3:1457:18313:25379 chrX 1278192 N chrX 1278544 N DUP 5
A00297:158:HT275DSXX:4:1134:1099:3020 chrX 1278192 N chrX 1278544 N DUP 5
A00404:155:HV27LDSXX:1:1655:23637:23390 chrX 1278192 N chrX 1278544 N DUP 5
A00404:155:HV27LDSXX:4:2441:30707:8829 chrX 1278192 N chrX 1278544 N DUP 5
A00297:158:HT275DSXX:3:1352:29441:16971 chrX 1278192 N chrX 1278544 N DUP 5
A00404:156:HV37TDSXX:1:1615:10059:23234 chrX 1278192 N chrX 1278544 N DUP 5
A00404:156:HV37TDSXX:1:2615:11487:26115 chrX 1278192 N chrX 1278544 N DUP 5
A00404:156:HV37TDSXX:4:2677:24876:5087 chrX 1278192 N chrX 1278544 N DUP 5
A00404:155:HV27LDSXX:1:2253:15718:35603 chrX 1278192 N chrX 1278544 N DUP 5
A00404:156:HV37TDSXX:2:1524:21630:20917 chrX 1278566 N chrX 1278918 N DEL 10
A00404:155:HV27LDSXX:1:1426:2989:21136 chrX 1278192 N chrX 1278544 N DUP 5
A00404:156:HV37TDSXX:2:1329:11071:6417 chrX 1278192 N chrX 1278544 N DUP 5
A00404:156:HV37TDSXX:2:1329:13141:6621 chrX 1278192 N chrX 1278544 N DUP 5
A00297:158:HT275DSXX:2:2248:11840:17926 chrX 1278192 N chrX 1278544 N DUP 5
A00297:158:HT275DSXX:2:2248:11885:17597 chrX 1278192 N chrX 1278544 N DUP 5
A00297:158:HT275DSXX:2:2170:11885:28745 chrX 1278192 N chrX 1278544 N DUP 6
A00404:155:HV27LDSXX:4:1310:26350:29340 chrX 1278192 N chrX 1278544 N DUP 8
A00297:158:HT275DSXX:1:1570:19199:23531 chrX 1278192 N chrX 1278544 N DUP 10
A00297:158:HT275DSXX:1:1570:20112:21981 chrX 1278192 N chrX 1278544 N DUP 10
A00297:158:HT275DSXX:3:2343:7943:27680 chrX 1278192 N chrX 1278544 N DUP 10
A00404:156:HV37TDSXX:3:2412:29315:28119 chrX 1278192 N chrX 1278544 N DUP 10
A00297:158:HT275DSXX:3:1456:20139:13479 chrX 1278192 N chrX 1278544 N DUP 10
A00297:158:HT275DSXX:3:1456:20148:13463 chrX 1278192 N chrX 1278544 N DUP 10
A00404:155:HV27LDSXX:4:1133:1506:9048 chrX 1278192 N chrX 1278544 N DUP 10
A00404:156:HV37TDSXX:1:1515:14669:32659 chrX 1278192 N chrX 1278544 N DUP 10
A00404:155:HV27LDSXX:2:1133:24578:19789 chrX 1278192 N chrX 1278544 N DUP 10
A00404:156:HV37TDSXX:4:1563:32325:15389 chrX 1278192 N chrX 1278544 N DUP 10
A00297:158:HT275DSXX:3:2671:10031:15295 chrX 1278192 N chrX 1278544 N DUP 10
A00297:158:HT275DSXX:1:2457:21052:28432 chrX 1278192 N chrX 1278544 N DUP 10
A00404:156:HV37TDSXX:1:2654:27688:22357 chrX 1278192 N chrX 1278544 N DUP 10
A00297:158:HT275DSXX:1:1231:2573:18662 chrX 1278193 N chrX 1278545 N DUP 10
A00404:155:HV27LDSXX:3:1567:17508:30749 chrX 1278202 N chrX 1278554 N DUP 5
A00404:155:HV27LDSXX:4:2513:28673:16266 chrX 1278284 N chrX 1278989 N DEL 10
A00297:158:HT275DSXX:2:2135:8567:6715 chrX 1278277 N chrX 1278631 N DEL 5
A00297:158:HT275DSXX:1:1228:11677:21966 chrX 1278609 N chrX 1278959 N DUP 5
A00404:155:HV27LDSXX:3:2278:24126:35697 chrX 1278277 N chrX 1278631 N DEL 5
A00404:156:HV37TDSXX:4:1315:13621:4413 chrX 1278277 N chrX 1278631 N DEL 5
A00404:156:HV37TDSXX:4:1315:13621:4413 chrX 1278277 N chrX 1278631 N DEL 5
A00404:155:HV27LDSXX:1:1205:32732:15937 chrX 1278277 N chrX 1278631 N DEL 5
A00297:158:HT275DSXX:1:1123:22878:1063 chrX 1278277 N chrX 1278631 N DEL 5
A00404:155:HV27LDSXX:3:1402:9679:2534 chrX 1278277 N chrX 1278631 N DEL 5
A00297:158:HT275DSXX:3:1566:10755:34992 chrX 1278277 N chrX 1278631 N DEL 5
A00404:155:HV27LDSXX:4:2444:19931:23672 chrX 1277925 N chrX 1278636 N DEL 5
A00404:155:HV27LDSXX:4:2444:22200:21715 chrX 1277925 N chrX 1278636 N DEL 5
A00297:158:HT275DSXX:3:2343:7943:27680 chrX 1277929 N chrX 1278640 N DEL 5
A00404:155:HV27LDSXX:1:2245:3387:1532 chrX 1277930 N chrX 1278641 N DEL 5
A00297:158:HT275DSXX:1:1131:19786:5165 chrX 1278349 N chrX 1278703 N DEL 5
A00297:158:HT275DSXX:4:1134:1099:3020 chrX 1278129 N chrX 1278833 N DUP 3
A00404:155:HV27LDSXX:1:1324:31277:15608 chrX 1278129 N chrX 1278833 N DUP 7
A00404:155:HV27LDSXX:1:1205:32732:15937 chrX 1277767 N chrX 1278848 N DEL 6
A00404:156:HV37TDSXX:2:1524:21630:20917 chrX 1278210 N chrX 1278915 N DEL 11
A00297:158:HT275DSXX:2:1126:28131:32550 chrX 1278147 N chrX 1278852 N DEL 5
A00297:158:HT275DSXX:1:1231:2573:18662 chrX 1278292 N chrX 1278997 N DEL 10
A00297:158:HT275DSXX:3:1325:27344:10144 chrX 1278296 N chrX 1279001 N DEL 5
A00404:156:HV37TDSXX:1:2569:12057:19648 chr1 21348675 N chr1 21348934 N DEL 1
A00297:158:HT275DSXX:1:1349:28330:5087 chr1 21348674 N chr1 21348930 N DEL 5
A00404:155:HV27LDSXX:2:2176:31665:36198 chr1 21348674 N chr1 21348930 N DEL 5
A00404:155:HV27LDSXX:4:2452:7446:26944 chrX 1895657 N chrX 1896008 N DEL 1
A00297:158:HT275DSXX:2:1365:19162:14387 chrX 1895657 N chrX 1896008 N DEL 3
A00404:155:HV27LDSXX:1:2536:22399:2581 chrX 1895827 N chrX 1896016 N DEL 18
A00297:158:HT275DSXX:1:2647:21802:3051 chr1 241675075 N chr1 241675216 N DUP 13
A00404:155:HV27LDSXX:1:2513:10285:15452 chr1 241675075 N chr1 241675216 N DUP 15
A00404:155:HV27LDSXX:3:2439:20781:26459 chr1 241675075 N chr1 241675216 N DUP 15
A00404:155:HV27LDSXX:2:1643:4725:4100 chr1 241675075 N chr1 241675254 N DUP 1
A00404:156:HV37TDSXX:3:1649:10628:27226 chr1 241675075 N chr1 241675254 N DUP 2
A00404:155:HV27LDSXX:4:1501:24876:36338 chr17 8363923 N chr17 8363980 N DEL 9
A00404:155:HV27LDSXX:3:1609:9055:24533 chr8 139872513 N chr8 139872594 N DEL 5
A00404:156:HV37TDSXX:4:1401:18168:21433 chr8 139872573 N chr8 139872770 N DEL 5
A00404:156:HV37TDSXX:4:1257:5195:2503 chr8 139872426 N chr8 139872543 N DEL 10
A00404:156:HV37TDSXX:2:2362:25861:8985 chr8 139872877 N chr8 139873078 N DEL 43
A00297:158:HT275DSXX:3:1117:6994:6120 chr8 139872626 N chr8 139872877 N DUP 8
A00404:156:HV37TDSXX:1:2660:32190:11741 chr8 139872427 N chr8 139872940 N DEL 1
A00297:158:HT275DSXX:1:2433:27326:5196 chr8 139872926 N chr8 139873053 N DUP 10
A00404:156:HV37TDSXX:3:2559:19253:23062 chr8 139872484 N chr8 139873129 N DEL 15
A00297:158:HT275DSXX:3:2550:6867:19053 chr8 139873090 N chr8 139873201 N DUP 8
A00297:158:HT275DSXX:3:1475:31647:22983 chr8 139872678 N chr8 139873131 N DEL 20
A00297:158:HT275DSXX:3:1475:31846:23234 chr8 139872678 N chr8 139873131 N DEL 20
A00404:156:HV37TDSXX:1:2313:31295:36432 chr8 139872678 N chr8 139873131 N DEL 20
A00404:155:HV27LDSXX:1:2539:7265:11788 chr8 139872485 N chr8 139873130 N DEL 17
A00404:156:HV37TDSXX:4:2101:26368:17472 chr8 139872484 N chr8 139873129 N DEL 20
A00404:155:HV27LDSXX:2:2652:13042:2440 chr8 139872484 N chr8 139873129 N DEL 20
A00404:156:HV37TDSXX:1:2327:21233:28025 chr8 139872810 N chr8 139873131 N DEL 13
A00297:158:HT275DSXX:1:2169:25626:22075 chr14 57333940 N chr14 57334262 N DEL 13
A00404:155:HV27LDSXX:4:2271:2908:28792 chr14 57333996 N chr14 57334316 N DUP 2
A00297:158:HT275DSXX:1:2236:29505:30013 chr14 57333977 N chr14 57334200 N DUP 1
A00297:158:HT275DSXX:1:2236:29677:29371 chr14 57333977 N chr14 57334200 N DUP 1
A00297:158:HT275DSXX:3:1224:32117:18787 chr14 57333977 N chr14 57334200 N DUP 2
A00297:158:HT275DSXX:2:2347:5457:5838 chr14 57333977 N chr14 57334200 N DUP 4
A00404:156:HV37TDSXX:4:1132:13268:22216 chr14 57333977 N chr14 57334200 N DUP 7
A00297:158:HT275DSXX:2:2247:6406:2754 chr14 57333977 N chr14 57334200 N DUP 7
A00297:158:HT275DSXX:2:2465:21838:20870 chr14 57334001 N chr14 57334225 N DEL 7
A00297:158:HT275DSXX:2:2465:21920:20697 chr14 57334001 N chr14 57334225 N DEL 7
A00297:158:HT275DSXX:2:1214:27281:22529 chr14 57334002 N chr14 57334226 N DEL 7
A00404:155:HV27LDSXX:1:2204:22254:35180 chr14 57334001 N chr14 57334225 N DEL 7
A00297:158:HT275DSXX:3:2357:17436:14090 chr11 2367339 N chr11 2367448 N DEL 45
A00297:158:HT275DSXX:3:2357:17436:14090 chr11 2367339 N chr11 2367448 N DEL 39
A00297:158:HT275DSXX:2:2415:3360:33771 chr19 2200856 N chr19 2200929 N DEL 48
A00404:156:HV37TDSXX:3:1316:30572:22247 chr19 2200875 N chr19 2201000 N DUP 5
A00297:158:HT275DSXX:2:1439:5746:6903 chr19 2201081 N chr19 2201154 N DEL 5
A00297:158:HT275DSXX:4:2131:5828:11303 chr19 2201081 N chr19 2201154 N DEL 5
A00404:155:HV27LDSXX:1:2316:2211:11741 chr19 2201081 N chr19 2201154 N DEL 5
A00404:156:HV37TDSXX:1:1617:7012:21746 chr19 2201108 N chr19 2201235 N DEL 16
A00404:156:HV37TDSXX:1:2173:1407:30702 chr19 2201145 N chr19 2201324 N DUP 10
A00404:155:HV27LDSXX:4:2671:7925:10551 chr19 2201135 N chr19 2201278 N DUP 10
A00297:158:HT275DSXX:2:1625:22453:3020 chr19 2201108 N chr19 2201235 N DEL 7
A00404:156:HV37TDSXX:3:2640:11306:14215 chr19 2201216 N chr19 2201269 N DUP 15
A00404:155:HV27LDSXX:1:1134:27688:4413 chr19 2201162 N chr19 2201307 N DEL 10
A00297:158:HT275DSXX:2:2216:15682:10426 chr19 2201120 N chr19 2201229 N DEL 10
A00404:155:HV27LDSXX:1:2149:24189:11318 chr19 2200882 N chr19 2201243 N DEL 5
A00404:156:HV37TDSXX:1:1166:17517:28541 chr19 2200874 N chr19 2201145 N DEL 7
A00297:158:HT275DSXX:2:1101:15980:30389 chr19 2201145 N chr19 2201324 N DUP 10
A00404:156:HV37TDSXX:2:1102:26521:22341 chr19 2201216 N chr19 2201269 N DUP 15
A00404:155:HV27LDSXX:1:2316:2211:11741 chr19 2201145 N chr19 2201324 N DUP 12
A00297:158:HT275DSXX:3:2328:5186:33708 chr19 2201162 N chr19 2201307 N DEL 10
A00297:158:HT275DSXX:3:1532:19976:25598 chr19 2201162 N chr19 2201307 N DEL 10
A00404:156:HV37TDSXX:4:1335:22770:19852 chr19 2201041 N chr19 2201276 N DEL 1
A00297:158:HT275DSXX:1:2206:10294:18975 chr19 2201162 N chr19 2201307 N DEL 10
A00404:156:HV37TDSXX:2:2675:5412:2159 chr19 2200936 N chr19 2201279 N DEL 5
A00404:156:HV37TDSXX:3:2157:22471:21840 chr19 2201253 N chr19 2201362 N DEL 5
A00297:158:HT275DSXX:2:2636:24632:36573 chr19 2201162 N chr19 2201307 N DEL 11
A00404:156:HV37TDSXX:3:2276:14624:26256 chr19 2201260 N chr19 2201315 N DEL 8
A00404:156:HV37TDSXX:1:2128:9372:34851 chr19 2200946 N chr19 2201307 N DEL 8
A00297:158:HT275DSXX:4:1108:3188:24737 chr19 2200958 N chr19 2201319 N DEL 3
A00297:158:HT275DSXX:2:1101:15980:30389 chr19 2200958 N chr19 2201319 N DEL 3
A00404:156:HV37TDSXX:4:1602:28655:35712 chr19 2201180 N chr19 2201343 N DEL 5
A00404:155:HV27LDSXX:2:1560:29767:17722 chr19 2201180 N chr19 2201343 N DEL 5
A00297:158:HT275DSXX:3:2533:10068:23719 chr19 2201000 N chr19 2201379 N DEL 10
A00404:155:HV27LDSXX:4:1658:1470:36918 chr19 2200877 N chr19 2201382 N DEL 5
A00297:158:HT275DSXX:2:2216:15682:10426 chr19 2200881 N chr19 2201404 N DEL 5
A00404:156:HV37TDSXX:3:1423:32823:33223 chr19 2201010 N chr19 2201533 N DEL 5
A00297:158:HT275DSXX:3:1532:19976:25598 chr19 2200854 N chr19 2201557 N DEL 4
A00297:158:HT275DSXX:2:1534:10836:30686 chr19 2200855 N chr19 2201558 N DEL 3
A00404:156:HV37TDSXX:2:2401:10267:15608 chr19 2200855 N chr19 2201558 N DEL 3
A00404:155:HV27LDSXX:1:1620:12581:36057 chr4 3668056 N chr4 3668131 N DEL 5
A00297:158:HT275DSXX:3:1316:6605:17253 chr4 3668079 N chr4 3668133 N DEL 8
A00297:158:HT275DSXX:1:1665:9254:35524 chr4 3668079 N chr4 3668133 N DEL 8
A00404:156:HV37TDSXX:4:2413:14525:2315 chr4 3668088 N chr4 3668165 N DUP 11
A00404:155:HV27LDSXX:1:2245:19506:22874 chr4 3668088 N chr4 3668165 N DUP 10
A00404:156:HV37TDSXX:3:1476:28908:23531 chr4 3668088 N chr4 3668165 N DUP 10
A00404:156:HV37TDSXX:2:2309:29152:21261 chr4 3668088 N chr4 3668165 N DUP 10
A00297:158:HT275DSXX:3:1543:25518:7827 chr7 102334819 N chr7 102334892 N DUP 10
A00404:155:HV27LDSXX:1:1617:11153:34053 chr22 50748385 N chr22 50748561 N DEL 5
A00404:156:HV37TDSXX:4:1538:31259:9345 chr22 50748425 N chr22 50748930 N DEL 5
A00404:156:HV37TDSXX:1:2459:6750:19570 chr22 50748425 N chr22 50748551 N DEL 5
A00297:158:HT275DSXX:1:1515:19479:36010 chr22 50748459 N chr22 50749065 N DEL 2
A00297:158:HT275DSXX:1:2263:10691:15624 chr22 50748434 N chr22 50749040 N DEL 7
A00404:156:HV37TDSXX:4:2175:28818:35869 chr22 50748507 N chr22 50748937 N DEL 5
A00297:158:HT275DSXX:2:2253:26232:8782 chr22 50748507 N chr22 50748937 N DEL 5
A00404:155:HV27LDSXX:4:1116:17571:18051 chr22 50748507 N chr22 50748937 N DEL 5
A00404:156:HV37TDSXX:3:1417:9227:24361 chr22 50748507 N chr22 50748937 N DEL 5
A00404:155:HV27LDSXX:1:2554:5294:24596 chr22 50748507 N chr22 50748937 N DEL 5
A00404:156:HV37TDSXX:1:1350:23357:27853 chr22 50748507 N chr22 50748937 N DEL 5
A00297:158:HT275DSXX:1:1320:18936:25050 chr22 50748507 N chr22 50748937 N DEL 5
A00297:158:HT275DSXX:1:1275:28158:3756 chr22 50748534 N chr22 50748636 N DEL 5
A00404:156:HV37TDSXX:2:2478:26377:34710 chr22 50748534 N chr22 50748636 N DEL 5
A00297:158:HT275DSXX:1:1478:24668:35352 chr22 50748534 N chr22 50748636 N DEL 5
A00404:155:HV27LDSXX:2:1240:25003:10535 chr22 50748534 N chr22 50748636 N DEL 5
A00404:155:HV27LDSXX:2:1240:25021:10535 chr22 50748534 N chr22 50748636 N DEL 5
A00404:155:HV27LDSXX:4:2254:21169:26819 chr22 50748534 N chr22 50748636 N DEL 5
A00297:158:HT275DSXX:1:2166:12653:25974 chr22 50748614 N chr22 50748919 N DEL 7
A00404:155:HV27LDSXX:3:1565:3152:29935 chr22 50748534 N chr22 50748636 N DEL 5
A00404:156:HV37TDSXX:3:2254:24487:24768 chr22 50748534 N chr22 50748636 N DEL 5
A00404:155:HV27LDSXX:2:2556:31204:20932 chr22 50748534 N chr22 50748636 N DEL 5
A00404:155:HV27LDSXX:1:2654:23628:25347 chr22 50748536 N chr22 50748787 N DUP 5
A00404:156:HV37TDSXX:1:1533:32579:3208 chr22 50748536 N chr22 50748787 N DUP 5
A00404:155:HV27LDSXX:2:1305:25898:23672 chr22 50748536 N chr22 50748787 N DUP 5
A00404:156:HV37TDSXX:3:2523:29270:13260 chr22 50748536 N chr22 50748787 N DUP 5
A00297:158:HT275DSXX:3:1655:28718:17347 chr22 50748536 N chr22 50748787 N DUP 5
A00404:155:HV27LDSXX:3:2414:16586:33348 chr22 50748536 N chr22 50748787 N DUP 5
A00404:156:HV37TDSXX:2:2532:6551:17785 chr22 50748536 N chr22 50748787 N DUP 5
A00404:156:HV37TDSXX:4:2114:21947:35900 chr22 50748492 N chr22 50748543 N DEL 5
A00404:155:HV27LDSXX:4:2523:5385:8343 chr22 50748493 N chr22 50748544 N DEL 5
A00404:156:HV37TDSXX:2:2529:32624:17848 chr22 50748495 N chr22 50748546 N DEL 5
A00404:155:HV27LDSXX:3:2374:20311:35227 chr22 50748422 N chr22 50748548 N DEL 3
A00404:155:HV27LDSXX:3:2374:23050:32988 chr22 50748422 N chr22 50748548 N DEL 3
A00404:155:HV27LDSXX:1:2319:6397:27821 chr22 50748590 N chr22 50749018 N DUP 5
A00297:158:HT275DSXX:4:2212:11532:22936 chr22 50748749 N chr22 50749051 N DUP 10
A00404:155:HV27LDSXX:3:2236:11876:1736 chr22 50748812 N chr22 50748940 N DEL 5
A00404:155:HV27LDSXX:4:1415:25843:7576 chr22 50748885 N chr22 50748937 N DEL 12
A00404:155:HV27LDSXX:1:2510:29993:30076 chr22 50748791 N chr22 50748969 N DEL 5
A00297:158:HT275DSXX:2:2625:13856:28213 chr22 50748414 N chr22 50748590 N DEL 5
A00404:156:HV37TDSXX:2:2532:6551:17785 chr22 50748658 N chr22 50748887 N DEL 11
A00404:155:HV27LDSXX:2:2678:23321:1799 chr22 50748658 N chr22 50748887 N DEL 11
A00404:155:HV27LDSXX:4:2356:31313:36902 chr22 50748663 N chr22 50748892 N DEL 11
A00404:156:HV37TDSXX:2:2223:9607:25801 chr22 50748658 N chr22 50748887 N DEL 11
A00404:156:HV37TDSXX:2:2228:27480:32957 chr22 50748887 N chr22 50749011 N DUP 19
A00404:155:HV27LDSXX:3:2501:14009:12352 chr22 50748658 N chr22 50748887 N DEL 11
A00297:158:HT275DSXX:1:2330:8214:29653 chr22 50748809 N chr22 50749088 N DEL 15
A00404:156:HV37TDSXX:2:2327:23285:32205 chr22 50748420 N chr22 50749101 N DEL 2
A00404:156:HV37TDSXX:2:1416:17309:26052 chr22 50748482 N chr22 50749113 N DEL 10
A00297:158:HT275DSXX:3:2418:22191:8140 chr22 50748582 N chr22 50749138 N DEL 5
A00404:155:HV27LDSXX:1:1225:10384:27837 chr22 50748477 N chr22 50749133 N DEL 12
A00297:158:HT275DSXX:4:1628:24551:2456 chr22 50748507 N chr22 50749138 N DEL 5
A00404:155:HV27LDSXX:4:2307:21495:10692 chr2 234544794 N chr2 234544924 N DEL 18
A00404:155:HV27LDSXX:3:1547:19081:22545 chr2 234544833 N chr2 234544889 N DUP 24
A00404:155:HV27LDSXX:3:1547:19434:22185 chr2 234544833 N chr2 234544889 N DUP 24
A00404:156:HV37TDSXX:1:1319:12906:29888 chr2 234544833 N chr2 234544889 N DUP 24
A00297:158:HT275DSXX:1:2245:20889:14528 chr2 234544750 N chr2 234544843 N DEL 14
A00404:156:HV37TDSXX:1:1168:25807:33160 chr2 234544826 N chr2 234544892 N DEL 13
A00404:156:HV37TDSXX:1:1278:2103:34507 chr2 234544831 N chr2 234544897 N DEL 8
A00297:158:HT275DSXX:1:2602:25310:7091 chr2 234544947 N chr2 234545054 N DEL 5
A00404:155:HV27LDSXX:4:2473:29677:36793 chr2 234544950 N chr2 234545057 N DEL 5
A00404:155:HV27LDSXX:3:2663:13648:6277 chr2 234544831 N chr2 234545059 N DEL 3
A00297:158:HT275DSXX:4:1309:31232:27148 chr18 76611836 N chr18 76612058 N DUP 27
A00404:156:HV37TDSXX:2:2111:27471:3850 chr18 76611836 N chr18 76612058 N DUP 25
A00404:156:HV37TDSXX:2:2111:27471:3850 chr18 76611834 N chr18 76611918 N DUP 16
A00404:155:HV27LDSXX:4:1347:1027:8750 chr18 76611926 N chr18 76611990 N DEL 5
A00404:155:HV27LDSXX:4:1126:12418:29982 chr18 76611848 N chr18 76611985 N DUP 20
A00297:158:HT275DSXX:4:1308:32407:5290 chr18 76611840 N chr18 76611932 N DEL 5
A00404:155:HV27LDSXX:3:1248:15519:6637 chr8 4386373 N chr8 4386502 N DEL 5
A00404:156:HV37TDSXX:2:2478:21920:5008 chr8 4386409 N chr8 4386536 N DUP 5
A00404:156:HV37TDSXX:2:2541:23610:25504 chr14 104576865 N chr14 104577062 N DEL 11
A00404:156:HV37TDSXX:4:2241:8531:21151 chr14 104576978 N chr14 104577175 N DEL 38
A00297:158:HT275DSXX:3:1253:15808:7858 chr14 104576875 N chr14 104577121 N DEL 5
A00404:156:HV37TDSXX:4:2268:12581:11099 chr14 104576933 N chr14 104577179 N DEL 30
A00404:155:HV27LDSXX:1:1164:1561:7858 chr14 104576938 N chr14 104577184 N DEL 5
A00297:158:HT275DSXX:1:2101:20374:24095 chr14 104576839 N chr14 104577230 N DEL 5
A00404:156:HV37TDSXX:4:1671:20618:28964 chr5 176252474 N chr5 176252630 N DUP 5
A00404:156:HV37TDSXX:1:1147:19822:10864 chr5 176252474 N chr5 176252746 N DUP 1
A00404:156:HV37TDSXX:2:2121:27624:3458 chr4 16110328 N chr4 16110395 N DUP 13
A00404:155:HV27LDSXX:3:1545:30463:12790 chr4 16110396 N chr4 16110460 N DEL 11
A00404:156:HV37TDSXX:4:1419:11532:2550 chr4 16110324 N chr4 16110417 N DEL 10
A00404:155:HV27LDSXX:2:1539:10872:14779 chr4 16110314 N chr4 16110424 N DEL 5
A00297:158:HT275DSXX:2:1429:25735:15937 chr4 16110375 N chr4 16110460 N DEL 7
A00404:155:HV27LDSXX:3:1542:2040:7811 chr4 16110373 N chr4 16110472 N DEL 12
A00404:156:HV37TDSXX:3:2368:27877:19366 chr4 16110358 N chr4 16110460 N DEL 7
A00297:158:HT275DSXX:3:2118:5466:8453 chr4 16110373 N chr4 16110472 N DEL 12
A00297:158:HT275DSXX:3:2118:5547:5024 chr4 16110373 N chr4 16110472 N DEL 12
A00297:158:HT275DSXX:3:2118:6045:9267 chr4 16110373 N chr4 16110472 N DEL 12
A00404:156:HV37TDSXX:4:2556:15338:29778 chr4 16110358 N chr4 16110460 N DEL 7
A00404:155:HV27LDSXX:2:1357:25183:29105 chr4 16110373 N chr4 16110472 N DEL 12
A00297:158:HT275DSXX:3:1434:4164:29215 chr4 16110355 N chr4 16110471 N DEL 7
A00404:155:HV27LDSXX:2:1623:12301:19977 chr4 16110355 N chr4 16110471 N DEL 7
A00297:158:HT275DSXX:2:1444:16342:15953 chr4 16110356 N chr4 16110472 N DEL 12
A00297:158:HT275DSXX:2:2443:12165:28166 chr4 16110356 N chr4 16110472 N DEL 12
A00404:156:HV37TDSXX:2:2659:2419:4679 chr4 16110321 N chr4 16110460 N DEL 11
A00297:158:HT275DSXX:1:2544:10321:35837 chr13 102234436 N chr13 102234589 N DEL 5
A00404:155:HV27LDSXX:3:1534:23014:3897 chr13 102234436 N chr13 102234589 N DEL 7
A00404:156:HV37TDSXX:1:1157:16984:32878 chr13 102234436 N chr13 102234589 N DEL 7
A00404:156:HV37TDSXX:2:1158:9064:26678 chr13 102234436 N chr13 102234589 N DEL 10
A00404:155:HV27LDSXX:3:2261:6045:36573 chr13 102234436 N chr13 102234589 N DEL 12
A00297:158:HT275DSXX:3:1146:30210:17080 chr13 102234436 N chr13 102234589 N DEL 14
A00297:158:HT275DSXX:4:1668:30951:16799 chr13 102234398 N chr13 102234589 N DEL 10
A00404:156:HV37TDSXX:1:1521:20663:12352 chr17 72900271 N chr17 72900327 N DEL 16
A00404:155:HV27LDSXX:1:1357:16731:10238 chr17 72900291 N chr17 72900367 N DEL 5
A00404:155:HV27LDSXX:4:1244:1958:36041 chr15 50645163 N chr15 50645589 N DEL 10
A00404:155:HV27LDSXX:4:2275:9824:6605 chr15 88941521 N chr15 88941573 N DEL 1
A00297:158:HT275DSXX:3:2230:20112:8923 chr15 88941494 N chr15 88941594 N DUP 2
A00297:158:HT275DSXX:2:1303:2058:20932 chr15 88941434 N chr15 88941612 N DUP 1
A00404:155:HV27LDSXX:2:1475:20057:29778 chr3 153646744 N chr3 153646832 N DEL 10
A00404:156:HV37TDSXX:4:1510:17653:7106 chr3 153646744 N chr3 153646832 N DEL 12
A00404:155:HV27LDSXX:3:2506:13711:21543 chr3 153646744 N chr3 153646832 N DEL 14
A00297:158:HT275DSXX:2:2316:21576:1939 chr3 153646689 N chr3 153646846 N DEL 1
A00297:158:HT275DSXX:4:2115:9326:10222 chr3 153646753 N chr3 153646841 N DEL 6
A00404:156:HV37TDSXX:2:1250:19144:19085 chr3 153646747 N chr3 153646835 N DEL 12
A00404:155:HV27LDSXX:2:2537:30879:13103 chr3 153646753 N chr3 153646841 N DEL 9
A00404:156:HV37TDSXX:1:2335:9390:32409 chr7 128689720 N chr7 128689801 N DEL 5
A00297:158:HT275DSXX:1:2430:10954:4366 chr7 128689737 N chr7 128689858 N DEL 18
A00404:155:HV27LDSXX:1:1152:11767:34929 chr7 128689750 N chr7 128689871 N DEL 2
A00404:155:HV27LDSXX:1:1152:11785:34929 chr7 128689750 N chr7 128689871 N DEL 2
A00404:155:HV27LDSXX:1:1152:12283:35196 chr7 128689750 N chr7 128689871 N DEL 2
A00297:158:HT275DSXX:1:2574:13422:11584 chr19 11488775 N chr19 11489078 N DEL 12
A00297:158:HT275DSXX:2:1601:24523:7639 chr19 11488788 N chr19 11489391 N DEL 22
A00404:156:HV37TDSXX:2:1541:8585:25723 chr9 126899253 N chr9 126899486 N DEL 1
A00297:158:HT275DSXX:1:2313:21097:2456 chr9 126899274 N chr9 126899504 N DUP 3
A00297:158:HT275DSXX:3:2466:14751:34741 chr15 35081691 N chr15 35082561 N DEL 10
A00297:158:HT275DSXX:3:2466:14751:34741 chr15 35081681 N chr15 35081951 N DEL 44
A00404:156:HV37TDSXX:4:1149:12427:33505 chr15 35081708 N chr15 35081783 N DUP 26
A00297:158:HT275DSXX:2:2371:23999:34601 chr15 35081877 N chr15 35082331 N DEL 5
A00404:156:HV37TDSXX:1:2268:9742:13510 chr15 35081960 N chr15 35082561 N DEL 5
A00297:158:HT275DSXX:2:2127:5746:28510 chr15 35081974 N chr15 35082648 N DEL 5
A00297:158:HT275DSXX:4:2211:27127:17910 chr15 35081974 N chr15 35082648 N DEL 5
A00404:155:HV27LDSXX:4:1524:7193:15765 chr15 35081974 N chr15 35082648 N DEL 5
A00404:155:HV27LDSXX:4:1524:7238:15843 chr15 35081974 N chr15 35082648 N DEL 5
A00404:155:HV27LDSXX:3:2421:26549:33974 chr15 35081987 N chr15 35082586 N DUP 5
A00404:156:HV37TDSXX:3:2168:15167:14732 chr15 35081987 N chr15 35082586 N DUP 5
A00404:155:HV27LDSXX:4:2258:12391:27868 chr15 35081987 N chr15 35082586 N DUP 5
A00297:158:HT275DSXX:3:1404:29405:4194 chr15 35082197 N chr15 35082501 N DEL 2
A00297:158:HT275DSXX:4:2211:27127:17910 chr15 35082088 N chr15 35082200 N DUP 5
A00404:155:HV27LDSXX:3:2119:24487:32283 chr15 35082268 N chr15 35082425 N DEL 3
A00404:156:HV37TDSXX:1:2275:28772:20917 chr15 35081718 N chr15 35082283 N DUP 7
A00404:155:HV27LDSXX:2:1436:26386:36918 chr15 35082215 N chr15 35082517 N DUP 5
A00404:155:HV27LDSXX:2:2351:25346:22968 chr15 35082215 N chr15 35082517 N DUP 5
A00404:155:HV27LDSXX:3:2370:20573:21652 chr15 35082215 N chr15 35082517 N DUP 5
A00404:156:HV37TDSXX:1:2211:8621:2174 chr15 35082117 N chr15 35082231 N DEL 4
A00297:158:HT275DSXX:4:2303:9001:2957 chr15 35081853 N chr15 35082304 N DEL 5
A00404:155:HV27LDSXX:2:1309:27190:33959 chr15 35082411 N chr15 35082706 N DEL 5
A00297:158:HT275DSXX:1:2459:29179:35023 chr15 35082411 N chr15 35082706 N DEL 5
A00297:158:HT275DSXX:1:1412:24424:28573 chr15 35081960 N chr15 35082337 N DEL 5
A00297:158:HT275DSXX:4:2549:19099:19570 chr15 35082572 N chr15 35082720 N DEL 11
A00404:155:HV27LDSXX:1:1265:8648:23234 chr15 35081989 N chr15 35082482 N DEL 5
A00404:156:HV37TDSXX:2:2566:30734:24032 chr15 35082615 N chr15 35083030 N DEL 7
A00297:158:HT275DSXX:4:1608:6614:14356 chr15 35081723 N chr15 35082853 N DEL 6
A00404:156:HV37TDSXX:2:2256:5213:1501 chr15 35082800 N chr15 35082914 N DEL 45
A00297:158:HT275DSXX:1:2416:14778:4726 chr15 35082333 N chr15 35082934 N DEL 5
A00297:158:HT275DSXX:3:1406:1678:5400 chr15 35082770 N chr15 35083040 N DEL 20
A00404:156:HV37TDSXX:2:2566:30734:24032 chr15 35081903 N chr15 35083034 N DEL 2
A00404:156:HV37TDSXX:1:2159:25147:20776 chr19 8682864 N chr19 8682945 N DEL 4
A00297:158:HT275DSXX:3:2632:31557:23766 chr9 41104741 N chr9 41104822 N DEL 11
A00404:156:HV37TDSXX:2:2274:3387:34475 chr9 41104872 N chr9 41104953 N DEL 5
A00297:158:HT275DSXX:1:1510:28257:11976 chr9 41104785 N chr9 41104864 N DUP 10
A00297:158:HT275DSXX:4:1143:9887:29387 chr9 41104904 N chr9 41104983 N DUP 8
A00404:155:HV27LDSXX:1:2547:16803:34945 chr9 41104903 N chr9 41104982 N DUP 25
A00404:156:HV37TDSXX:2:2639:1226:16673 chr9 41104893 N chr9 41104972 N DUP 5
A00404:156:HV37TDSXX:4:2572:23972:32424 chr9 41104903 N chr9 41104982 N DUP 19
A00404:156:HV37TDSXX:3:2117:13259:8484 chr9 41104932 N chr9 41105012 N DEL 12
A00404:156:HV37TDSXX:1:1274:20681:29700 chr9 41104764 N chr9 41105004 N DEL 1
A00297:158:HT275DSXX:4:1672:26033:32706 chr9 41104932 N chr9 41105012 N DEL 10
A00404:156:HV37TDSXX:1:2654:17038:36667 chr9 41104934 N chr9 41105014 N DEL 10
A00404:155:HV27LDSXX:1:2316:15917:9674 chr9 41104937 N chr9 41105017 N DEL 8
A00404:156:HV37TDSXX:1:2620:23330:24987 chr19 13554293 N chr19 13554458 N DEL 5
A00297:158:HT275DSXX:2:2563:32371:32816 chr9 137429932 N chr9 137430307 N DEL 12
A00297:158:HT275DSXX:3:2611:5448:4006 chr9 137430100 N chr9 137430309 N DEL 5
A00404:156:HV37TDSXX:2:2258:8558:19695 chr9 137429936 N chr9 137430311 N DEL 5
A00297:158:HT275DSXX:2:2563:32371:32816 chr9 137429944 N chr9 137430319 N DEL 3
A00404:156:HV37TDSXX:4:1373:6696:5509 chr6 131591019 N chr6 131591381 N DEL 24
A00297:158:HT275DSXX:1:2630:5728:1611 chr5 177979518 N chr5 177979635 N DUP 9
A00404:156:HV37TDSXX:2:1216:26539:26349 chr5 177979573 N chr5 177979642 N DEL 7
A00404:156:HV37TDSXX:2:1649:17481:7341 chr5 177979670 N chr5 177979729 N DUP 26
A00297:158:HT275DSXX:2:2544:14687:24267 chr5 177979636 N chr5 177979709 N DUP 12
A00404:155:HV27LDSXX:2:2118:3179:12947 chr5 177979636 N chr5 177979709 N DUP 12
A00404:155:HV27LDSXX:2:2118:3314:12618 chr5 177979636 N chr5 177979709 N DUP 12
A00404:155:HV27LDSXX:2:2118:4444:10911 chr5 177979636 N chr5 177979709 N DUP 12
A00297:158:HT275DSXX:3:1260:10321:35775 chr5 177979519 N chr5 177979636 N DEL 16
A00297:158:HT275DSXX:2:2148:30309:25175 chr5 177979521 N chr5 177979638 N DEL 13
A00297:158:HT275DSXX:4:2354:30734:26600 chr5 177979525 N chr5 177979642 N DEL 9
A00404:155:HV27LDSXX:4:2371:12328:25723 chr5 177979528 N chr5 177979643 N DEL 8
A00404:155:HV27LDSXX:3:2375:29677:10520 chr9 134712159 N chr9 134712339 N DUP 3
A00297:158:HT275DSXX:1:1371:29640:13056 chr14 67193154 N chr14 67193223 N DEL 5
A00297:158:HT275DSXX:1:2151:28158:19946 chr6 69121747 N chr6 69122095 N DEL 5
A00404:156:HV37TDSXX:1:2448:5547:36025 chr6 69121835 N chr6 69121913 N DUP 3
A00404:156:HV37TDSXX:1:2152:19849:10598 chr6 69121843 N chr6 69121922 N DUP 5
A00404:155:HV27LDSXX:3:2539:29677:35509 chr6 69121843 N chr6 69121922 N DUP 5
A00297:158:HT275DSXX:1:1258:26341:18145 chr6 69121843 N chr6 69121922 N DUP 5
A00404:155:HV27LDSXX:3:1123:4119:10473 chr6 69121843 N chr6 69121922 N DUP 5
A00297:158:HT275DSXX:4:1213:9968:33442 chr6 69121843 N chr6 69121922 N DUP 5
A00297:158:HT275DSXX:4:1607:16504:36370 chr6 69121844 N chr6 69121923 N DUP 5
A00404:156:HV37TDSXX:4:1608:10285:12320 chr6 69121843 N chr6 69121922 N DUP 5
A00404:155:HV27LDSXX:2:1307:20003:35947 chr6 69121843 N chr6 69121922 N DUP 5
A00404:155:HV27LDSXX:2:1307:20681:36151 chr6 69121843 N chr6 69121922 N DUP 5
A00404:155:HV27LDSXX:2:2307:15582:35869 chr6 69121843 N chr6 69121922 N DUP 5
A00404:155:HV27LDSXX:1:2264:11017:26647 chr6 69121843 N chr6 69121922 N DUP 5
A00404:155:HV27LDSXX:1:2515:14163:31751 chr6 69122026 N chr6 69122140 N DEL 5
A00404:155:HV27LDSXX:2:1212:26241:14904 chr6 69122026 N chr6 69122140 N DEL 5
A00404:156:HV37TDSXX:4:2371:13819:3129 chr6 69121860 N chr6 69121941 N DEL 1
A00404:155:HV27LDSXX:4:1552:5602:20525 chr6 69122042 N chr6 69122154 N DUP 1
A00404:155:HV27LDSXX:4:2662:22263:4570 chr6 69122015 N chr6 69122167 N DUP 5
A00297:158:HT275DSXX:2:2172:23746:32127 chr11 67996205 N chr11 67996287 N DEL 5
A00297:158:HT275DSXX:4:1276:4860:14387 chr16 80926717 N chr16 80926768 N DUP 10
A00297:158:HT275DSXX:4:1432:14570:30170 chr8 110728468 N chr8 110728534 N DEL 10
A00404:156:HV37TDSXX:3:2267:25030:34444 chr8 110728468 N chr8 110728534 N DEL 10
A00404:156:HV37TDSXX:2:1277:31467:7607 chr8 110728466 N chr8 110728537 N DEL 10
A00297:158:HT275DSXX:4:2350:17273:19977 chrY 26668533 N chrY 26668681 N DUP 5
A00297:158:HT275DSXX:1:1605:20130:36260 chrY 26668586 N chrY 26668697 N DEL 10
A00404:155:HV27LDSXX:2:2347:24198:10300 chrY 26668588 N chrY 26668704 N DEL 5
A00404:156:HV37TDSXX:2:1369:13250:3490 chrY 26668584 N chrY 26668705 N DEL 1
A00404:156:HV37TDSXX:2:2653:7871:4163 chr10 3251930 N chr10 3252019 N DEL 8
A00297:158:HT275DSXX:2:1648:26729:10614 chr10 3251953 N chr10 3252350 N DEL 15
A00404:155:HV27LDSXX:1:1507:11514:19648 chr10 3252108 N chr10 3252329 N DEL 6
A00404:156:HV37TDSXX:1:1127:11758:13119 chr10 3252193 N chr10 3252326 N DEL 10
A00297:158:HT275DSXX:2:1569:19144:21652 chr10 3252216 N chr10 3252524 N DEL 5
A00404:156:HV37TDSXX:2:2344:24017:30342 chr10 3252086 N chr10 3252305 N DUP 1
A00404:155:HV27LDSXX:2:1548:31394:11177 chr10 3251878 N chr10 3252187 N DEL 12
A00404:156:HV37TDSXX:1:1543:26630:33113 chr10 3251937 N chr10 3252246 N DEL 5
A00404:155:HV27LDSXX:4:2478:13675:26428 chr10 3252377 N chr10 3252859 N DEL 5
A00404:155:HV27LDSXX:1:1507:11514:19648 chr10 3252108 N chr10 3252329 N DEL 14
A00404:156:HV37TDSXX:2:2439:19976:28510 chr10 3252124 N chr10 3252430 N DUP 5
A00404:155:HV27LDSXX:1:1538:28067:20228 chr10 3252240 N chr10 3252810 N DEL 18
A00297:158:HT275DSXX:4:2132:31665:10895 chr8 139830348 N chr8 139830404 N DUP 4
A00404:155:HV27LDSXX:3:1673:24297:3552 chr8 139830348 N chr8 139830404 N DUP 9
A00404:155:HV27LDSXX:4:1178:21739:7357 chr8 139830348 N chr8 139830404 N DUP 9
A00404:155:HV27LDSXX:4:2178:16315:7420 chr8 139830348 N chr8 139830404 N DUP 9
A00297:158:HT275DSXX:2:1110:11243:1955 chr8 139830348 N chr8 139830404 N DUP 9
A00404:156:HV37TDSXX:4:1207:23122:1047 chr8 139830348 N chr8 139830404 N DUP 9
A00297:158:HT275DSXX:1:2541:10547:17848 chr8 139830387 N chr8 139830443 N DEL 9
A00404:156:HV37TDSXX:1:1569:22218:6840 chr8 139830387 N chr8 139830443 N DEL 9
A00404:155:HV27LDSXX:4:1610:1913:15483 chr8 139830387 N chr8 139830443 N DEL 9
A00297:158:HT275DSXX:1:1462:21694:20901 chr8 139830387 N chr8 139830443 N DEL 9
A00404:156:HV37TDSXX:2:1135:2437:19586 chrX 71645169 N chrX 71645256 N DUP 5
A00404:155:HV27LDSXX:3:2439:10529:30780 chr18 71568880 N chr18 71568935 N DUP 17
A00404:156:HV37TDSXX:2:1464:8314:29982 chr18 71568880 N chr18 71568935 N DUP 16
A00297:158:HT275DSXX:1:2674:29875:17816 chr18 71568892 N chr18 71568969 N DEL 2
A00297:158:HT275DSXX:4:2203:22471:37027 chr18 71568893 N chr18 71568970 N DEL 1
A00404:156:HV37TDSXX:4:2220:6741:33426 chr1 91168742 N chr1 91168797 N DUP 28
A00297:158:HT275DSXX:2:1409:30011:28573 chr1 91168801 N chr1 91168854 N DEL 13
A00404:156:HV37TDSXX:1:2560:30020:32690 chr1 91168801 N chr1 91168854 N DEL 13
A00404:156:HV37TDSXX:2:1534:8278:10160 chr1 91168801 N chr1 91168854 N DEL 13
A00404:156:HV37TDSXX:2:2243:30318:20369 chr1 91168880 N chr1 91168931 N DUP 6
A00404:156:HV37TDSXX:4:2248:11812:25582 chr1 91168880 N chr1 91168931 N DUP 7
A00404:156:HV37TDSXX:4:1505:32353:24267 chr1 91168773 N chr1 91168854 N DEL 13
A00297:158:HT275DSXX:1:2426:29035:33520 chr1 91168800 N chr1 91168889 N DEL 2
A00404:156:HV37TDSXX:4:2302:29595:5901 chr1 91168951 N chr1 91169132 N DEL 4
A00404:155:HV27LDSXX:3:2330:17155:9283 chr1 91169193 N chr1 91169274 N DUP 7
A00404:156:HV37TDSXX:2:2656:18367:27853 chr1 91169193 N chr1 91169274 N DUP 7
A00404:155:HV27LDSXX:3:1340:17852:29653 chr1 91169193 N chr1 91169274 N DUP 7
A00297:158:HT275DSXX:1:1207:10565:34757 chr1 91169193 N chr1 91169274 N DUP 7
A00297:158:HT275DSXX:4:2321:30237:10895 chr1 91169193 N chr1 91169274 N DUP 7
A00404:155:HV27LDSXX:4:1267:28067:26741 chr1 91169193 N chr1 91169274 N DUP 7
A00297:158:HT275DSXX:1:2372:5972:9956 chr1 91169193 N chr1 91169274 N DUP 7
A00404:156:HV37TDSXX:1:1255:16034:2863 chr1 91169163 N chr1 91169288 N DUP 3
A00404:156:HV37TDSXX:2:1621:13078:8860 chr1 91169193 N chr1 91169274 N DUP 7
A00404:155:HV27LDSXX:2:2108:29505:5744 chr9 81697902 N chr9 81698194 N DEL 4
A00297:158:HT275DSXX:2:1474:20446:12508 chr10 92556597 N chr10 92556731 N DUP 1
A00404:156:HV37TDSXX:4:2459:3929:9330 chr8 27865725 N chr8 27865904 N DEL 5
A00404:155:HV27LDSXX:2:1650:30056:18756 chr8 27865726 N chr8 27865905 N DUP 1
A00297:158:HT275DSXX:4:1631:5403:30733 chrX 779171 N chrX 779238 N DEL 3
A00404:156:HV37TDSXX:1:2159:21169:26412 chrX 779179 N chrX 779609 N DEL 10
A00404:156:HV37TDSXX:3:1415:22390:29434 chrX 779171 N chrX 779400 N DEL 13
A00404:155:HV27LDSXX:4:1329:7148:9455 chrX 779174 N chrX 779399 N DEL 37
A00404:155:HV27LDSXX:4:2329:5755:16939 chrX 779174 N chrX 779399 N DEL 37
A00404:155:HV27LDSXX:4:1329:7157:9471 chrX 779178 N chrX 779399 N DEL 41
A00404:155:HV27LDSXX:4:1216:27724:31125 chrX 779253 N chrX 779511 N DEL 5
A00404:155:HV27LDSXX:3:2441:21793:25113 chrX 779204 N chrX 779621 N DUP 11
A00404:155:HV27LDSXX:2:1110:12292:24158 chrX 779202 N chrX 779619 N DUP 13
A00404:155:HV27LDSXX:1:1603:29333:30749 chrX 779213 N chrX 779315 N DUP 4
A00404:155:HV27LDSXX:2:1641:32796:35086 chrX 779213 N chrX 779315 N DUP 4
A00297:158:HT275DSXX:3:1560:31575:8171 chrX 779187 N chrX 779246 N DEL 7
A00404:156:HV37TDSXX:3:1538:7780:29183 chrX 779275 N chrX 779436 N DUP 10
A00404:156:HV37TDSXX:3:1337:28736:15843 chrX 779275 N chrX 779436 N DUP 10
A00404:156:HV37TDSXX:4:2274:5999:26631 chrX 779202 N chrX 779306 N DEL 13
A00297:158:HT275DSXX:1:1656:15673:17989 chrX 779419 N chrX 779675 N DUP 30
A00404:155:HV27LDSXX:2:1372:9489:10128 chrX 779236 N chrX 779551 N DUP 14
A00404:156:HV37TDSXX:2:2655:11279:5776 chrX 779474 N chrX 779526 N DEL 5
A00404:155:HV27LDSXX:2:1227:2654:15107 chrX 779216 N chrX 779529 N DEL 10
A00404:156:HV37TDSXX:4:1468:14326:25614 chrX 779555 N chrX 779625 N DUP 2
A00297:158:HT275DSXX:1:1423:23312:27023 chrX 779569 N chrX 779639 N DUP 5
A00404:155:HV27LDSXX:2:1429:26142:4742 chrX 779183 N chrX 779682 N DUP 9
A00297:158:HT275DSXX:2:2312:11659:6621 chr11 28430357 N chr11 28430632 N DEL 3
A00404:156:HV37TDSXX:2:2452:8965:6151 chr11 28430349 N chr11 28430624 N DEL 11
A00404:156:HV37TDSXX:2:2452:8965:6151 chr11 28430349 N chr11 28430624 N DEL 28
A00404:155:HV27LDSXX:3:2568:9028:14309 chr11 28430361 N chr11 28430459 N DUP 5
A00404:155:HV27LDSXX:1:1412:23384:19163 chr11 28430459 N chr11 28430684 N DEL 5
A00404:156:HV37TDSXX:3:2102:3115:7983 chr11 28430408 N chr11 28430505 N DUP 7
A00297:158:HT275DSXX:1:2472:29866:27821 chr11 28430508 N chr11 28430684 N DEL 7
A00404:155:HV27LDSXX:4:2206:23619:5666 chr11 28430422 N chr11 28430520 N DEL 7
A00404:155:HV27LDSXX:3:1136:24768:3615 chr11 28430423 N chr11 28430521 N DEL 7
A00404:156:HV37TDSXX:3:1304:29053:14074 chr11 28430530 N chr11 28430705 N DUP 1
A00404:155:HV27LDSXX:1:2355:26802:10144 chr11 28430425 N chr11 28430649 N DUP 2
A00404:155:HV27LDSXX:2:1549:12048:24424 chr9 137669472 N chr9 137669586 N DEL 8
A00404:155:HV27LDSXX:3:1469:1063:27508 chr9 137669474 N chr9 137669699 N DEL 14
A00404:156:HV37TDSXX:2:1202:1154:10097 chr9 137669470 N chr9 137669544 N DEL 12
A00404:156:HV37TDSXX:3:1257:15682:24017 chr9 137669470 N chr9 137669544 N DEL 13
A00404:156:HV37TDSXX:4:1538:5159:9643 chr9 137669470 N chr9 137669544 N DEL 20
A00404:156:HV37TDSXX:2:2309:5773:34695 chr9 137669470 N chr9 137669544 N DEL 20
A00404:155:HV27LDSXX:4:2101:6063:18662 chr9 137669470 N chr9 137669544 N DEL 23
A00404:155:HV27LDSXX:4:2244:30544:25394 chr9 137669529 N chr9 137669605 N DUP 6
A00404:155:HV27LDSXX:2:1405:30581:19914 chr9 137669534 N chr9 137669724 N DUP 7
A00404:155:HV27LDSXX:2:2141:21043:22529 chr9 137669496 N chr9 137669645 N DUP 11
A00404:156:HV37TDSXX:4:1457:22806:33880 chr9 137669572 N chr9 137669722 N DUP 14
A00404:155:HV27LDSXX:4:2332:1434:18881 chr9 137669527 N chr9 137669714 N DUP 19
A00404:155:HV27LDSXX:4:2332:2112:19742 chr9 137669527 N chr9 137669714 N DUP 19
A00404:155:HV27LDSXX:4:2332:3766:18599 chr9 137669527 N chr9 137669714 N DUP 19
A00297:158:HT275DSXX:2:2530:10936:18396 chr9 137669563 N chr9 137669641 N DEL 5
A00404:155:HV27LDSXX:4:2123:32452:24314 chr9 137669546 N chr9 137669661 N DEL 2
A00404:155:HV27LDSXX:3:2654:2944:29794 chr18 77400064 N chr18 77400144 N DEL 5
A00404:155:HV27LDSXX:1:1222:11369:28134 chr18 77400083 N chr18 77400161 N DUP 5
A00404:156:HV37TDSXX:4:1354:21603:22153 chr16 32843101 N chr16 32843313 N DEL 10
A00297:158:HT275DSXX:3:1209:15139:6793 chr16 32843101 N chr16 32843313 N DEL 10
A00404:155:HV27LDSXX:4:1601:25545:8688 chr16 32843043 N chr16 32843122 N DEL 1
A00404:155:HV27LDSXX:4:1601:27317:9815 chr16 32843043 N chr16 32843122 N DEL 1
A00404:155:HV27LDSXX:4:2667:5855:25911 chr16 32843041 N chr16 32843120 N DEL 3
A00404:155:HV27LDSXX:2:1371:8070:26991 chr16 32843042 N chr16 32843121 N DEL 2
A00404:155:HV27LDSXX:2:1371:8088:26929 chr16 32843042 N chr16 32843121 N DEL 2
A00297:158:HT275DSXX:4:1506:20139:25848 chr5 26793752 N chr5 26793803 N DEL 5
A00404:156:HV37TDSXX:4:1614:17264:30107 chr22 47212949 N chr22 47213027 N DUP 5
A00404:155:HV27LDSXX:4:2372:32334:13651 chr22 47213024 N chr22 47213076 N DUP 5
A00297:158:HT275DSXX:2:1140:8748:20369 chr22 47212959 N chr22 47213072 N DEL 5
A00297:158:HT275DSXX:2:1140:9164:7247 chr22 47213173 N chr22 47213414 N DEL 5
A00404:156:HV37TDSXX:3:1376:27814:3004 chr22 47212961 N chr22 47213074 N DEL 5
A00404:156:HV37TDSXX:1:1510:21350:14638 chr22 47213180 N chr22 47213553 N DEL 5
A00404:155:HV27LDSXX:4:1432:16170:2096 chr22 47213035 N chr22 47213261 N DUP 5
A00404:155:HV27LDSXX:3:1163:10926:12085 chr22 47213021 N chr22 47213201 N DEL 5
A00297:158:HT275DSXX:4:2504:14244:5243 chr22 47213024 N chr22 47213204 N DEL 5
A00404:155:HV27LDSXX:3:1341:15338:33536 chr22 47213067 N chr22 47213227 N DEL 3
A00297:158:HT275DSXX:1:1470:20600:24737 chr22 47213139 N chr22 47213382 N DUP 2
A00297:158:HT275DSXX:1:1470:21603:16579 chr22 47213139 N chr22 47213382 N DUP 2
A00404:155:HV27LDSXX:1:2357:15456:29105 chr22 47212991 N chr22 47213398 N DEL 8
A00404:155:HV27LDSXX:2:1123:32063:9768 chr22 47212931 N chr22 47213505 N DUP 18
A00404:155:HV27LDSXX:4:1350:7265:1329 chr22 47213200 N chr22 47213461 N DEL 24
A00297:158:HT275DSXX:1:1348:25427:17190 chrX 68592929 N chrX 68592986 N DUP 27
A00297:158:HT275DSXX:4:1502:22354:17785 chrX 68592902 N chrX 68592956 N DUP 19
A00404:155:HV27LDSXX:3:1457:25880:18537 chrX 68592932 N chrX 68593019 N DUP 11
A00297:158:HT275DSXX:4:2626:31114:27571 chr7 158126293 N chr7 158126816 N DEL 9
A00297:158:HT275DSXX:1:2407:4562:18850 chr7 158126348 N chr7 158126652 N DEL 5
A00404:155:HV27LDSXX:3:2216:15257:2926 chr7 158126235 N chr7 158126801 N DEL 14
A00297:158:HT275DSXX:4:2614:15203:25504 chr7 158126775 N chr7 158126863 N DEL 5
A00404:156:HV37TDSXX:4:2429:3097:33191 chr7 158126713 N chr7 158126801 N DEL 5
A00297:158:HT275DSXX:2:2420:10140:35931 chr7 158126514 N chr7 158126864 N DEL 7
A00404:156:HV37TDSXX:4:1407:3134:22952 chr7 158126191 N chr7 158126801 N DEL 5
A00404:155:HV27LDSXX:3:2216:15257:2926 chr7 158126196 N chr7 158126806 N DEL 5
A00404:155:HV27LDSXX:1:1320:28546:18114 chr21 28314953 N chr21 28315065 N DEL 2
A00404:156:HV37TDSXX:4:1569:3775:23782 chr21 28314953 N chr21 28315065 N DEL 2
A00297:158:HT275DSXX:3:1107:30617:19507 chr12 28863698 N chr12 28863865 N DEL 3
A00297:158:HT275DSXX:3:1107:31394:19601 chr12 28863698 N chr12 28863865 N DEL 3
A00297:158:HT275DSXX:2:2642:31665:30749 chr5 11240275 N chr5 11240384 N DUP 12
A00297:158:HT275DSXX:2:2642:31665:30749 chr5 11240275 N chr5 11240384 N DUP 13
A00297:158:HT275DSXX:2:2321:27317:36276 chr5 11240401 N chr5 11240878 N DUP 4
A00297:158:HT275DSXX:3:2233:25111:4648 chr5 11240691 N chr5 11240844 N DEL 9
A00404:156:HV37TDSXX:2:2546:27959:25144 chr5 11240288 N chr5 11240621 N DEL 5
A00404:155:HV27LDSXX:4:1318:24388:2268 chr5 11240739 N chr5 11241130 N DEL 11
A00404:155:HV27LDSXX:4:1318:24388:2268 chr5 11240739 N chr5 11241130 N DEL 12
A00297:158:HT275DSXX:4:2367:21133:18364 chr5 11240294 N chr5 11240701 N DEL 9
A00404:155:HV27LDSXX:4:1414:32425:34538 chr5 11240436 N chr5 11240710 N DEL 4
A00404:155:HV27LDSXX:3:2349:20283:12508 chr5 11240917 N chr5 11241003 N DUP 5
A00297:158:HT275DSXX:1:1576:14895:7091 chr5 11240301 N chr5 11241154 N DEL 5
A00297:158:HT275DSXX:2:2567:27896:27884 chr5 11240811 N chr5 11241230 N DEL 1
A00404:156:HV37TDSXX:4:1552:2166:4053 chr12 124358068 N chr12 124358249 N DUP 5
A00404:156:HV37TDSXX:1:2267:3387:10520 chr16 89619614 N chr16 89619672 N DUP 11
A00404:155:HV27LDSXX:1:1365:3007:3505 chr16 89619628 N chr16 89619687 N DUP 5
A00404:155:HV27LDSXX:4:2631:22191:36417 chr16 89619625 N chr16 89619723 N DUP 1
A00404:156:HV37TDSXX:4:1664:7066:34804 chr16 89619850 N chr16 89619914 N DEL 8
A00404:155:HV27LDSXX:4:1556:13612:14325 chr11 76934811 N chr11 76934863 N DUP 12
A00404:155:HV27LDSXX:1:2611:3748:7012 chr11 76934811 N chr11 76934863 N DUP 16
A00404:155:HV27LDSXX:3:1135:19569:30091 chr11 76934825 N chr11 76934877 N DUP 1
A00297:158:HT275DSXX:4:1431:8929:15264 chr11 76934824 N chr11 76934876 N DUP 2
A00404:156:HV37TDSXX:2:2656:17390:4022 chr21 43313197 N chr21 43313290 N DUP 15
A00404:156:HV37TDSXX:2:2113:8983:11162 chrX 147489113 N chrX 147489274 N DEL 7
A00404:155:HV27LDSXX:3:2417:28791:27712 chrX 147489113 N chrX 147489274 N DEL 7
A00404:155:HV27LDSXX:4:2657:1561:37012 chr18 61970198 N chr18 61971204 N DEL 12
A00297:158:HT275DSXX:3:2367:3766:19225 chr18 61970198 N chr18 61971204 N DEL 12
A00404:155:HV27LDSXX:4:2417:26567:23766 chr18 61970198 N chr18 61971204 N DEL 12
A00297:158:HT275DSXX:3:2123:30906:26271 chr18 61970198 N chr18 61971204 N DEL 12
A00404:155:HV27LDSXX:1:2475:15248:31469 chr18 61971182 N chr18 61971610 N DUP 11
A00297:158:HT275DSXX:3:2473:5195:8547 chr16 64876213 N chr16 64876276 N DUP 2
A00404:156:HV37TDSXX:4:1359:27308:30530 chr16 64876213 N chr16 64876276 N DUP 2
A00297:158:HT275DSXX:1:2444:22119:21198 chr16 64876213 N chr16 64876276 N DUP 5
A00404:155:HV27LDSXX:1:1357:11668:6324 chr16 64876213 N chr16 64876276 N DUP 8
A00297:158:HT275DSXX:4:2172:12246:28401 chr16 64876213 N chr16 64876308 N DUP 21
A00404:156:HV37TDSXX:1:2131:6659:27054 chr16 64876222 N chr16 64876285 N DUP 20
A00404:155:HV27LDSXX:1:2344:6099:30311 chr16 64876213 N chr16 64876276 N DUP 23
A00404:156:HV37TDSXX:4:1406:14488:21010 chr16 64876213 N chr16 64876276 N DUP 27
A00404:155:HV27LDSXX:3:1158:13367:32910 chr16 64876213 N chr16 64876276 N DUP 27
A00404:155:HV27LDSXX:1:2276:14669:33442 chr16 64876206 N chr16 64876303 N DEL 9
A00404:156:HV37TDSXX:1:1313:12120:31000 chr16 64876228 N chr16 64876309 N DEL 3
A00297:158:HT275DSXX:4:1175:29749:33755 chr16 64876211 N chr16 64876308 N DEL 4
A00297:158:HT275DSXX:2:1260:7997:12806 chr3 10642163 N chr3 10642232 N DUP 7
A00404:156:HV37TDSXX:2:2132:10050:3396 chr2 169786290 N chr2 169786416 N DUP 1
A00404:155:HV27LDSXX:1:1666:27145:32440 chr2 169786394 N chr2 169786623 N DEL 3
A00297:158:HT275DSXX:1:1221:1787:11882 chr2 87092042 N chr2 87092141 N DUP 5
A00404:155:HV27LDSXX:2:2343:18430:32565 chr4 186239656 N chr4 186239864 N DUP 5
A00404:155:HV27LDSXX:1:1111:16315:2378 chr1 39111476 N chr1 39111662 N DUP 5
A00404:155:HV27LDSXX:4:1137:32597:33207 chr9 6728468 N chr9 6728778 N DUP 5
A00404:156:HV37TDSXX:1:2273:16278:30624 chr9 6728480 N chr9 6728792 N DEL 5
A00404:155:HV27LDSXX:2:2662:2175:1564 chr19 12312690 N chr19 12312855 N DUP 5
A00404:156:HV37TDSXX:4:2122:23737:28886 chr19 12312839 N chr19 12313144 N DEL 42
A00297:158:HT275DSXX:2:2530:1841:14700 chr19 12313024 N chr19 12313325 N DEL 10
A00404:156:HV37TDSXX:3:1220:6307:18051 chr20 58695164 N chr20 58695370 N DEL 5
A00404:155:HV27LDSXX:4:1506:25400:21245 chr20 58695164 N chr20 58695370 N DEL 7
A00404:156:HV37TDSXX:3:2528:31991:22639 chr20 58695164 N chr20 58695370 N DEL 28
A00404:155:HV27LDSXX:1:1313:8621:14199 chr20 58695179 N chr20 58695295 N DUP 4
A00404:156:HV37TDSXX:3:1471:17418:6825 chr20 58695174 N chr20 58695225 N DUP 9
A00404:155:HV27LDSXX:2:1416:4661:30639 chr20 58695378 N chr20 58695437 N DUP 5
A00404:155:HV27LDSXX:2:1152:4725:8484 chr20 58695394 N chr20 58695455 N DEL 5
A00404:155:HV27LDSXX:4:1502:27516:19899 chr20 58695398 N chr20 58695459 N DEL 5
A00297:158:HT275DSXX:3:1152:10402:7012 chr5 1870800 N chr5 1870913 N DUP 13
A00404:155:HV27LDSXX:4:1565:2663:15186 chr19 57606594 N chr19 57606931 N DEL 10
A00404:156:HV37TDSXX:2:2403:12943:2707 chr19 57606890 N chr19 57606973 N DUP 5
A00404:155:HV27LDSXX:4:1565:2663:15186 chr19 57606594 N chr19 57606931 N DEL 22
A00404:156:HV37TDSXX:2:2266:31620:24345 chr19 57607164 N chr19 57607417 N DEL 5
A00404:156:HV37TDSXX:3:2536:12481:9580 chr19 57606572 N chr19 57607413 N DEL 5
A00297:158:HT275DSXX:3:2678:32696:10864 chr11 42682141 N chr11 42682330 N DEL 11
A00297:158:HT275DSXX:4:1116:25961:27915 chr11 42682143 N chr11 42682330 N DEL 12
A00404:155:HV27LDSXX:2:1658:1570:27727 chr11 42682141 N chr11 42682330 N DEL 31
A00404:156:HV37TDSXX:2:2623:2465:5196 chr11 42682252 N chr11 42682347 N DEL 5
A00297:158:HT275DSXX:1:2656:21169:5024 chr11 42682252 N chr11 42682347 N DEL 5
A00404:155:HV27LDSXX:3:1266:14371:18771 chr11 42682268 N chr11 42682403 N DEL 5
A00404:155:HV27LDSXX:4:1108:8693:30044 chr11 42682268 N chr11 42682407 N DUP 8
A00297:158:HT275DSXX:2:1168:23701:23469 chr11 42682222 N chr11 42682317 N DUP 9
A00404:155:HV27LDSXX:3:1507:3432:14356 chr11 42682214 N chr11 42682401 N DUP 12
A00297:158:HT275DSXX:4:2308:25165:7560 chr11 42682291 N chr11 42682342 N DEL 7
A00404:156:HV37TDSXX:4:2341:15546:8437 chr11 42682222 N chr11 42682451 N DUP 16
A00404:155:HV27LDSXX:4:1134:29957:19617 chr11 42682243 N chr11 42682342 N DEL 7
A00404:156:HV37TDSXX:4:2536:27055:9580 chr11 42682243 N chr11 42682342 N DEL 7
A00404:155:HV27LDSXX:3:2306:6451:33583 chr11 42682246 N chr11 42682345 N DEL 7
A00404:156:HV37TDSXX:1:1143:30300:29637 chr11 42682248 N chr11 42682347 N DEL 7
A00404:155:HV27LDSXX:2:1434:4643:34147 chr11 42682248 N chr11 42682347 N DEL 7
A00404:155:HV27LDSXX:1:1221:9426:4163 chr17 20984965 N chr17 20985190 N DUP 3
A00404:155:HV27LDSXX:1:2364:5547:11224 chr17 20984870 N chr17 20985073 N DUP 5
A00297:158:HT275DSXX:2:2453:5285:19695 chr17 20985062 N chr17 20985368 N DEL 11
A00404:155:HV27LDSXX:1:2660:27561:15405 chr17 20984892 N chr17 20984997 N DEL 4
A00297:158:HT275DSXX:2:2319:30147:33818 chr17 20985128 N chr17 20985307 N DEL 5
A00297:158:HT275DSXX:2:2171:23384:25488 chr17 20985128 N chr17 20985307 N DEL 5
A00404:155:HV27LDSXX:4:1521:12572:7576 chr17 20985128 N chr17 20985307 N DEL 5
A00404:155:HV27LDSXX:1:2641:16993:22686 chr17 20984912 N chr17 20985068 N DEL 5
A00297:158:HT275DSXX:4:1507:14950:29481 chr17 20985239 N chr17 20985596 N DUP 12
A00404:156:HV37TDSXX:4:2354:14199:36104 chr17 20984888 N chr17 20985219 N DEL 7
A00404:155:HV27LDSXX:2:1630:26657:36980 chr17 20985108 N chr17 20985363 N DUP 5
A00297:158:HT275DSXX:1:2263:31810:9298 chr17 20985088 N chr17 20985264 N DEL 3
A00404:156:HV37TDSXX:2:2467:25599:26318 chr17 20985090 N chr17 20985268 N DEL 8
A00404:155:HV27LDSXX:3:2624:30228:24158 chr17 20984892 N chr17 20985270 N DEL 9
A00297:158:HT275DSXX:2:1433:31530:36746 chr17 20985314 N chr17 20985391 N DUP 5
A00297:158:HT275DSXX:1:1658:18249:26334 chr17 20985266 N chr17 20985445 N DUP 7
A00297:158:HT275DSXX:2:1425:29749:15280 chr17 20985266 N chr17 20985445 N DUP 7
A00297:158:HT275DSXX:4:1428:12545:20369 chr17 20985266 N chr17 20985445 N DUP 7
A00404:155:HV27LDSXX:3:2254:25346:8531 chr17 20985113 N chr17 20985370 N DEL 8
A00404:156:HV37TDSXX:1:2241:3577:28228 chr17 20985279 N chr17 20985457 N DUP 4
A00297:158:HT275DSXX:3:1649:21847:17785 chr17 20985266 N chr17 20985446 N DUP 12
A00404:155:HV27LDSXX:1:1506:22444:21668 chr17 20985251 N chr17 20985429 N DUP 5
A00404:155:HV27LDSXX:2:2106:32226:36292 chr17 20985251 N chr17 20985429 N DUP 5
A00297:158:HT275DSXX:1:1610:15718:29622 chr17 20985251 N chr17 20985429 N DUP 5
A00297:158:HT275DSXX:1:2560:17336:4304 chr17 20985262 N chr17 20985393 N DEL 3
A00404:156:HV37TDSXX:2:2347:27896:6903 chr17 20985251 N chr17 20985429 N DUP 5
A00404:156:HV37TDSXX:3:1461:18394:4914 chr17 20985251 N chr17 20985429 N DUP 5
A00297:158:HT275DSXX:1:2560:17336:4304 chr17 20985264 N chr17 20985395 N DEL 1
A00404:156:HV37TDSXX:1:2222:11324:11115 chr17 20985251 N chr17 20985429 N DUP 5
A00404:155:HV27LDSXX:3:1565:11614:20697 chr17 20985251 N chr17 20985429 N DUP 5
A00297:158:HT275DSXX:2:2453:5285:19695 chr17 20985251 N chr17 20985429 N DUP 5
A00404:155:HV27LDSXX:4:1553:19289:29481 chr17 20985251 N chr17 20985429 N DUP 5
A00404:156:HV37TDSXX:1:1462:3893:36292 chr17 20985251 N chr17 20985429 N DUP 5
A00404:156:HV37TDSXX:1:1462:4001:36793 chr17 20985251 N chr17 20985429 N DUP 5
A00297:158:HT275DSXX:3:2414:1696:33301 chr17 20985251 N chr17 20985429 N DUP 5
A00297:158:HT275DSXX:1:2519:2121:17597 chr17 20985252 N chr17 20985430 N DUP 5
A00404:155:HV27LDSXX:3:2464:18719:1438 chr17 20985251 N chr17 20985429 N DUP 5
A00404:155:HV27LDSXX:2:2346:20609:31297 chr17 20984920 N chr17 20985251 N DEL 5
A00297:158:HT275DSXX:4:2112:13684:22060 chr17 20984925 N chr17 20985256 N DEL 5
A00404:155:HV27LDSXX:4:2156:31982:28635 chr17 20985103 N chr17 20985460 N DEL 1
A00297:158:HT275DSXX:2:2162:1488:1908 chr17 20985103 N chr17 20985460 N DEL 1
A00404:155:HV27LDSXX:4:1650:24071:2660 chr17 20985414 N chr17 20985467 N DEL 6
A00404:156:HV37TDSXX:4:2162:7012:9220 chr17 20985129 N chr17 20985487 N DEL 5
A00404:155:HV27LDSXX:2:1147:30427:36996 chr17 20985132 N chr17 20985490 N DEL 5
A00404:155:HV27LDSXX:2:2475:5810:13495 chr17 20985406 N chr17 20985584 N DUP 3
A00404:156:HV37TDSXX:2:1640:12843:1752 chr17 20985406 N chr17 20985584 N DUP 3
A00404:156:HV37TDSXX:3:2235:17219:21198 chr17 20985335 N chr17 20985513 N DUP 3
A00297:158:HT275DSXX:3:2631:7898:6089 chr17 20985043 N chr17 20985624 N DUP 5
A00404:155:HV27LDSXX:4:2651:29017:17268 chr17 20985365 N chr17 20985589 N DUP 13
A00297:158:HT275DSXX:2:1248:2157:15186 chr17 20985543 N chr17 20985640 N DUP 5
A00297:158:HT275DSXX:1:2419:12246:36824 chr17 20985541 N chr17 20985638 N DUP 10
A00297:158:HT275DSXX:1:2419:12472:36777 chr17 20985541 N chr17 20985638 N DUP 10
A00297:158:HT275DSXX:1:2639:3323:34460 chr17 20985543 N chr17 20985640 N DUP 5
A00404:156:HV37TDSXX:1:1261:18665:13620 chr17 20985091 N chr17 20985625 N DEL 5
A00297:158:HT275DSXX:1:1265:16360:31641 chr17 20985091 N chr17 20985625 N DEL 5
A00297:158:HT275DSXX:1:1267:13503:1266 chr17 20985091 N chr17 20985625 N DEL 5
A00404:155:HV27LDSXX:4:1451:17445:8406 chr17 20984891 N chr17 20985629 N DEL 5
A00404:156:HV37TDSXX:2:2633:26187:26772 chr17 20984892 N chr17 20985630 N DEL 5
A00297:158:HT275DSXX:2:1447:30047:11443 chr22 31366466 N chr22 31366809 N DEL 2
A00404:155:HV27LDSXX:2:2153:3992:11193 chr16 84949429 N chr16 84949554 N DUP 12
A00404:156:HV37TDSXX:4:1664:5864:6386 chr16 84949548 N chr16 84949601 N DUP 7
A00404:156:HV37TDSXX:3:2134:9824:15342 chr16 84949548 N chr16 84949601 N DUP 7
A00297:158:HT275DSXX:2:2312:25663:4319 chr10 16147992 N chr10 16148171 N DEL 5
A00297:158:HT275DSXX:2:2165:29894:1438 chr19 4145659 N chr19 4145896 N DUP 7
A00297:158:HT275DSXX:2:1218:12780:21089 chr16 79825391 N chr16 79825464 N DEL 14
A00404:156:HV37TDSXX:2:1636:31539:28213 chr16 79825302 N chr16 79825555 N DEL 5
A00404:156:HV37TDSXX:2:1503:27046:14700 chr13 107680871 N chr13 107680963 N DEL 9
A00404:156:HV37TDSXX:2:1503:28013:14904 chr13 107680871 N chr13 107680963 N DEL 9
A00297:158:HT275DSXX:3:1466:20482:31861 chr13 107680871 N chr13 107680963 N DEL 9
A00404:155:HV27LDSXX:4:2473:22146:8625 chr13 107680871 N chr13 107680963 N DEL 9
A00404:155:HV27LDSXX:4:1410:32063:28432 chr13 107680871 N chr13 107680963 N DEL 9
A00404:155:HV27LDSXX:4:2410:31277:25191 chr13 107680871 N chr13 107680963 N DEL 9
A00404:155:HV27LDSXX:4:2410:31394:24925 chr13 107680871 N chr13 107680963 N DEL 9
A00297:158:HT275DSXX:3:2223:15781:15107 chr13 107680871 N chr13 107680963 N DEL 9
A00404:156:HV37TDSXX:3:1161:4047:14262 chr13 107680871 N chr13 107680963 N DEL 9
A00404:156:HV37TDSXX:1:1277:17363:23077 chr13 107680903 N chr13 107680995 N DUP 8
A00404:156:HV37TDSXX:4:2506:14344:35916 chr13 107680910 N chr13 107681002 N DUP 1
A00404:156:HV37TDSXX:4:2545:10357:10755 chr13 107680906 N chr13 107680998 N DUP 5
A00404:156:HV37TDSXX:4:2545:10673:11083 chr13 107680906 N chr13 107680998 N DUP 5
A00297:158:HT275DSXX:3:2552:23963:13150 chrX 543239 N chrX 543559 N DEL 10
A00297:158:HT275DSXX:1:1434:32588:14090 chrX 543206 N chrX 543526 N DEL 5
A00297:158:HT275DSXX:1:2677:8549:1986 chr1 195848550 N chr1 195848602 N DEL 5
A00404:155:HV27LDSXX:4:1662:10890:11741 chr7 5449426 N chr7 5449621 N DEL 14
A00404:155:HV27LDSXX:4:1662:9905:12790 chr7 5449407 N chr7 5449600 N DEL 18
A00404:156:HV37TDSXX:4:2560:2519:16814 chr7 5449382 N chr7 5449503 N DUP 9
A00404:155:HV27LDSXX:3:1237:18828:33943 chr7 5449370 N chr7 5449461 N DUP 9
A00297:158:HT275DSXX:3:1613:29776:36213 chr7 5449384 N chr7 5449609 N DUP 21
A00404:156:HV37TDSXX:4:2640:8712:10347 chr7 5449375 N chr7 5449432 N DUP 7
A00404:156:HV37TDSXX:3:1638:1588:29825 chr7 5449370 N chr7 5449431 N DUP 9
A00404:155:HV27LDSXX:4:1602:13449:4335 chr7 5449375 N chr7 5449432 N DUP 7
A00404:155:HV27LDSXX:2:1678:16848:34084 chr7 5449382 N chr7 5449473 N DUP 9
A00404:156:HV37TDSXX:3:1601:8603:19460 chr7 5449384 N chr7 5449609 N DUP 24
A00404:156:HV37TDSXX:2:1268:28854:6496 chr7 5449400 N chr7 5449461 N DUP 9
A00404:155:HV27LDSXX:3:2647:5855:29168 chr7 5449400 N chr7 5449505 N DUP 5
A00404:156:HV37TDSXX:4:1319:9399:27195 chr7 5449400 N chr7 5449491 N DUP 9
A00297:158:HT275DSXX:1:2148:14371:32581 chr7 5449370 N chr7 5449431 N DUP 9
A00404:155:HV27LDSXX:3:2551:10185:8891 chr7 5449370 N chr7 5449491 N DUP 9
A00404:155:HV27LDSXX:4:1333:7771:18865 chr7 5449375 N chr7 5449612 N DUP 12
A00404:155:HV27LDSXX:1:1127:29405:12461 chr7 5449541 N chr7 5449610 N DUP 13
A00297:158:HT275DSXX:2:1676:31376:21386 chr7 5449404 N chr7 5449597 N DEL 19
A00404:156:HV37TDSXX:2:1351:29053:27665 chr7 5449409 N chr7 5449602 N DEL 9
A00297:158:HT275DSXX:1:1127:18159:20322 chr7 5449396 N chr7 5449621 N DEL 5
A00404:156:HV37TDSXX:1:1111:12924:6715 chr7 5449397 N chr7 5449622 N DEL 5
A00404:155:HV27LDSXX:1:2307:4526:3724 chr7 5449397 N chr7 5449622 N DEL 5
A00297:158:HT275DSXX:3:2511:21829:20384 chr17 82959093 N chr17 82959185 N DEL 10
A00297:158:HT275DSXX:3:2639:27308:34569 chr17 82959082 N chr17 82959174 N DEL 12
A00404:155:HV27LDSXX:1:2670:7609:26663 chr17 82959106 N chr17 82959198 N DEL 2
A00404:155:HV27LDSXX:4:1624:18602:32080 chr17 82959137 N chr17 82959283 N DEL 16
A00404:155:HV27LDSXX:2:2404:14814:29997 chr16 86857918 N chr16 86858092 N DUP 10
A00297:158:HT275DSXX:4:1220:13241:2127 chr16 86857919 N chr16 86858093 N DUP 8
A00297:158:HT275DSXX:3:2115:22869:5682 chr4 3617620 N chr4 3617843 N DEL 37
A00404:156:HV37TDSXX:2:2112:10827:20995 chr8 97587486 N chr8 97587543 N DEL 11
A00297:158:HT275DSXX:2:2248:29622:8860 chr8 97587500 N chr8 97587583 N DEL 21
A00404:155:HV27LDSXX:4:1211:8052:23171 chr8 97587518 N chr8 97587603 N DUP 15
A00297:158:HT275DSXX:1:2234:13376:25473 chr8 97587518 N chr8 97587603 N DUP 16
A00404:155:HV27LDSXX:4:1372:10926:10488 chr8 97587517 N chr8 97587602 N DUP 5
A00404:156:HV37TDSXX:3:1631:23249:33802 chr8 97587538 N chr8 97587665 N DUP 9
A00404:156:HV37TDSXX:1:2677:19705:15765 chr8 97587538 N chr8 97587665 N DUP 7
A00404:156:HV37TDSXX:2:1341:7780:1282 chr8 97587517 N chr8 97587674 N DUP 10
A00297:158:HT275DSXX:2:2202:13485:23375 chr8 97587548 N chr8 97587603 N DEL 7
A00404:156:HV37TDSXX:3:2534:3568:4633 chr8 97587604 N chr8 97587681 N DEL 18
A00404:156:HV37TDSXX:4:2254:29622:27993 chr8 97587571 N chr8 97587672 N DEL 19
A00404:155:HV27LDSXX:1:2209:27462:22999 chr8 97587606 N chr8 97587683 N DEL 16
A00297:158:HT275DSXX:3:2601:5999:13823 chr8 97587616 N chr8 97587693 N DEL 10
A00404:155:HV27LDSXX:1:2164:2618:18834 chr8 97587574 N chr8 97587675 N DEL 7
A00404:156:HV37TDSXX:4:1267:2555:10645 chr8 97587584 N chr8 97587689 N DEL 7
A00404:155:HV27LDSXX:2:1525:14371:31078 chr8 97587535 N chr8 97587696 N DEL 4
A00404:155:HV27LDSXX:2:1572:21278:5713 chr8 97587537 N chr8 97587698 N DEL 2
A00404:156:HV37TDSXX:1:1340:16740:14356 chr15 45293406 N chr15 45293521 N DUP 4
A00404:155:HV27LDSXX:4:2125:7862:2174 chr15 45293502 N chr15 45293581 N DUP 1
A00297:158:HT275DSXX:3:2341:23565:9706 chr7 74496270 N chr7 74496421 N DEL 5
A00404:155:HV27LDSXX:4:2207:3902:23844 chr3 262084 N chr3 262533 N DUP 1
A00404:155:HV27LDSXX:4:2408:10592:13542 chr3 262084 N chr3 262533 N DUP 1
A00404:155:HV27LDSXX:1:2601:3486:9940 chr3 262085 N chr3 262401 N DEL 5
A00404:156:HV37TDSXX:1:1319:30553:32612 chr3 262123 N chr3 262574 N DEL 5
A00404:156:HV37TDSXX:2:1467:27154:34585 chr3 262096 N chr3 262680 N DUP 5
A00297:158:HT275DSXX:2:1101:27995:29716 chr3 262123 N chr3 262529 N DEL 5
A00404:156:HV37TDSXX:3:1678:25382:20243 chr3 262123 N chr3 262529 N DEL 5
A00404:155:HV27LDSXX:3:1327:30337:27853 chr3 262096 N chr3 262680 N DUP 5
A00404:155:HV27LDSXX:3:1143:11731:6339 chr3 262123 N chr3 262529 N DEL 5
A00404:155:HV27LDSXX:1:2344:4517:11287 chr3 262123 N chr3 262529 N DEL 5
A00404:155:HV27LDSXX:2:2239:4056:33160 chr3 262096 N chr3 262680 N DUP 5
A00404:155:HV27LDSXX:4:1539:30789:9157 chr3 262079 N chr3 262528 N DUP 5
A00404:155:HV27LDSXX:2:2460:5050:15624 chr3 262123 N chr3 262529 N DEL 5
A00404:156:HV37TDSXX:3:1304:16902:31109 chr3 262168 N chr3 262529 N DEL 5
A00297:158:HT275DSXX:2:1122:15365:14826 chr3 262073 N chr3 262162 N DUP 5
A00297:158:HT275DSXX:3:2504:3812:15139 chr3 262123 N chr3 262574 N DEL 5
A00404:155:HV27LDSXX:3:1327:30337:27853 chr3 262123 N chr3 262574 N DEL 5
A00404:156:HV37TDSXX:3:2457:22453:22498 chr3 262134 N chr3 262585 N DEL 4
A00404:156:HV37TDSXX:3:2457:22462:23359 chr3 262134 N chr3 262585 N DEL 4
A00404:156:HV37TDSXX:4:2667:3604:34194 chr3 262096 N chr3 262680 N DUP 5
A00404:156:HV37TDSXX:2:2609:6189:34820 chr3 262123 N chr3 262574 N DEL 5
A00404:155:HV27LDSXX:4:1155:12581:2613 chr3 262439 N chr3 262528 N DUP 5
A00297:158:HT275DSXX:3:1469:6325:35556 chr3 262087 N chr3 262403 N DEL 5
A00404:155:HV27LDSXX:4:2207:3902:23844 chr3 262168 N chr3 262529 N DEL 2
A00404:155:HV27LDSXX:3:1563:2781:34804 chr3 262484 N chr3 262573 N DUP 10
A00404:155:HV27LDSXX:3:1541:9435:22122 chr3 262484 N chr3 262573 N DUP 10
A00404:155:HV27LDSXX:4:2213:28926:4241 chr3 262484 N chr3 262573 N DUP 9
A00404:155:HV27LDSXX:2:2478:25247:26271 chr3 262123 N chr3 262529 N DEL 5
A00404:155:HV27LDSXX:2:2268:27371:11005 chr3 262125 N chr3 262531 N DEL 5
A00297:158:HT275DSXX:4:1227:28971:5760 chr3 262168 N chr3 262529 N DEL 5
A00404:155:HV27LDSXX:4:2155:9236:10379 chr3 262130 N chr3 262536 N DEL 5
A00297:158:HT275DSXX:3:1407:5647:6292 chr3 262484 N chr3 262573 N DUP 10
A00404:156:HV37TDSXX:2:2436:20654:26146 chr3 262484 N chr3 262573 N DUP 6
A00404:155:HV27LDSXX:3:1302:28682:14810 chr3 262092 N chr3 262498 N DEL 1
A00297:158:HT275DSXX:1:2447:32579:26412 chr3 262123 N chr3 262529 N DEL 5
A00404:155:HV27LDSXX:4:2625:8947:11005 chr3 262123 N chr3 262529 N DEL 5
A00404:155:HV27LDSXX:3:1544:26720:25441 chr3 262082 N chr3 262531 N DUP 3
A00404:155:HV27LDSXX:3:1563:2781:34804 chr3 262082 N chr3 262531 N DUP 3
A00404:155:HV27LDSXX:3:1541:9435:22122 chr3 262484 N chr3 262573 N DUP 10
A00297:158:HT275DSXX:2:1402:16360:18991 chr3 262110 N chr3 262559 N DUP 2
A00404:155:HV27LDSXX:3:1143:11731:6339 chr3 262081 N chr3 262530 N DUP 4
A00297:158:HT275DSXX:1:2365:5801:16235 chr3 262128 N chr3 262579 N DEL 5
A00404:155:HV27LDSXX:1:1271:31765:23156 chr3 262129 N chr3 262580 N DEL 5
A00404:155:HV27LDSXX:1:1271:32081:23328 chr3 262129 N chr3 262580 N DEL 5
A00404:155:HV27LDSXX:1:1271:32090:23312 chr3 262129 N chr3 262580 N DEL 5
A00297:158:HT275DSXX:4:1313:9525:24596 chr3 262140 N chr3 262681 N DEL 10
A00297:158:HT275DSXX:4:1313:9525:24596 chr3 262140 N chr3 262681 N DEL 6
A00404:156:HV37TDSXX:2:1157:32479:25394 chr3 262140 N chr3 262681 N DEL 5
A00404:156:HV37TDSXX:1:2522:29532:9111 chr7 80932003 N chr7 80932084 N DUP 10
A00404:156:HV37TDSXX:2:1270:16676:20917 chr6 167590510 N chr6 167590625 N DUP 5
A00404:156:HV37TDSXX:2:2356:29658:24267 chr6 167590366 N chr6 167590612 N DUP 5
A00297:158:HT275DSXX:1:1271:15148:6120 chr6 167590366 N chr6 167590612 N DUP 5
A00404:155:HV27LDSXX:3:1570:18123:19413 chr6 167590399 N chr6 167590519 N DEL 5
A00404:156:HV37TDSXX:3:2250:4047:13197 chr6 167590549 N chr6 167590676 N DUP 5
A00404:156:HV37TDSXX:1:2541:17381:3787 chr6 167590366 N chr6 167590612 N DUP 5
A00404:156:HV37TDSXX:3:2301:25798:32581 chr6 167590605 N chr6 167590732 N DUP 27
A00404:156:HV37TDSXX:4:1238:9037:33019 chr6 167590604 N chr6 167590737 N DEL 36
A00404:155:HV27LDSXX:4:2663:22525:20995 chr6 167590549 N chr6 167590676 N DUP 10
A00404:155:HV27LDSXX:1:2578:12228:18443 chr6 167590558 N chr6 167590685 N DUP 5
A00297:158:HT275DSXX:2:1321:13096:31751 chr6 167590605 N chr6 167590732 N DUP 18
A00404:155:HV27LDSXX:3:2404:29396:20369 chr6 167590440 N chr6 167590560 N DEL 2
A00297:158:HT275DSXX:1:1363:26160:29888 chr6 167590560 N chr6 167590687 N DUP 4
A00297:158:HT275DSXX:3:2271:27353:4335 chr6 167590549 N chr6 167590676 N DUP 1
A00297:158:HT275DSXX:3:1674:26332:18912 chr6 167590626 N chr6 167590871 N DUP 2
A00297:158:HT275DSXX:1:1246:15320:31469 chr6 167590549 N chr6 167590676 N DUP 7
A00404:155:HV27LDSXX:2:2647:12671:12571 chr6 167590549 N chr6 167590676 N DUP 34
A00404:156:HV37TDSXX:2:2134:17119:21997 chr6 167590549 N chr6 167590676 N DUP 36
A00404:156:HV37TDSXX:3:1263:13602:21198 chr6 167590549 N chr6 167590676 N DUP 34
A00404:156:HV37TDSXX:1:1269:18837:25974 chr6 167590744 N chr6 167590857 N DUP 5
A00404:156:HV37TDSXX:3:2552:30400:23610 chr6 167590745 N chr6 167590858 N DUP 5
A00404:156:HV37TDSXX:4:2604:15510:35587 chr6 167590615 N chr6 167590748 N DEL 4
A00404:156:HV37TDSXX:3:2556:11550:35775 chr15 33336576 N chr15 33336641 N DEL 2
A00297:158:HT275DSXX:1:1310:14488:24392 chr15 33336577 N chr15 33336634 N DEL 6
A00297:158:HT275DSXX:2:1667:25852:8030 chr9 136718306 N chr9 136718379 N DEL 7
A00404:155:HV27LDSXX:1:1646:32886:35055 chr9 136718306 N chr9 136718379 N DEL 7
A00404:156:HV37TDSXX:1:2528:15890:2550 chr9 136718306 N chr9 136718379 N DEL 8
A00404:156:HV37TDSXX:4:1460:7139:6402 chr9 136718306 N chr9 136718379 N DEL 11
A00404:156:HV37TDSXX:1:2278:8929:33144 chr9 136718306 N chr9 136718379 N DEL 14
A00404:156:HV37TDSXX:1:2278:9543:31798 chr9 136718306 N chr9 136718379 N DEL 14
A00404:156:HV37TDSXX:1:1359:11134:13761 chr9 136718261 N chr9 136718370 N DEL 32
A00404:156:HV37TDSXX:2:1366:26982:20979 chr9 136718331 N chr9 136718404 N DEL 29
A00404:155:HV27LDSXX:4:1455:22444:19570 chr9 136718331 N chr9 136718404 N DEL 27
A00404:156:HV37TDSXX:2:1457:14904:18035 chr9 136718331 N chr9 136718404 N DEL 22
A00404:156:HV37TDSXX:2:2457:16260:25927 chr9 136718331 N chr9 136718404 N DEL 22
A00404:155:HV27LDSXX:2:2407:8350:19680 chr9 136718331 N chr9 136718404 N DEL 14
A00297:158:HT275DSXX:2:2264:17996:22921 chr9 136718332 N chr9 136718405 N DEL 6
A00297:158:HT275DSXX:3:1475:7057:8359 chr9 136718334 N chr9 136718407 N DEL 5
A00297:158:HT275DSXX:1:1435:7066:23156 chr9 136718337 N chr9 136718410 N DEL 5
A00297:158:HT275DSXX:3:2144:32398:26475 chr9 136718341 N chr9 136718414 N DEL 5
A00404:155:HV27LDSXX:2:2401:5782:7999 chr9 136718342 N chr9 136718415 N DEL 4
A00297:158:HT275DSXX:4:1619:17897:12132 chr4 2244069 N chr4 2244154 N DUP 2
A00404:156:HV37TDSXX:3:1471:4119:35086 chr4 2244055 N chr4 2244192 N DEL 4
A00297:158:HT275DSXX:4:2462:16984:15969 chr2 90326300 N chr2 90326460 N DEL 4
A00297:158:HT275DSXX:4:2223:17589:12696 chr2 90326308 N chr2 90326466 N DUP 4
A00404:155:HV27LDSXX:1:1337:21676:9659 chr17 44405599 N chr17 44405896 N DEL 5
A00404:155:HV27LDSXX:1:1337:21676:9659 chr17 44405599 N chr17 44405896 N DEL 15
A00404:155:HV27LDSXX:3:2133:19407:11428 chr15 84240344 N chr15 84240408 N DEL 4
A00404:155:HV27LDSXX:3:2542:11695:18427 chr15 84240516 N chr15 84240595 N DEL 5
A00404:156:HV37TDSXX:4:1620:1443:30859 chr15 84240523 N chr15 84240602 N DEL 5
A00404:156:HV37TDSXX:1:1573:4354:34021 chr15 40136443 N chr15 40136593 N DEL 5
A00404:155:HV27LDSXX:2:1107:22562:6245 chr14 86287220 N chr14 86287285 N DEL 15
A00404:155:HV27LDSXX:2:2107:20564:14873 chr14 86287220 N chr14 86287285 N DEL 15
A00404:155:HV27LDSXX:4:1123:24017:23547 chr14 86287220 N chr14 86287285 N DEL 25
A00404:155:HV27LDSXX:1:1405:18267:6324 chr14 86287220 N chr14 86287285 N DEL 22
A00404:155:HV27LDSXX:4:2219:29595:36401 chr12 70203032 N chr12 70203285 N DUP 9
A00297:158:HT275DSXX:2:1378:29487:35368 chr12 70203111 N chr12 70203238 N DEL 5
A00297:158:HT275DSXX:1:2450:19180:22592 chr12 70202916 N chr12 70203342 N DEL 6
A00297:158:HT275DSXX:3:2306:27588:10974 chr12 70202927 N chr12 70203353 N DEL 4
A00404:155:HV27LDSXX:1:1246:10140:14262 chr2 167201290 N chr2 167201357 N DEL 12
A00404:155:HV27LDSXX:4:1334:21233:10864 chr2 167201423 N chr2 167201482 N DUP 38
A00404:155:HV27LDSXX:4:2151:31458:14732 chr2 167201423 N chr2 167201482 N DUP 33
A00297:158:HT275DSXX:1:2515:10529:34006 chr2 167201436 N chr2 167201499 N DUP 2
A00404:155:HV27LDSXX:3:1261:18692:22310 chr2 167201427 N chr2 167201486 N DUP 11
A00404:156:HV37TDSXX:4:2431:19813:21433 chr2 167201427 N chr2 167201486 N DUP 11
A00297:158:HT275DSXX:3:2632:29243:3881 chr19 50975316 N chr19 50975766 N DEL 23
A00404:155:HV27LDSXX:4:2378:14597:28776 chr19 50975233 N chr19 50975401 N DEL 3
A00404:155:HV27LDSXX:3:1301:30544:16376 chr8 6177587 N chr8 6177732 N DEL 5
A00297:158:HT275DSXX:3:2129:4996:1219 chr8 6177587 N chr8 6177732 N DEL 5
A00404:155:HV27LDSXX:1:2570:9028:26553 chr8 6177587 N chr8 6177732 N DEL 5
A00297:158:HT275DSXX:1:1145:14163:5196 chr8 6177520 N chr8 6177593 N DEL 1
A00297:158:HT275DSXX:1:1145:14226:10629 chr8 6177520 N chr8 6177593 N DEL 1
A00404:155:HV27LDSXX:1:1158:14498:16391 chr8 6177513 N chr8 6177586 N DEL 3
A00297:158:HT275DSXX:3:2117:30752:20964 chr8 6177513 N chr8 6177586 N DEL 3
A00404:156:HV37TDSXX:1:1537:13467:5087 chr8 6177525 N chr8 6177708 N DUP 7
A00404:156:HV37TDSXX:4:2409:22987:28150 chr8 6177626 N chr8 6177734 N DEL 13
A00404:155:HV27LDSXX:2:2339:20672:7044 chr8 6177517 N chr8 6177734 N DEL 13
A00404:156:HV37TDSXX:4:2353:12843:29496 chr8 6177520 N chr8 6177737 N DEL 12
A00297:158:HT275DSXX:2:1329:30834:25175 chr8 6177602 N chr8 6177747 N DEL 2
A00297:158:HT275DSXX:3:2130:1389:7560 chr10 133156878 N chr10 133156979 N DEL 5
A00404:155:HV27LDSXX:2:2263:11433:7200 chr2 238902672 N chr2 238903809 N DEL 9
A00404:155:HV27LDSXX:3:1367:26883:32080 chr2 238902676 N chr2 238903804 N DEL 10
A00297:158:HT275DSXX:3:1439:30472:29309 chr2 238902679 N chr2 238903805 N DEL 10
A00297:158:HT275DSXX:4:2608:3649:22185 chr2 238902706 N chr2 238903806 N DEL 5
A00404:156:HV37TDSXX:2:2210:11975:1125 chr2 238902727 N chr2 238903808 N DEL 5
A00404:156:HV37TDSXX:4:1555:3468:8343 chr2 238902728 N chr2 238903804 N DEL 8
A00404:155:HV27LDSXX:1:1140:11496:31328 chr2 238902741 N chr2 238903803 N DEL 7
A00404:155:HV27LDSXX:1:2666:2392:17347 chr2 238902749 N chr2 238903819 N DUP 5
A00297:158:HT275DSXX:3:1369:1895:20932 chr2 238902757 N chr2 238903808 N DEL 5
A00404:155:HV27LDSXX:3:1566:25771:15060 chr2 238902766 N chr2 238903809 N DEL 10
A00297:158:HT275DSXX:2:2547:28682:7451 chr2 238902794 N chr2 238903808 N DEL 4
A00404:156:HV37TDSXX:2:2578:1958:11710 chr2 238902800 N chr2 238903804 N DEL 5
A00297:158:HT275DSXX:4:2139:22679:2754 chr2 238902821 N chr2 238903807 N DEL 7
A00404:156:HV37TDSXX:4:2271:1904:15468 chr2 238902813 N chr2 238903809 N DEL 7
A00404:155:HV27LDSXX:2:2451:29243:4883 chr2 238902831 N chr2 238903806 N DEL 5
A00297:158:HT275DSXX:4:2139:22679:2754 chr2 238902839 N chr2 238903809 N DEL 6
A00404:155:HV27LDSXX:1:2370:5737:8891 chr2 238902850 N chr2 238903797 N DEL 5
A00404:155:HV27LDSXX:3:1268:12391:6918 chr2 238902859 N chr2 238903804 N DEL 6
A00297:158:HT275DSXX:3:2437:20491:4476 chr2 238902893 N chr2 238903802 N DEL 7
A00404:155:HV27LDSXX:2:2519:27624:5087 chr2 238902911 N chr2 238903793 N DEL 10
A00297:158:HT275DSXX:4:2562:27010:19210 chr2 238902825 N chr2 238903809 N DEL 7
A00297:158:HT275DSXX:3:1441:1018:19570 chr2 238902989 N chr2 238903809 N DEL 7
A00297:158:HT275DSXX:3:2437:20491:4476 chr2 238903005 N chr2 238903808 N DEL 5
A00404:156:HV37TDSXX:2:2251:4924:14967 chr2 238903007 N chr2 238903809 N DEL 6
A00404:155:HV27LDSXX:4:1373:7663:27821 chr2 238902912 N chr2 238903808 N DEL 10
A00297:158:HT275DSXX:4:1574:18593:21449 chr2 238902869 N chr2 238903809 N DEL 5
A00297:158:HT275DSXX:1:1271:9353:4257 chr2 238902822 N chr2 238903804 N DEL 7
A00404:156:HV37TDSXX:4:2426:27245:15765 chr2 238902869 N chr2 238903803 N DEL 5
A00297:158:HT275DSXX:2:2207:6207:28213 chr2 238902920 N chr2 238903802 N DEL 6
A00404:156:HV37TDSXX:2:1415:17092:24706 chr2 238902836 N chr2 238903804 N DEL 6
A00404:155:HV27LDSXX:1:2322:19967:30154 chr2 238902831 N chr2 238903806 N DEL 5
A00404:156:HV37TDSXX:3:2677:23610:27665 chr2 238903041 N chr2 238903809 N DEL 6
A00404:156:HV37TDSXX:3:2677:23610:27665 chr2 238903032 N chr2 238903342 N DEL 5
A00297:158:HT275DSXX:1:1212:31015:8766 chr2 238903357 N chr2 238903809 N DEL 10
A00404:156:HV37TDSXX:4:2412:21305:31438 chr2 238903383 N chr2 238903809 N DEL 10
A00297:158:HT275DSXX:1:1271:9353:4257 chr2 238903404 N chr2 238903809 N DEL 7
A00404:155:HV27LDSXX:3:1653:14714:35587 chr2 238903442 N chr2 238903806 N DEL 4
A00404:156:HV37TDSXX:1:1245:19741:10160 chr2 238903442 N chr2 238903804 N DEL 5
A00404:155:HV27LDSXX:1:1658:22390:18349 chr2 238903461 N chr2 238903808 N DEL 5
A00297:158:HT275DSXX:2:2448:7907:16219 chr2 238903505 N chr2 238903809 N DEL 7
A00297:158:HT275DSXX:1:2351:9100:8265 chr2 238903521 N chr2 238903808 N DEL 5
A00297:158:HT275DSXX:4:1323:11704:22013 chr2 238903560 N chr2 238903820 N DUP 5
A00404:155:HV27LDSXX:1:2464:26765:5885 chr2 238902826 N chr2 238903809 N DEL 1
A00404:155:HV27LDSXX:1:2312:30852:16783 chr2 238903606 N chr2 238903800 N DEL 9
A00404:155:HV27LDSXX:3:1134:18927:34679 chr2 238903622 N chr2 238903814 N DUP 4
A00404:156:HV37TDSXX:1:2229:6659:29935 chr2 238902815 N chr2 238903808 N DEL 7
A00404:155:HV27LDSXX:2:2636:10700:31078 chr2 238903430 N chr2 238903808 N DEL 5
A00297:158:HT275DSXX:2:1413:21730:25473 chr4 123538674 N chr4 123538835 N DEL 5
A00297:158:HT275DSXX:4:2117:22742:4398 chr4 123538674 N chr4 123538835 N DEL 5
A00404:156:HV37TDSXX:3:2663:26323:1235 chr4 123538674 N chr4 123538835 N DEL 5
A00404:156:HV37TDSXX:3:2663:26621:1783 chr4 123538674 N chr4 123538835 N DEL 5
A00297:158:HT275DSXX:1:2268:29731:36417 chr4 123538674 N chr4 123538835 N DEL 5
A00404:155:HV27LDSXX:3:1545:18846:5447 chr4 123538693 N chr4 123538852 N DUP 5
A00297:158:HT275DSXX:4:2309:30662:8061 chr4 123538584 N chr4 123538704 N DEL 4
A00404:155:HV27LDSXX:4:2513:1976:1376 chr4 123538585 N chr4 123538705 N DEL 3
A00404:156:HV37TDSXX:1:1126:1886:24768 chr2 6184498 N chr2 6184589 N DUP 21
A00297:158:HT275DSXX:4:1419:21730:6214 chr2 6184498 N chr2 6184589 N DUP 21
A00404:155:HV27LDSXX:1:1167:27679:3803 chr2 6184498 N chr2 6184589 N DUP 21
A00297:158:HT275DSXX:2:1116:2510:13291 chr2 6184515 N chr2 6184592 N DEL 7
A00404:156:HV37TDSXX:2:2365:8730:32205 chr16 67222611 N chr16 67222779 N DUP 3
A00404:156:HV37TDSXX:1:1428:24460:32487 chr16 67222610 N chr16 67222778 N DEL 4
A00404:156:HV37TDSXX:1:2602:9480:24111 chr10 71869450 N chr10 71869625 N DUP 10
A00404:155:HV27LDSXX:3:1119:27688:33004 chr22 10628951 N chr22 10629082 N DEL 2
A00404:156:HV37TDSXX:3:1335:15962:21621 chr22 10628951 N chr22 10629082 N DEL 4
A00404:155:HV27LDSXX:4:2230:7229:8938 chr22 10628951 N chr22 10629082 N DEL 5
A00404:155:HV27LDSXX:3:1326:31385:27508 chr22 10628977 N chr22 10629056 N DEL 10
A00404:156:HV37TDSXX:4:1568:21151:34679 chr21 44763814 N chr21 44763952 N DEL 5
A00404:156:HV37TDSXX:2:1458:18756:9455 chr21 44763821 N chr21 44763974 N DUP 11
A00297:158:HT275DSXX:1:1161:1723:34319 chr21 44763829 N chr21 44763982 N DUP 6
A00297:158:HT275DSXX:1:2409:26928:20948 chr21 44763940 N chr21 44764478 N DEL 10
A00404:155:HV27LDSXX:1:2163:18855:30671 chr21 44763821 N chr21 44764099 N DEL 23
A00404:155:HV27LDSXX:1:2163:18855:30671 chr21 44763821 N chr21 44764099 N DEL 17
A00297:158:HT275DSXX:2:2255:5864:33066 chr21 44763841 N chr21 44764102 N DEL 12
A00404:155:HV27LDSXX:3:2218:8196:20478 chr21 44764120 N chr21 44764242 N DEL 10
A00404:155:HV27LDSXX:1:2411:15212:34444 chr21 44764120 N chr21 44764242 N DEL 5
A00404:155:HV27LDSXX:2:2114:29550:5885 chr21 44763950 N chr21 44764400 N DUP 5
A00404:156:HV37TDSXX:4:1577:28348:16360 chr21 44764209 N chr21 44764537 N DEL 24
A00297:158:HT275DSXX:4:2510:17110:15342 chr16 3016774 N chr16 3016942 N DEL 39
A00404:156:HV37TDSXX:1:1561:13829:20744 chr2 3263812 N chr2 3263879 N DEL 8
A00297:158:HT275DSXX:3:1402:29722:5995 chr16 33619501 N chr16 33619582 N DEL 25
A00404:156:HV37TDSXX:1:2134:13160:15264 chr16 33619517 N chr16 33619620 N DEL 1
A00404:155:HV27LDSXX:2:2244:26232:11757 chr16 33619508 N chr16 33619653 N DEL 4
A00404:156:HV37TDSXX:4:2307:27733:33270 chr17 37565595 N chr17 37565868 N DEL 10
A00404:156:HV37TDSXX:2:1658:4128:10113 chr17 37565625 N chr17 37565700 N DUP 1
A00404:155:HV27LDSXX:4:1256:19750:8954 chr17 37565620 N chr17 37565775 N DUP 5
A00404:156:HV37TDSXX:2:1658:4128:10113 chr17 37565659 N chr17 37565851 N DUP 5
A00404:156:HV37TDSXX:1:2521:4752:6339 chr17 37565713 N chr17 37565947 N DEL 52
A00297:158:HT275DSXX:2:1212:11912:13573 chr3 8502417 N chr3 8502470 N DUP 9
A00404:156:HV37TDSXX:4:2462:29921:17644 chr3 8502417 N chr3 8502470 N DUP 9
A00404:156:HV37TDSXX:3:1318:16685:28228 chr3 8502497 N chr3 8502571 N DUP 26
A00404:156:HV37TDSXX:3:2663:23800:7200 chr3 8502408 N chr3 8502474 N DUP 17
A00297:158:HT275DSXX:3:2440:9516:2910 chrX 2224801 N chrX 2225106 N DUP 1
A00404:155:HV27LDSXX:4:2402:25970:5384 chrX 2224971 N chrX 2225104 N DUP 2
A00404:155:HV27LDSXX:2:2457:26277:16908 chr12 88715537 N chr12 88715586 N DUP 23
A00404:155:HV27LDSXX:2:1248:20509:14434 chr12 88715537 N chr12 88715586 N DUP 29
A00297:158:HT275DSXX:3:2603:26648:24752 chr12 88715537 N chr12 88715586 N DUP 21
A00404:155:HV27LDSXX:1:2127:8151:33677 chr12 88715537 N chr12 88715586 N DUP 38
A00404:155:HV27LDSXX:1:2127:8739:33755 chr12 88715537 N chr12 88715586 N DUP 38
A00404:155:HV27LDSXX:3:1462:23448:14763 chr20 51455973 N chr20 51456282 N DEL 11
A00404:156:HV37TDSXX:2:1101:13539:8688 chr20 51455980 N chr20 51456039 N DUP 2
A00404:155:HV27LDSXX:4:2178:4255:8453 chr20 51455924 N chr20 51456087 N DUP 10
A00297:158:HT275DSXX:2:1242:25889:25034 chr20 51455866 N chr20 51456093 N DUP 10
A00404:155:HV27LDSXX:2:2428:19153:30906 chr20 51456059 N chr20 51456110 N DUP 5
A00404:156:HV37TDSXX:3:1367:28908:36464 chr20 51455887 N chr20 51456056 N DEL 5
A00404:155:HV27LDSXX:4:2649:27299:16611 chr2 92080839 N chr2 92081178 N DUP 10
A00404:156:HV37TDSXX:1:1139:1741:12399 chr2 92080977 N chr2 92081146 N DUP 5
A00404:156:HV37TDSXX:3:2406:30644:2675 chr2 92080687 N chr2 92081162 N DEL 5
A00404:155:HV27LDSXX:1:2521:17879:21840 chr2 92080765 N chr2 92081178 N DEL 2
A00404:155:HV27LDSXX:3:1644:16821:14685 chr2 92080770 N chr2 92081435 N DEL 5
A00297:158:HT275DSXX:2:2153:15121:11741 chr18 36064664 N chr18 36064747 N DEL 1
A00297:158:HT275DSXX:3:2428:10357:30514 chr7 128361151 N chr7 128361266 N DEL 2
A00297:158:HT275DSXX:1:1319:4318:15358 chr17 1665460 N chr17 1665765 N DEL 10
A00297:158:HT275DSXX:3:1175:13006:27868 chr17 1665427 N chr17 1665732 N DEL 25
A00297:158:HT275DSXX:1:2511:27507:8641 chr17 1665981 N chr17 1666302 N DEL 10
A00404:155:HV27LDSXX:2:1343:27218:10958 chr21 7257635 N chr21 7257784 N DUP 5
A00404:155:HV27LDSXX:2:1343:27570:10848 chr21 7257635 N chr21 7257784 N DUP 5
A00297:158:HT275DSXX:3:1662:32497:35603 chr21 7257761 N chr21 7257830 N DUP 5
A00297:158:HT275DSXX:1:2343:8576:36636 chr21 7257761 N chr21 7257830 N DUP 6
A00404:155:HV27LDSXX:4:1423:8522:23923 chr21 7257690 N chr21 7257864 N DUP 2
A00404:155:HV27LDSXX:2:2378:24460:10254 chr21 7257690 N chr21 7257864 N DUP 3
A00404:155:HV27LDSXX:4:1559:3125:21183 chr21 7257690 N chr21 7257864 N DUP 4
A00297:158:HT275DSXX:3:2468:10077:29778 chr21 7257686 N chr21 7257885 N DUP 5
A00297:158:HT275DSXX:2:1213:14832:17534 chr21 7257686 N chr21 7257885 N DUP 5
A00404:156:HV37TDSXX:2:1571:16559:2456 chr21 7257903 N chr21 7257959 N DEL 5
A00404:156:HV37TDSXX:4:1378:6569:12618 chr7 45016564 N chr7 45016868 N DEL 28
A00404:156:HV37TDSXX:1:2508:10529:27211 chr7 45016564 N chr7 45016868 N DEL 27
A00404:156:HV37TDSXX:4:1378:6569:12618 chr7 45016564 N chr7 45016868 N DEL 20
A00404:155:HV27LDSXX:3:2146:3034:13730 chr7 45016623 N chr7 45016927 N DEL 5
A00404:156:HV37TDSXX:2:1338:21133:3270 chr12 1604910 N chr12 1604962 N DEL 5
A00404:155:HV27LDSXX:2:2201:18810:14058 chr16 28416953 N chr16 28417212 N DEL 2
A00404:156:HV37TDSXX:1:2342:30110:15843 chr16 28416895 N chr16 28416945 N DUP 5
A00297:158:HT275DSXX:3:2551:7464:35274 chr16 28416937 N chr16 28417065 N DUP 5
A00404:155:HV27LDSXX:3:1251:5647:31000 chr16 28416953 N chr16 28417212 N DEL 17
A00404:155:HV27LDSXX:4:2175:17237:15311 chr16 28417045 N chr16 28417302 N DEL 3
A00404:155:HV27LDSXX:1:2676:27353:2675 chr16 28416958 N chr16 28417086 N DUP 1
A00404:156:HV37TDSXX:2:2134:23683:24220 chr16 28417059 N chr16 28417367 N DEL 15
A00297:158:HT275DSXX:4:1547:2311:6464 chr16 28416924 N chr16 28417052 N DUP 5
A00297:158:HT275DSXX:1:1472:12762:10535 chr16 28416723 N chr16 28416972 N DEL 3
A00297:158:HT275DSXX:3:1233:7808:9533 chr16 28416844 N chr16 28417014 N DEL 10
A00297:158:HT275DSXX:2:2578:11993:33473 chr16 28417146 N chr16 28417276 N DEL 8
A00404:155:HV27LDSXX:1:1216:7482:29324 chr16 28416942 N chr16 28417200 N DUP 7
A00297:158:HT275DSXX:1:2645:30563:16219 chr16 28416942 N chr16 28417200 N DUP 7
A00404:155:HV27LDSXX:2:1265:3992:13041 chr16 28416942 N chr16 28417200 N DUP 7
A00297:158:HT275DSXX:1:1667:28330:3583 chr16 28416942 N chr16 28417200 N DUP 7
A00404:155:HV27LDSXX:1:2251:17725:18067 chr16 28416942 N chr16 28417200 N DUP 7
A00404:156:HV37TDSXX:4:1642:16251:35806 chr16 28416942 N chr16 28417200 N DUP 7
A00404:156:HV37TDSXX:4:1131:31096:24565 chr16 28417064 N chr16 28417143 N DEL 2
A00404:156:HV37TDSXX:2:2223:25039:25911 chr16 28417063 N chr16 28417142 N DEL 3
A00404:155:HV27LDSXX:3:2454:19922:19398 chr16 28416967 N chr16 28417226 N DEL 1
A00297:158:HT275DSXX:1:2303:30454:20823 chr16 28416966 N chr16 28417225 N DEL 2
A00297:158:HT275DSXX:1:2303:30807:21089 chr16 28416966 N chr16 28417225 N DEL 2
A00404:156:HV37TDSXX:4:2645:30120:26256 chr16 28416904 N chr16 28417292 N DEL 5
A00297:158:HT275DSXX:1:2267:10610:9784 chr16 28416905 N chr16 28417293 N DEL 5
A00404:156:HV37TDSXX:2:2134:23683:24220 chr16 28417059 N chr16 28417367 N DEL 10
A00404:156:HV37TDSXX:4:1423:9833:6370 chr13 49377943 N chr13 49378177 N DEL 5
A00297:158:HT275DSXX:3:2675:18358:30467 chr13 49378031 N chr13 49378345 N DEL 16
A00297:158:HT275DSXX:2:2660:4001:19914 chr13 49378282 N chr13 49378361 N DUP 7
A00404:155:HV27LDSXX:1:1267:5629:6699 chr12 107895241 N chr12 107895424 N DEL 5
A00404:156:HV37TDSXX:3:1141:32597:29606 chr12 107895241 N chr12 107895424 N DEL 5
A00404:155:HV27LDSXX:1:2116:7139:20901 chr12 107895259 N chr12 107895440 N DUP 4
A00404:156:HV37TDSXX:2:1337:29451:14794 chr12 107895259 N chr12 107895440 N DUP 4
A00404:156:HV37TDSXX:2:1272:6343:35994 chr2 89787877 N chr2 89787929 N DEL 5
A00404:156:HV37TDSXX:3:2421:10682:30639 chr2 89787856 N chr2 89787934 N DEL 5
A00404:155:HV27LDSXX:2:1107:24099:29919 chr10 37054888 N chr10 37054978 N DUP 16
A00404:156:HV37TDSXX:3:2178:19877:26710 chr7 109447778 N chr7 109447856 N DEL 10
A00404:156:HV37TDSXX:3:2178:20039:26804 chr7 109447778 N chr7 109447856 N DEL 10
A00297:158:HT275DSXX:2:2502:24026:32706 chr15 101757099 N chr15 101757189 N DUP 1
A00404:156:HV37TDSXX:2:1174:28601:24940 chr15 101757080 N chr15 101757170 N DUP 14
A00404:155:HV27LDSXX:3:1373:1380:27430 chr15 101757141 N chr15 101757231 N DUP 5
A00404:156:HV37TDSXX:4:1568:32470:19617 chr15 101757154 N chr15 101757493 N DEL 5
A00297:158:HT275DSXX:3:1352:1280:33364 chr15 101757179 N chr15 101757269 N DUP 2
A00404:155:HV27LDSXX:1:2604:26910:10989 chr15 101757096 N chr15 101757188 N DEL 3
A00297:158:HT275DSXX:1:2309:24352:13448 chr15 101757176 N chr15 101757266 N DUP 5
A00404:155:HV27LDSXX:2:1475:21676:32957 chr15 101757226 N chr15 101757316 N DUP 3
A00404:155:HV27LDSXX:1:1654:10710:18004 chr15 101757141 N chr15 101757233 N DEL 5
A00404:156:HV37TDSXX:3:1666:18050:31250 chr15 101757317 N chr15 101757654 N DUP 5
A00404:156:HV37TDSXX:3:1469:28076:29481 chr15 101757274 N chr15 101757364 N DUP 5
A00404:156:HV37TDSXX:3:1466:14470:2879 chr15 101757134 N chr15 101757317 N DEL 5
A00297:158:HT275DSXX:3:1452:19461:21512 chr15 101757144 N chr15 101757327 N DEL 10
A00297:158:HT275DSXX:3:1204:14488:24706 chr15 101757143 N chr15 101757326 N DEL 5
A00297:158:HT275DSXX:2:1352:4481:18677 chr15 101757263 N chr15 101757355 N DEL 15
A00297:158:HT275DSXX:3:2171:22761:34741 chr15 101757165 N chr15 101757348 N DEL 20
A00404:155:HV27LDSXX:1:1207:19334:27492 chr15 101757237 N chr15 101757329 N DEL 3
A00404:156:HV37TDSXX:1:1614:5222:4210 chr15 101757331 N chr15 101757395 N DUP 5
A00404:156:HV37TDSXX:1:2273:5168:14137 chr15 101757100 N chr15 101757437 N DUP 5
A00404:155:HV27LDSXX:2:1506:30499:23657 chr15 101757403 N chr15 101757495 N DEL 20
A00404:156:HV37TDSXX:1:2438:11053:10895 chr15 101757148 N chr15 101757485 N DUP 5
A00404:156:HV37TDSXX:1:2222:1931:23437 chr15 101757153 N chr15 101757401 N DEL 18
A00297:158:HT275DSXX:3:1640:5095:18865 chr15 101757175 N chr15 101757423 N DEL 15
A00404:156:HV37TDSXX:3:2664:11713:29857 chr15 101757492 N chr15 101757673 N DUP 10
A00404:155:HV27LDSXX:2:2559:23095:7701 chr15 101757495 N chr15 101757676 N DUP 10
A00404:156:HV37TDSXX:2:1658:6388:25520 chr15 101757156 N chr15 101757586 N DEL 7
A00404:156:HV37TDSXX:4:2156:32154:27398 chr12 39711793 N chr12 39711852 N DUP 7
A00404:155:HV27LDSXX:3:2224:13485:33082 chr12 39711966 N chr12 39712045 N DEL 5
A00404:155:HV27LDSXX:1:1125:27073:29403 chr13 91571938 N chr13 91572011 N DEL 1
A00404:155:HV27LDSXX:2:2522:2808:35289 chr13 91571931 N chr13 91572028 N DUP 9
A00404:156:HV37TDSXX:2:1442:4544:8797 chr13 91571989 N chr13 91572040 N DUP 21
A00404:155:HV27LDSXX:4:1246:21703:4476 chr13 91571989 N chr13 91572040 N DUP 20
A00404:155:HV27LDSXX:1:2150:11026:23281 chr13 91571989 N chr13 91572040 N DUP 13
A00404:155:HV27LDSXX:1:1578:15736:1532 chr13 91571989 N chr13 91572040 N DUP 17
A00404:155:HV27LDSXX:3:1137:29215:26694 chr13 91571989 N chr13 91572040 N DUP 13
A00404:155:HV27LDSXX:4:1317:3405:14591 chr13 69956029 N chr13 69956265 N DEL 2
A00404:155:HV27LDSXX:1:1561:3622:12806 chr7 36515749 N chr7 36515938 N DUP 5
A00404:156:HV37TDSXX:4:2536:16875:3912 chr7 36515812 N chr7 36516152 N DUP 1
A00404:155:HV27LDSXX:2:1446:29152:11835 chr13 22023401 N chr13 22023469 N DEL 5
A00404:155:HV27LDSXX:4:1536:17354:15890 chr13 22023354 N chr13 22023495 N DUP 19
A00404:156:HV37TDSXX:1:1241:32524:35462 chr13 22023354 N chr13 22023495 N DUP 19
A00404:156:HV37TDSXX:2:2466:21016:29434 chr13 22023317 N chr13 22023408 N DEL 5
A00404:155:HV27LDSXX:4:2302:9860:32189 chr13 22023548 N chr13 22023659 N DUP 13
A00404:156:HV37TDSXX:1:2129:4227:33833 chr13 22023551 N chr13 22023702 N DUP 10
A00404:156:HV37TDSXX:3:1537:20464:27164 chr13 22023547 N chr13 22023658 N DUP 14
A00404:156:HV37TDSXX:3:2121:13367:14309 chr13 22023606 N chr13 22023663 N DEL 10
A00297:158:HT275DSXX:2:2311:29197:4022 chr13 22023606 N chr13 22023663 N DEL 10
A00404:155:HV27LDSXX:3:1453:28122:23766 chr13 22023606 N chr13 22023663 N DEL 10
A00404:156:HV37TDSXX:3:1427:5132:16799 chr13 22023606 N chr13 22023663 N DEL 10
A00404:156:HV37TDSXX:2:2466:21016:29434 chr13 22023606 N chr13 22023663 N DEL 10
A00404:155:HV27LDSXX:3:2232:6858:19445 chr13 22023578 N chr13 22023663 N DEL 10
A00404:155:HV27LDSXX:4:1464:7817:24361 chr13 22023578 N chr13 22023663 N DEL 10
A00404:155:HV27LDSXX:4:1464:8314:25535 chr13 22023578 N chr13 22023663 N DEL 10
A00404:156:HV37TDSXX:4:1431:20934:4085 chr13 22023675 N chr13 22023735 N DUP 3
A00297:158:HT275DSXX:3:1178:9489:19366 chrX 124471342 N chrX 124471423 N DUP 2
A00404:156:HV37TDSXX:2:2626:14606:34303 chr7 6975720 N chr7 6975837 N DEL 5
A00404:155:HV27LDSXX:4:2575:20600:6856 chrX 24309854 N chrX 24309918 N DUP 12
A00404:155:HV27LDSXX:1:2123:14498:12978 chr6 62838344 N chr6 62838574 N DEL 2
A00404:155:HV27LDSXX:1:2123:18005:14137 chr6 62838344 N chr6 62838574 N DEL 2
A00404:156:HV37TDSXX:3:1637:11993:16814 chr6 62838577 N chr6 62838728 N DUP 2
A00297:158:HT275DSXX:3:1524:12283:20572 chr22 42538647 N chr22 42538779 N DEL 7
A00297:158:HT275DSXX:4:1401:19190:24612 chr22 20251649 N chr22 20251995 N DEL 5
A00404:156:HV37TDSXX:2:2149:21314:2957 chr22 20251863 N chr22 20252003 N DUP 5
A00404:155:HV27LDSXX:1:1443:1669:10927 chr22 20251850 N chr22 20252044 N DUP 2
A00404:156:HV37TDSXX:2:2127:2917:8234 chr22 20252027 N chr22 20252173 N DEL 5
A00297:158:HT275DSXX:4:2432:20763:7420 chr22 20252027 N chr22 20252173 N DEL 5
A00297:158:HT275DSXX:4:2432:22218:17550 chr22 20251730 N chr22 20252173 N DEL 7
A00404:155:HV27LDSXX:4:1673:17336:6433 chr1 143262745 N chr1 143262796 N DUP 1
A00404:155:HV27LDSXX:4:1661:29288:24126 chr1 143262759 N chr1 143262905 N DUP 5
A00404:156:HV37TDSXX:4:1211:11831:4507 chr1 143262701 N chr1 143262870 N DUP 10
A00297:158:HT275DSXX:2:1409:3134:8766 chr1 143262659 N chr1 143262782 N DUP 5
A00404:156:HV37TDSXX:2:1646:16794:19210 chr1 143262773 N chr1 143262893 N DUP 5
A00404:156:HV37TDSXX:2:1142:14705:23578 chr1 143262766 N chr1 143262912 N DUP 5
A00404:156:HV37TDSXX:3:2372:8124:34319 chr4 38753827 N chr4 38754015 N DUP 4
A00404:156:HV37TDSXX:3:2107:15519:19476 chr4 38753843 N chr4 38754033 N DEL 5
A00404:155:HV27LDSXX:3:1668:26874:35853 chr8 939201 N chr8 939313 N DEL 13
A00297:158:HT275DSXX:4:1473:19596:12258 chr8 939225 N chr8 939300 N DUP 5
A00404:155:HV27LDSXX:4:2213:29866:17769 chr8 939303 N chr8 939493 N DUP 5
A00297:158:HT275DSXX:3:1562:26386:6793 chr8 939303 N chr8 939982 N DEL 4
A00297:158:HT275DSXX:3:1613:30553:5650 chr8 939928 N chr8 940003 N DEL 4
A00297:158:HT275DSXX:2:2366:18023:29199 chr8 939202 N chr8 939351 N DUP 10
A00297:158:HT275DSXX:4:2656:27100:35274 chr8 939202 N chr8 939351 N DUP 10
A00297:158:HT275DSXX:3:1421:7283:15515 chr8 939202 N chr8 939275 N DUP 5
A00404:156:HV37TDSXX:1:1327:7048:3239 chr8 939266 N chr8 939945 N DEL 14
A00404:155:HV27LDSXX:4:1659:22290:7592 chr8 939351 N chr8 939993 N DEL 4
A00404:156:HV37TDSXX:1:1244:24008:5368 chr8 939504 N chr8 939994 N DEL 4
A00404:156:HV37TDSXX:1:2119:31919:34100 chrX 125321528 N chrX 125321842 N DUP 5
A00404:156:HV37TDSXX:2:1206:24758:34695 chrX 125321577 N chrX 125321956 N DEL 5
A00297:158:HT275DSXX:4:2334:32145:18490 chrX 125321580 N chrX 125321959 N DEL 9
A00297:158:HT275DSXX:4:2443:4960:17190 chrX 125322057 N chrX 125322367 N DEL 5
A00404:155:HV27LDSXX:3:1512:31222:24251 chrX 125321897 N chrX 125322207 N DEL 16
A00404:156:HV37TDSXX:2:1475:3821:27931 chrX 125321607 N chrX 125322232 N DEL 10
A00297:158:HT275DSXX:3:1575:2709:25347 chr11 57716621 N chr11 57716893 N DEL 10
A00404:155:HV27LDSXX:1:2635:15013:19319 chr11 57716621 N chr11 57716893 N DEL 5
A00297:158:HT275DSXX:3:1522:12192:2190 chr11 57716666 N chr11 57716938 N DEL 2
A00404:155:HV27LDSXX:3:2370:18530:4241 chr11 57716558 N chr11 57716684 N DUP 11
A00297:158:HT275DSXX:3:1515:3360:10848 chr11 57716561 N chr11 57716687 N DUP 2
A00404:155:HV27LDSXX:2:2406:26901:14481 chr11 57716667 N chr11 57716937 N DUP 5
A00404:156:HV37TDSXX:1:2249:18738:15562 chr11 57716538 N chr11 57716984 N DUP 7
A00404:155:HV27LDSXX:2:1458:18602:35493 chr11 57716667 N chr11 57716937 N DUP 6
A00404:155:HV27LDSXX:2:2458:14055:5447 chr11 57716667 N chr11 57716937 N DUP 6
A00404:155:HV27LDSXX:4:1578:1334:1078 chr11 57716667 N chr11 57716937 N DUP 5
A00297:158:HT275DSXX:4:1354:27932:5337 chr11 57716667 N chr11 57716937 N DUP 5
A00404:155:HV27LDSXX:2:1472:2844:36260 chr11 57716667 N chr11 57716937 N DUP 5
A00404:156:HV37TDSXX:2:2625:17662:13823 chr11 57716667 N chr11 57716937 N DUP 5
A00297:158:HT275DSXX:3:1252:7355:29042 chr11 57716538 N chr11 57716759 N DUP 5
A00297:158:HT275DSXX:1:2241:21097:9251 chr11 57716678 N chr11 57716948 N DUP 4
A00404:156:HV37TDSXX:4:2674:18249:32283 chr11 57716584 N chr11 57716758 N DEL 5
A00404:155:HV27LDSXX:3:2504:2058:32550 chr11 57716633 N chr11 57716856 N DEL 15
A00404:155:HV27LDSXX:2:1232:12346:9940 chr11 57716576 N chr11 57716848 N DEL 5
A00404:156:HV37TDSXX:1:1239:28185:31109 chr11 57716666 N chr11 57716938 N DEL 5
A00404:156:HV37TDSXX:1:1239:28185:31109 chr11 57716666 N chr11 57716938 N DEL 5
A00404:155:HV27LDSXX:1:1244:21667:29997 chr11 57716760 N chr11 57717035 N DEL 26
A00404:155:HV27LDSXX:1:1244:21667:29997 chr11 57716760 N chr11 57717035 N DEL 31
A00297:158:HT275DSXX:4:1534:30409:17926 chr10 130197490 N chr10 130197940 N DEL 14
A00404:156:HV37TDSXX:3:2563:31693:34679 chr10 130197531 N chr10 130197997 N DEL 26
A00297:158:HT275DSXX:2:2525:15646:1908 chr10 130197595 N chr10 130197939 N DEL 41
A00404:156:HV37TDSXX:1:1648:29631:23970 chr10 130197528 N chr10 130197668 N DUP 2
A00404:155:HV27LDSXX:3:1201:16929:4507 chr10 130197925 N chr10 130198026 N DUP 5
A00404:156:HV37TDSXX:2:2538:29613:10817 chr10 130197925 N chr10 130198026 N DUP 5
A00404:156:HV37TDSXX:4:2516:31458:32330 chr10 130197925 N chr10 130198026 N DUP 5
A00297:158:HT275DSXX:4:2409:13792:8437 chr10 130198058 N chr10 130198262 N DUP 5
A00297:158:HT275DSXX:2:2410:3821:28307 chr10 130197867 N chr10 130198072 N DEL 1
A00404:156:HV37TDSXX:2:2511:16993:16892 chr10 130197867 N chr10 130198072 N DEL 1
A00404:156:HV37TDSXX:2:2511:17291:17033 chr10 130197867 N chr10 130198072 N DEL 1
A00404:156:HV37TDSXX:3:1310:24569:29951 chr10 130197990 N chr10 130198300 N DEL 42
A00404:155:HV27LDSXX:2:2122:21423:21746 chr4 7076343 N chr4 7076461 N DEL 12
A00404:156:HV37TDSXX:2:1572:21197:8202 chr4 7076315 N chr4 7076416 N DUP 5
A00297:158:HT275DSXX:2:1215:11125:22169 chr4 7076315 N chr4 7076416 N DUP 6
A00404:155:HV27LDSXX:4:2403:13196:36746 chr4 7076331 N chr4 7076405 N DEL 14
A00404:155:HV27LDSXX:4:2403:17879:33927 chr4 7076331 N chr4 7076405 N DEL 14
A00404:156:HV37TDSXX:4:1573:6442:11271 chr4 7076332 N chr4 7076406 N DEL 11
A00404:156:HV37TDSXX:4:2546:19831:37027 chr4 7076335 N chr4 7076409 N DEL 10
A00297:158:HT275DSXX:2:2319:22137:21480 chr10 56083618 N chr10 56083683 N DUP 7
A00404:155:HV27LDSXX:4:1366:27661:32362 chr10 56083618 N chr10 56083683 N DUP 7
A00297:158:HT275DSXX:4:1114:13214:35117 chr10 56083618 N chr10 56083683 N DUP 7
A00404:156:HV37TDSXX:1:1563:22236:14418 chr10 56083618 N chr10 56083683 N DUP 7
A00297:158:HT275DSXX:3:1165:21567:24972 chr10 56083618 N chr10 56083683 N DUP 7
A00404:155:HV27LDSXX:4:2448:4065:18740 chr12 49880116 N chr12 49880463 N DUP 17
A00297:158:HT275DSXX:3:1444:11785:27821 chr12 49880116 N chr12 49880463 N DUP 17
A00404:155:HV27LDSXX:3:1669:4074:8672 chr12 49880116 N chr12 49880463 N DUP 17
A00404:155:HV27LDSXX:2:2267:18656:33113 chr12 49880117 N chr12 49880318 N DUP 14
A00404:155:HV27LDSXX:4:1570:1570:4053 chr12 49880118 N chr12 49880319 N DUP 13
A00404:156:HV37TDSXX:2:2258:8693:2112 chr12 49880122 N chr12 49880323 N DUP 9
A00404:155:HV27LDSXX:3:2458:5972:3035 chr12 49880104 N chr12 49880591 N DUP 3
A00297:158:HT275DSXX:2:1167:5629:36072 chr1 143216024 N chr1 143216176 N DUP 4
A00404:155:HV27LDSXX:1:2429:32687:22842 chr1 143215991 N chr1 143216165 N DUP 5
A00404:155:HV27LDSXX:1:1361:20817:1720 chr1 143216013 N chr1 143216113 N DUP 2
A00297:158:HT275DSXX:2:2507:30210:20776 chr1 143216042 N chr1 143216220 N DUP 5
A00297:158:HT275DSXX:3:1351:31937:2785 chr1 143216049 N chr1 143216227 N DUP 2
A00404:155:HV27LDSXX:4:2660:3712:17722 chr13 114007446 N chr13 114007519 N DUP 16
A00404:155:HV27LDSXX:3:2202:13069:3114 chr13 114007367 N chr13 114007499 N DEL 7
A00404:156:HV37TDSXX:2:1443:5565:28823 chr18 78449140 N chr18 78449258 N DEL 5
A00404:156:HV37TDSXX:1:1237:5791:16689 chr18 78449140 N chr18 78449258 N DEL 5
A00404:155:HV27LDSXX:3:1212:19226:24361 chr18 78449140 N chr18 78449258 N DEL 5
A00404:156:HV37TDSXX:4:2138:14000:6261 chr18 78449158 N chr18 78449274 N DUP 3
A00404:156:HV37TDSXX:4:2138:14525:6856 chr18 78449158 N chr18 78449274 N DUP 3
A00297:158:HT275DSXX:1:1201:10565:13839 chr6 89125947 N chr6 89126832 N DEL 1
A00404:155:HV27LDSXX:2:1303:27245:12070 chr6 89125947 N chr6 89126830 N DEL 3
A00297:158:HT275DSXX:1:1306:9561:21840 chr19 49818793 N chr19 49819127 N DEL 5
A00404:156:HV37TDSXX:1:1249:31204:17832 chr12 117103547 N chr12 117103658 N DUP 5
A00404:156:HV37TDSXX:2:1444:14751:9251 chr12 117103614 N chr12 117103815 N DUP 5
A00404:155:HV27LDSXX:4:1105:30138:23249 chr12 117103715 N chr12 117103772 N DEL 5
A00404:155:HV27LDSXX:4:1105:32190:21731 chr12 117103715 N chr12 117103772 N DEL 5
A00404:155:HV27LDSXX:3:1442:28899:5196 chr12 117103715 N chr12 117103772 N DEL 5
A00404:155:HV27LDSXX:2:1358:2465:23797 chr12 117103715 N chr12 117103772 N DEL 5
A00404:156:HV37TDSXX:4:1260:16966:25238 chr12 48842696 N chr12 48842823 N DUP 7
A00404:155:HV27LDSXX:3:1442:17101:24314 chr12 48842671 N chr12 48842799 N DEL 7
A00404:156:HV37TDSXX:4:1618:13566:7357 chr12 48842686 N chr12 48842863 N DEL 5
A00404:155:HV27LDSXX:3:1249:6867:36088 chr16 84355194 N chr16 84355259 N DEL 7
A00297:158:HT275DSXX:4:1347:26901:27508 chr16 84355197 N chr16 84355502 N DEL 6
A00297:158:HT275DSXX:2:2569:28113:34773 chr16 84355334 N chr16 84355651 N DEL 4
A00404:155:HV27LDSXX:4:1209:29875:14434 chr16 84355230 N chr16 84355385 N DUP 5
A00297:158:HT275DSXX:4:2418:30255:4382 chr16 84355405 N chr16 84355654 N DEL 18
A00404:155:HV27LDSXX:2:2131:24731:28072 chr16 84355222 N chr16 84355567 N DEL 33
A00297:158:HT275DSXX:2:1635:28890:7498 chr3 40377599 N chr3 40377658 N DUP 20
A00404:155:HV27LDSXX:2:1501:3341:5838 chr5 149393066 N chr5 149393184 N DEL 10
A00404:156:HV37TDSXX:2:1378:30047:6308 chr19 44490096 N chr19 44490226 N DEL 7
A00404:155:HV27LDSXX:4:2469:6207:20666 chr11 86110020 N chr11 86110136 N DEL 5
A00297:158:HT275DSXX:2:1312:6180:26381 chr17 68050482 N chr17 68050540 N DEL 13
A00404:155:HV27LDSXX:1:2444:15826:11929 chr9 75021532 N chr9 75021589 N DUP 9
A00404:156:HV37TDSXX:4:2636:8919:24612 chrX 991792 N chrX 991870 N DUP 5
A00297:158:HT275DSXX:3:1361:18991:32722 chr9 137560962 N chr9 137561129 N DEL 4
A00297:158:HT275DSXX:3:2270:14507:17065 chr14 105690875 N chr14 105691034 N DEL 3
A00404:156:HV37TDSXX:4:2665:6027:1157 chr19 7871057 N chr19 7871127 N DEL 9
A00297:158:HT275DSXX:1:1315:26033:28823 chr19 7871057 N chr19 7871127 N DEL 17
A00404:156:HV37TDSXX:2:2625:2718:5791 chr19 7871057 N chr19 7871127 N DEL 18
A00297:158:HT275DSXX:4:1535:11776:5948 chr19 7871069 N chr19 7871137 N DUP 4
A00404:156:HV37TDSXX:1:1524:23746:11365 chr19 7871057 N chr19 7871127 N DEL 14
A00404:155:HV27LDSXX:3:1426:3378:11381 chr19 7871067 N chr19 7871137 N DEL 5
A00404:155:HV27LDSXX:4:1455:6090:7811 chr4 26492708 N chr4 26492865 N DEL 18
A00404:156:HV37TDSXX:3:2331:18313:19429 chr4 26492811 N chr4 26492944 N DEL 8
A00297:158:HT275DSXX:4:1560:12644:7482 chr4 26492653 N chr4 26492944 N DEL 5
A00297:158:HT275DSXX:4:2559:4924:2973 chr4 26492653 N chr4 26492944 N DEL 5
A00297:158:HT275DSXX:2:1519:1570:1172 chr4 26492670 N chr4 26492969 N DEL 18
A00404:156:HV37TDSXX:4:2478:31810:17942 chr4 26492653 N chr4 26492944 N DEL 5
A00404:155:HV27LDSXX:1:1123:5547:13103 chr4 26492837 N chr4 26492978 N DEL 18
A00404:156:HV37TDSXX:4:1464:11867:13557 chr4 26492663 N chr4 26492954 N DEL 5
A00297:158:HT275DSXX:2:2343:8974:8359 chr4 26492832 N chr4 26492973 N DEL 11
A00297:158:HT275DSXX:3:2208:14796:33035 chr4 26492876 N chr4 26493009 N DEL 3
A00404:155:HV27LDSXX:3:1530:23728:28401 chr4 26492714 N chr4 26493015 N DEL 1
A00404:156:HV37TDSXX:4:2223:31177:35916 chr4 26492710 N chr4 26493011 N DEL 5
A00297:158:HT275DSXX:1:2409:7157:17174 chr19 29129394 N chr19 29129712 N DEL 55
A00404:155:HV27LDSXX:4:2666:23538:14450 chr17 80511368 N chr17 80511454 N DEL 5
A00404:156:HV37TDSXX:2:1410:28791:15280 chr17 80511219 N chr17 80511478 N DUP 5
A00404:155:HV27LDSXX:4:2275:4363:1939 chr6 69513003 N chr6 69513060 N DEL 1
A00297:158:HT275DSXX:4:1574:12717:18067 chr3 184414656 N chr3 184414768 N DEL 5
A00297:158:HT275DSXX:4:1574:12771:18255 chr3 184414656 N chr3 184414768 N DEL 5
A00404:155:HV27LDSXX:2:1459:23077:26177 chr3 184414821 N chr3 184414884 N DUP 5
A00297:158:HT275DSXX:1:1156:20817:9204 chr22 45228827 N chr22 45229060 N DEL 5
A00404:155:HV27LDSXX:4:1410:19533:26678 chr22 45228844 N chr22 45229076 N DEL 22
A00404:156:HV37TDSXX:2:2454:8703:20697 chr22 45228853 N chr22 45229198 N DEL 1
A00297:158:HT275DSXX:1:1221:19126:14168 chr22 45228853 N chr22 45229198 N DEL 23
A00404:155:HV27LDSXX:2:2312:15311:35681 chr22 45228909 N chr22 45229258 N DEL 12
A00404:155:HV27LDSXX:2:2313:18023:25692 chr22 45228909 N chr22 45229258 N DEL 12
A00297:158:HT275DSXX:1:2548:12906:35117 chr22 45228867 N chr22 45228948 N DEL 2
A00297:158:HT275DSXX:4:2174:19922:5431 chr22 45229164 N chr22 45229478 N DUP 34
A00297:158:HT275DSXX:4:2174:20094:5666 chr22 45229164 N chr22 45229478 N DUP 34
A00404:156:HV37TDSXX:3:1432:25030:33035 chr22 45229080 N chr22 45229274 N DUP 12
A00404:155:HV27LDSXX:4:1652:8332:24659 chr22 45228925 N chr22 45229311 N DUP 20
A00404:155:HV27LDSXX:2:2173:24822:13542 chr22 45228925 N chr22 45229229 N DUP 10
A00297:158:HT275DSXX:2:1231:26874:31031 chr22 45229204 N chr22 45229442 N DEL 25
A00404:155:HV27LDSXX:2:2174:25762:24815 chr22 45228860 N chr22 45229442 N DEL 18
A00404:155:HV27LDSXX:1:1137:23927:19413 chr22 45229206 N chr22 45229444 N DEL 13
A00404:156:HV37TDSXX:4:2209:12518:5384 chr22 45228891 N chr22 45229472 N DEL 12
A00404:156:HV37TDSXX:1:1131:5819:17300 chr22 45228987 N chr22 45229488 N DEL 7
A00404:155:HV27LDSXX:4:2535:5086:5572 chr22 45228847 N chr22 45229470 N DEL 17
A00404:155:HV27LDSXX:1:1318:3640:35853 chr22 45228847 N chr22 45229470 N DEL 15
A00404:155:HV27LDSXX:2:2475:31340:3787 chr22 45228907 N chr22 45229489 N DEL 5
A00297:158:HT275DSXX:3:2543:29071:3208 chr22 45228910 N chr22 45229492 N DEL 5
A00297:158:HT275DSXX:1:2114:27145:28213 chr22 45228883 N chr22 45229502 N DEL 1
A00297:158:HT275DSXX:4:1112:2908:14481 chr19 4355641 N chr19 4355776 N DEL 5
A00297:158:HT275DSXX:4:1469:27715:13855 chr19 4355641 N chr19 4355776 N DEL 5
A00404:156:HV37TDSXX:1:2603:23909:26741 chr19 4355641 N chr19 4355776 N DEL 5
A00404:155:HV27LDSXX:1:1445:6985:2910 chr19 4355661 N chr19 4355794 N DUP 5
A00297:158:HT275DSXX:1:1515:16107:24126 chr19 4355661 N chr19 4355794 N DUP 5
A00297:158:HT275DSXX:1:2177:28510:21840 chr19 4355661 N chr19 4355794 N DUP 5
A00404:156:HV37TDSXX:1:2649:14027:25629 chr19 4355667 N chr19 4355800 N DUP 5
A00404:155:HV27LDSXX:1:1275:28872:11569 chr19 4355675 N chr19 4355808 N DUP 1
A00297:158:HT275DSXX:1:2102:8594:27868 chr7 1870352 N chr7 1870785 N DEL 15
A00404:155:HV27LDSXX:4:2469:18222:26600 chr7 1870352 N chr7 1870785 N DEL 19
A00404:156:HV37TDSXX:3:1262:14009:16548 chr7 1870548 N chr7 1870777 N DEL 11
A00404:156:HV37TDSXX:2:2137:18376:31219 chr7 1870581 N chr7 1871346 N DEL 5
A00297:158:HT275DSXX:1:2562:3667:3740 chr7 1870582 N chr7 1871574 N DUP 10
A00404:155:HV27LDSXX:3:2163:21911:23657 chr7 1870584 N chr7 1871576 N DUP 10
A00404:156:HV37TDSXX:2:2362:6560:12195 chr7 1870638 N chr7 1870789 N DUP 5
A00297:158:HT275DSXX:2:1266:17508:5447 chr7 1870644 N chr7 1870820 N DUP 5
A00404:155:HV27LDSXX:3:2120:17390:15483 chr7 1870751 N chr7 1871389 N DEL 5
A00404:156:HV37TDSXX:3:2540:5195:17347 chr7 1870733 N chr7 1871091 N DEL 6
A00404:155:HV27LDSXX:3:1404:24894:16047 chr7 1870409 N chr7 1870664 N DEL 5
A00404:155:HV27LDSXX:3:2203:4517:18333 chr7 1870385 N chr7 1870666 N DEL 5
A00297:158:HT275DSXX:2:2302:4490:7106 chr7 1870659 N chr7 1870785 N DUP 24
A00297:158:HT275DSXX:3:2658:1796:22827 chr7 1870646 N chr7 1870799 N DEL 3
A00297:158:HT275DSXX:1:1516:16676:37043 chr7 1870873 N chr7 1871841 N DEL 5
A00404:155:HV27LDSXX:1:1604:2799:13322 chr7 1870659 N chr7 1870887 N DUP 5
A00297:158:HT275DSXX:1:2443:21341:26710 chr7 1870747 N chr7 1870924 N DUP 13
A00297:158:HT275DSXX:3:1341:32579:15984 chr7 1870650 N chr7 1870954 N DUP 22
A00404:156:HV37TDSXX:3:1262:14009:16548 chr7 1870650 N chr7 1870954 N DUP 26
A00404:155:HV27LDSXX:1:1632:29279:23234 chr7 1870650 N chr7 1870954 N DUP 26
A00404:156:HV37TDSXX:4:2573:17562:6731 chr7 1871029 N chr7 1871285 N DEL 8
A00404:155:HV27LDSXX:2:2113:11903:25269 chr7 1870801 N chr7 1870981 N DEL 26
A00297:158:HT275DSXX:1:2278:22643:30968 chr7 1870801 N chr7 1870981 N DEL 26
A00297:158:HT275DSXX:2:1437:24297:31391 chr7 1870420 N chr7 1871007 N DEL 26
A00404:155:HV27LDSXX:3:1203:8712:31078 chr7 1870735 N chr7 1871042 N DEL 10
A00297:158:HT275DSXX:4:1154:6623:12587 chr7 1870420 N chr7 1871132 N DUP 5
A00404:156:HV37TDSXX:2:2170:31114:28823 chr7 1870733 N chr7 1871091 N DEL 5
A00404:156:HV37TDSXX:4:1149:12608:29152 chr7 1870733 N chr7 1871091 N DEL 5
A00404:156:HV37TDSXX:3:2131:29288:19116 chr7 1871042 N chr7 1871194 N DUP 5
A00404:155:HV27LDSXX:4:1169:27588:31892 chr7 1870386 N chr7 1871100 N DEL 10
A00297:158:HT275DSXX:1:2278:22643:30968 chr7 1871157 N chr7 1871589 N DUP 5
A00297:158:HT275DSXX:1:2602:3459:33348 chr7 1871142 N chr7 1871574 N DUP 5
A00297:158:HT275DSXX:4:1125:29894:30185 chr7 1871004 N chr7 1871156 N DUP 5
A00404:155:HV27LDSXX:4:2640:12789:23797 chr7 1871243 N chr7 1871346 N DEL 5
A00404:156:HV37TDSXX:2:1368:6063:1407 chr7 1871319 N chr7 1871549 N DEL 2
A00297:158:HT275DSXX:3:1137:24722:14497 chr7 1870582 N chr7 1871345 N DUP 5
A00297:158:HT275DSXX:4:1154:6623:12587 chr7 1870582 N chr7 1871345 N DUP 5
A00404:156:HV37TDSXX:3:1241:1949:35806 chr7 1871287 N chr7 1871642 N DUP 5
A00297:158:HT275DSXX:2:2302:4490:7106 chr7 1870775 N chr7 1871388 N DEL 15
A00404:155:HV27LDSXX:3:2163:21911:23657 chr7 1870775 N chr7 1871388 N DEL 10
A00297:158:HT275DSXX:4:2313:10764:15655 chr7 1870623 N chr7 1871388 N DEL 5
A00404:156:HV37TDSXX:4:2218:11288:24424 chr7 1870419 N chr7 1871388 N DEL 5
A00404:155:HV27LDSXX:4:1623:30662:13354 chr7 1870577 N chr7 1871393 N DEL 5
A00297:158:HT275DSXX:4:1642:8721:32972 chr7 1870419 N chr7 1871388 N DEL 5
A00404:155:HV27LDSXX:4:1623:30662:13354 chr7 1870368 N chr7 1871388 N DEL 5
A00297:158:HT275DSXX:3:2659:23628:2832 chr7 1870371 N chr7 1871391 N DEL 5
A00297:158:HT275DSXX:2:1148:31503:36511 chr7 1871473 N chr7 1871574 N DUP 20
A00297:158:HT275DSXX:2:1148:31503:36511 chr7 1871346 N chr7 1871625 N DUP 20
A00404:156:HV37TDSXX:3:1247:17996:8860 chr7 1871541 N chr7 1871820 N DEL 21
A00297:158:HT275DSXX:3:1415:30671:19445 chr7 1870635 N chr7 1871730 N DEL 19
A00404:156:HV37TDSXX:1:1624:27986:6621 chr7 1871575 N chr7 1871650 N DUP 7
A00297:158:HT275DSXX:4:2268:28800:34992 chr7 1870406 N chr7 1871680 N DEL 5
A00404:155:HV27LDSXX:1:1262:20754:31422 chr7 1870748 N chr7 1871868 N DEL 23
A00404:155:HV27LDSXX:3:1411:21811:30624 chr7 1871254 N chr7 1871890 N DEL 5
A00404:156:HV37TDSXX:4:1464:18674:16110 chr7 1871638 N chr7 1871892 N DEL 5
A00404:155:HV27LDSXX:4:2463:22742:28322 chr20 34659291 N chr20 34659515 N DUP 5
A00404:156:HV37TDSXX:1:1429:27525:36730 chr20 34659292 N chr20 34659516 N DUP 5
A00404:156:HV37TDSXX:3:2531:6343:20055 chr20 34659305 N chr20 34659529 N DUP 1
A00297:158:HT275DSXX:2:1647:8612:25739 chr20 34659395 N chr20 34659570 N DUP 3
A00297:158:HT275DSXX:1:1639:6424:21919 chr20 34659291 N chr20 34659515 N DUP 3
A00404:155:HV27LDSXX:2:1127:32759:16016 chr20 34659334 N chr20 34659433 N DEL 5
A00297:158:HT275DSXX:2:1320:18593:20196 chr20 34659339 N chr20 34659438 N DEL 5
A00404:156:HV37TDSXX:3:2448:18855:11350 chr20 34659345 N chr20 34659569 N DUP 2
A00404:155:HV27LDSXX:4:2225:2094:24189 chr20 34659425 N chr20 34659551 N DUP 4
A00297:158:HT275DSXX:2:1657:27606:24502 chr20 34659444 N chr20 34659570 N DUP 10
A00297:158:HT275DSXX:1:1458:8115:34804 chr20 34659374 N chr20 34659600 N DEL 5
A00404:156:HV37TDSXX:4:1351:30282:33458 chr20 34659382 N chr20 34659608 N DEL 1
A00404:156:HV37TDSXX:2:1232:21920:1188 chr11 47562389 N chr11 47562692 N DEL 2
A00404:155:HV27LDSXX:2:1369:4743:25207 chr9 136294059 N chr9 136294142 N DUP 2
A00297:158:HT275DSXX:1:2340:23348:19225 chr9 136294140 N chr9 136294267 N DUP 7
A00297:158:HT275DSXX:1:1571:20582:3192 chr9 136294148 N chr9 136294273 N DUP 10
A00404:155:HV27LDSXX:2:1155:17363:6073 chr9 136294140 N chr9 136294267 N DUP 9
A00297:158:HT275DSXX:2:1423:7735:26663 chr9 136294140 N chr9 136294267 N DUP 9
A00404:156:HV37TDSXX:1:2377:29767:28056 chr10 126143285 N chr10 126143392 N DUP 3
A00404:156:HV37TDSXX:4:1260:26440:5509 chr10 126143312 N chr10 126143403 N DUP 5
A00297:158:HT275DSXX:4:2639:13431:17989 chr10 126143253 N chr10 126143489 N DUP 5
A00404:156:HV37TDSXX:3:2473:26359:15170 chr6 169937320 N chr6 169937374 N DUP 3
A00404:156:HV37TDSXX:4:1537:4580:18286 chr6 169937308 N chr6 169937362 N DUP 5
A00404:156:HV37TDSXX:4:2235:20961:16313 chr6 169937308 N chr6 169937362 N DUP 5
A00404:156:HV37TDSXX:3:2127:19253:31516 chr6 169937308 N chr6 169937362 N DUP 8
A00297:158:HT275DSXX:2:1431:3405:36072 chr6 169937308 N chr6 169937362 N DUP 10
A00404:155:HV27LDSXX:1:1533:30825:36432 chr6 169937308 N chr6 169937362 N DUP 13
A00404:156:HV37TDSXX:1:1541:24117:23062 chr6 169937313 N chr6 169937369 N DEL 9
A00404:156:HV37TDSXX:2:1548:17960:19319 chr21 46068961 N chr21 46069018 N DEL 12
A00404:156:HV37TDSXX:4:1556:20880:36495 chr19 11276793 N chr19 11277223 N DUP 5
A00297:158:HT275DSXX:4:2542:18439:11381 chr19 11276817 N chr19 11277133 N DEL 11
A00404:155:HV27LDSXX:4:2177:13340:33332 chr19 11276898 N chr19 11277169 N DEL 19
A00404:155:HV27LDSXX:2:2337:31828:11146 chr19 11276965 N chr19 11277238 N DEL 5
A00404:155:HV27LDSXX:1:1272:25048:12587 chr19 11276807 N chr19 11277239 N DEL 5
A00404:155:HV27LDSXX:1:1272:25491:23093 chr19 11276807 N chr19 11277239 N DEL 5
A00404:155:HV27LDSXX:1:1272:25997:12477 chr19 11276807 N chr19 11277239 N DEL 5
A00297:158:HT275DSXX:4:1512:30228:11005 chr19 11276808 N chr19 11277240 N DEL 5
A00404:156:HV37TDSXX:4:2634:6741:23750 chrX 2137256 N chrX 2137389 N DEL 11
A00297:158:HT275DSXX:3:2111:5918:20071 chrX 2137256 N chrX 2137389 N DEL 6
A00404:156:HV37TDSXX:1:2251:15130:26349 chrX 2137149 N chrX 2137298 N DUP 5
A00404:156:HV37TDSXX:1:2322:23755:20525 chrX 2137149 N chrX 2137298 N DUP 5
A00404:156:HV37TDSXX:4:1606:12545:3646 chrX 2137313 N chrX 2137380 N DEL 21
A00404:156:HV37TDSXX:1:2322:23755:20525 chrX 2137275 N chrX 2137349 N DUP 34
A00297:158:HT275DSXX:2:2453:31494:10880 chr7 151948184 N chr7 151948286 N DUP 6
A00297:158:HT275DSXX:2:2453:32208:12054 chr7 151948184 N chr7 151948286 N DUP 6
A00404:156:HV37TDSXX:1:2336:12427:4351 chr7 151948226 N chr7 151948318 N DUP 10
A00404:156:HV37TDSXX:2:1538:14362:26021 chr10 700383 N chr10 700479 N DEL 7
A00297:158:HT275DSXX:4:1521:3070:29512 chr7 128513771 N chr7 128513909 N DEL 5
A00404:155:HV27LDSXX:1:1138:16740:31015 chr4 1194959 N chr4 1195129 N DEL 41
A00404:155:HV27LDSXX:2:1215:18982:23563 chr4 1195027 N chr4 1195216 N DEL 15
A00297:158:HT275DSXX:4:1217:5439:2268 chr4 1195016 N chr4 1195140 N DUP 5
A00404:155:HV27LDSXX:3:2265:21368:31015 chr4 1195060 N chr4 1195142 N DUP 5
A00404:155:HV27LDSXX:4:2415:21052:12680 chr4 1195060 N chr4 1195142 N DUP 5
A00404:155:HV27LDSXX:3:2502:28031:26115 chr4 1195116 N chr4 1195198 N DUP 9
A00404:155:HV27LDSXX:1:1427:27588:23062 chr4 1195112 N chr4 1195194 N DUP 11
A00404:155:HV27LDSXX:2:2439:7265:5650 chr4 1195152 N chr4 1195216 N DEL 5
A00404:156:HV37TDSXX:4:1526:7853:11209 chr4 1195152 N chr4 1195216 N DEL 5
A00297:158:HT275DSXX:1:2534:8024:32643 chr4 1195112 N chr4 1195194 N DUP 10
A00297:158:HT275DSXX:4:1540:32705:36495 chr4 1195112 N chr4 1195194 N DUP 12
A00404:156:HV37TDSXX:2:2447:20130:22232 chr4 1195112 N chr4 1195194 N DUP 34
A00297:158:HT275DSXX:3:2206:5936:35540 chr4 1194996 N chr4 1195187 N DEL 3
A00404:156:HV37TDSXX:1:2513:17427:13917 chr4 1195096 N chr4 1195222 N DEL 5
A00404:155:HV27LDSXX:1:2416:15338:2722 chr4 1195075 N chr4 1195222 N DEL 5
A00404:155:HV27LDSXX:4:1460:18548:2707 chr4 1195069 N chr4 1195216 N DEL 5
A00404:156:HV37TDSXX:3:1475:30327:13996 chr16 34014831 N chr16 34014900 N DUP 5
A00297:158:HT275DSXX:3:2329:30165:33818 chr16 57705696 N chr16 57706709 N DUP 3
A00404:156:HV37TDSXX:2:2520:14705:14465 chr16 57705525 N chr16 57705935 N DEL 3
A00404:155:HV27LDSXX:3:2234:17544:1157 chr16 57705518 N chr16 57705928 N DEL 10
A00297:158:HT275DSXX:1:2166:16197:30890 chr16 57706129 N chr16 57706355 N DUP 5
A00297:158:HT275DSXX:1:2445:22010:20040 chr16 57705697 N chr16 57706314 N DEL 5
A00404:155:HV27LDSXX:3:1476:4047:31297 chr16 57706338 N chr16 57707028 N DUP 3
A00297:158:HT275DSXX:3:2234:20726:18286 chr16 57706467 N chr16 57706826 N DEL 5
A00404:156:HV37TDSXX:2:2461:25482:16407 chr16 57706475 N chr16 57706834 N DEL 5
A00297:158:HT275DSXX:2:2170:18647:17221 chr16 57705814 N chr16 57706562 N DEL 3
A00297:158:HT275DSXX:4:1646:2609:3161 chr16 57706102 N chr16 57706671 N DEL 53
A00404:155:HV27LDSXX:4:2509:12861:24956 chr16 57706671 N chr16 57706948 N DUP 1
A00404:156:HV37TDSXX:3:2460:28501:15562 chr16 57706671 N chr16 57706980 N DUP 4
A00404:156:HV37TDSXX:3:2434:20518:27258 chr16 57705629 N chr16 57706874 N DEL 5
A00404:156:HV37TDSXX:3:2434:20518:27258 chr16 57705629 N chr16 57706874 N DEL 5
A00404:155:HV27LDSXX:4:2516:9869:20870 chr7 1481779 N chr7 1481888 N DEL 16
A00404:156:HV37TDSXX:1:2274:26259:28494 chr11 2291170 N chr11 2292466 N DEL 16
A00404:155:HV27LDSXX:1:2340:26015:12727 chr11 2291431 N chr11 2292513 N DEL 10
A00404:156:HV37TDSXX:3:1454:4544:15843 chr11 2291178 N chr11 2291398 N DEL 5
A00404:156:HV37TDSXX:2:1350:17101:28980 chr11 2291476 N chr11 2292778 N DUP 5
A00404:155:HV27LDSXX:2:1328:31358:28714 chr11 2291260 N chr11 2291534 N DEL 25
A00404:155:HV27LDSXX:3:1259:5339:7921 chr11 2291657 N chr11 2292739 N DUP 5
A00404:156:HV37TDSXX:4:2124:15004:6120 chr11 2291223 N chr11 2291658 N DEL 1
A00404:155:HV27LDSXX:2:1327:4734:9220 chr11 2291431 N chr11 2291708 N DEL 6
A00297:158:HT275DSXX:4:2220:19605:35540 chr11 2291750 N chr11 2291907 N DEL 10
A00404:155:HV27LDSXX:3:2675:8675:10692 chr11 2291461 N chr11 2292595 N DUP 10
A00404:156:HV37TDSXX:1:2646:7175:13542 chr11 2291523 N chr11 2292331 N DEL 5
A00404:155:HV27LDSXX:2:1328:31358:28714 chr11 2291260 N chr11 2291534 N DEL 19
A00297:158:HT275DSXX:2:1601:2537:29966 chr11 2291587 N chr11 2292285 N DEL 7
A00404:155:HV27LDSXX:1:1130:9679:18443 chr11 2291504 N chr11 2291615 N DEL 14
A00297:158:HT275DSXX:2:1167:9037:10942 chr11 2291425 N chr11 2292185 N DEL 7
A00297:158:HT275DSXX:2:1167:9037:10942 chr11 2291427 N chr11 2292187 N DEL 5
A00404:155:HV27LDSXX:1:1322:18032:34068 chr11 2291532 N chr11 2292233 N DEL 15
A00404:156:HV37TDSXX:4:1131:25762:11224 chr11 2291311 N chr11 2292666 N DEL 16
A00404:155:HV27LDSXX:2:2208:32099:25989 chr11 2291489 N chr11 2292297 N DEL 3
A00404:156:HV37TDSXX:1:2212:2853:30013 chr11 2292394 N chr11 2292727 N DEL 11
A00404:155:HV27LDSXX:2:2208:32099:25989 chr11 2292394 N chr11 2292615 N DEL 14
A00404:155:HV27LDSXX:3:2222:15275:17832 chr11 2292408 N chr11 2292571 N DUP 5
A00297:158:HT275DSXX:3:1264:21775:33035 chr11 2291494 N chr11 2291605 N DEL 8
A00404:156:HV37TDSXX:1:2212:2853:30013 chr11 2292394 N chr11 2292727 N DEL 13
A00297:158:HT275DSXX:3:1323:2139:10708 chr11 2291644 N chr11 2292558 N DUP 5
A00404:156:HV37TDSXX:1:2113:4969:6590 chr11 2291644 N chr11 2292558 N DUP 5
A00404:155:HV27LDSXX:2:1135:6126:27665 chr11 2291644 N chr11 2292558 N DUP 5
A00404:155:HV27LDSXX:3:2603:4146:17910 chr11 2291587 N chr11 2292503 N DEL 2
A00404:156:HV37TDSXX:1:2436:7491:25864 chr11 2291288 N chr11 2292533 N DEL 1
A00297:158:HT275DSXX:4:2659:6253:5901 chr11 2292509 N chr11 2292788 N DEL 22
A00404:155:HV27LDSXX:1:2148:26820:12430 chr11 2291214 N chr11 2292788 N DEL 5
A00404:155:HV27LDSXX:3:1149:9100:16532 chr11 2291207 N chr11 2292783 N DEL 12
A00297:158:HT275DSXX:3:1323:2139:10708 chr11 2291181 N chr11 2292811 N DEL 4
A00404:155:HV27LDSXX:2:2535:7084:24439 chr12 48842421 N chr12 48842599 N DEL 5
A00404:155:HV27LDSXX:2:1457:27552:9565 chr12 48842342 N chr12 48842516 N DUP 10
A00404:156:HV37TDSXX:4:2402:21838:13636 chr12 48842444 N chr12 48842571 N DUP 5
A00404:155:HV27LDSXX:1:1642:11659:16767 chr1 168472147 N chr1 168472320 N DEL 12
A00297:158:HT275DSXX:4:2447:2058:8907 chr1 168472161 N chr1 168472280 N DEL 15
A00297:158:HT275DSXX:3:1414:8929:24752 chr1 168472174 N chr1 168472253 N DUP 15
A00297:158:HT275DSXX:4:1130:3206:31563 chr1 168472137 N chr1 168472318 N DUP 17
A00404:156:HV37TDSXX:4:1138:10673:36166 chr1 168472246 N chr1 168472295 N DUP 7
A00404:155:HV27LDSXX:2:1134:24704:21010 chr1 168472246 N chr1 168472295 N DUP 2
A00404:156:HV37TDSXX:1:2125:4218:16000 chr1 168472203 N chr1 168472338 N DUP 13
A00404:156:HV37TDSXX:4:2550:22372:14873 chr1 168472146 N chr1 168472327 N DUP 8
A00404:156:HV37TDSXX:1:1304:18367:16047 chr1 168472125 N chr1 168472226 N DEL 11
A00404:156:HV37TDSXX:2:1445:28944:21590 chr1 168472119 N chr1 168472240 N DEL 1
A00404:155:HV27LDSXX:3:2406:23077:5353 chr1 168472118 N chr1 168472321 N DEL 7
A00404:156:HV37TDSXX:3:1233:22869:10410 chr1 168472244 N chr1 168472327 N DEL 4
A00404:156:HV37TDSXX:2:1466:1732:15577 chr1 168472129 N chr1 168472372 N DEL 3
A00404:156:HV37TDSXX:2:1466:2953:15248 chr1 168472129 N chr1 168472372 N DEL 3
A00404:155:HV27LDSXX:2:2169:18954:15405 chrX 940150 N chrX 940645 N DUP 7
A00404:155:HV27LDSXX:2:2117:15600:11068 chr20 62585206 N chr20 62585283 N DUP 4
A00404:155:HV27LDSXX:4:2172:6090:1642 chr20 62585300 N chr20 62585505 N DEL 5
A00404:155:HV27LDSXX:1:2622:4824:25755 chr20 62585223 N chr20 62585302 N DEL 5
A00404:155:HV27LDSXX:4:2426:16929:24549 chr20 62585223 N chr20 62585302 N DEL 5
A00297:158:HT275DSXX:1:1336:22155:6417 chr20 62585234 N chr20 62585313 N DEL 4
A00404:156:HV37TDSXX:2:2330:25247:19914 chr20 62585234 N chr20 62585313 N DEL 4
A00404:156:HV37TDSXX:4:2210:15483:11459 chr20 62585388 N chr20 62585573 N DUP 4
A00404:156:HV37TDSXX:1:2451:22525:34929 chr20 62585211 N chr20 62585410 N DEL 9
A00404:155:HV27LDSXX:4:1340:6090:4993 chr20 62585179 N chr20 62585430 N DEL 5
A00404:156:HV37TDSXX:4:2174:19253:4836 chr20 62585218 N chr20 62585439 N DEL 5
A00404:156:HV37TDSXX:1:1431:2627:18192 chr7 2388935 N chr7 2389187 N DEL 13
A00297:158:HT275DSXX:4:1369:21368:21840 chr7 2388946 N chr7 2389281 N DEL 6
A00404:156:HV37TDSXX:1:1259:23104:3709 chr7 2388935 N chr7 2389229 N DEL 2
A00404:156:HV37TDSXX:1:1259:23104:3709 chr7 2388935 N chr7 2389229 N DEL 11
A00404:156:HV37TDSXX:1:1431:2627:18192 chr7 2388935 N chr7 2389187 N DEL 32
A00297:158:HT275DSXX:3:2140:1886:2691 chr7 2388960 N chr7 2389081 N DUP 7
A00404:156:HV37TDSXX:3:2207:3360:28761 chr7 2389169 N chr7 2389420 N DEL 5
A00404:155:HV27LDSXX:1:1359:18656:10034 chr7 2389079 N chr7 2389292 N DEL 9
A00404:156:HV37TDSXX:3:1613:25880:1783 chr7 2389227 N chr7 2389478 N DEL 5
A00404:156:HV37TDSXX:3:1613:25880:1783 chr7 2389291 N chr7 2389542 N DEL 5
A00404:155:HV27LDSXX:4:2502:31530:22310 chr14 76734845 N chr14 76735198 N DEL 5
A00297:158:HT275DSXX:2:2320:12454:33301 chr14 76734865 N chr14 76735216 N DUP 5
A00297:158:HT275DSXX:1:2369:6903:8625 chr14 76734695 N chr14 76734866 N DEL 5
A00297:158:HT275DSXX:3:2234:25373:5916 chr14 76734868 N chr14 76735219 N DUP 5
A00404:156:HV37TDSXX:2:2370:20329:23703 chr14 76735080 N chr14 76735237 N DEL 35
A00297:158:HT275DSXX:2:1139:8965:1172 chr14 76734852 N chr14 76735205 N DEL 1
A00404:155:HV27LDSXX:4:2337:12825:17660 chr16 7229893 N chr16 7229948 N DEL 10
A00404:155:HV27LDSXX:1:1463:6533:17628 chr16 7229891 N chr16 7229964 N DEL 15
A00297:158:HT275DSXX:4:2264:4237:19914 chr16 7229893 N chr16 7229948 N DEL 15
A00404:155:HV27LDSXX:4:2550:2338:29371 chr16 7229912 N chr16 7230197 N DUP 22
A00297:158:HT275DSXX:3:1472:8024:32831 chr16 7229808 N chr16 7229934 N DEL 5
A00404:155:HV27LDSXX:1:1453:19108:26349 chr16 7229948 N chr16 7230179 N DUP 20
A00404:156:HV37TDSXX:2:1214:30373:4961 chr16 7229954 N chr16 7230185 N DUP 17
A00404:156:HV37TDSXX:4:1448:21477:7623 chr16 7230002 N chr16 7230179 N DUP 30
A00404:155:HV27LDSXX:2:1516:13901:18771 chr16 7230092 N chr16 7230197 N DUP 27
A00297:158:HT275DSXX:1:1667:29975:25911 chr16 7230092 N chr16 7230197 N DUP 30
A00404:156:HV37TDSXX:2:1301:14841:21746 chr16 7230092 N chr16 7230197 N DUP 30
A00297:158:HT275DSXX:1:1476:18882:11428 chr16 7229871 N chr16 7230056 N DEL 5
A00404:156:HV37TDSXX:2:2142:31901:14779 chr16 7229948 N chr16 7230179 N DUP 26
A00297:158:HT275DSXX:1:1670:20003:21731 chr16 7229859 N chr16 7230204 N DEL 14
A00404:156:HV37TDSXX:4:1344:11921:6292 chr16 7229799 N chr16 7230211 N DEL 5
A00297:158:HT275DSXX:1:2341:12210:17347 chr16 7229802 N chr16 7230214 N DEL 5
A00404:156:HV37TDSXX:2:1219:15121:25989 chr7 154779248 N chr7 154779352 N DUP 3
A00404:155:HV27LDSXX:1:1329:11369:33677 chr2 2185577 N chr2 2186280 N DEL 5
A00404:155:HV27LDSXX:2:2629:32551:19006 chr2 2185609 N chr2 2185808 N DEL 13
A00404:155:HV27LDSXX:1:1329:11369:33677 chr2 2185604 N chr2 2185803 N DEL 20
A00297:158:HT275DSXX:1:1201:20356:3176 chr2 2185623 N chr2 2185723 N DEL 8
A00297:158:HT275DSXX:1:2534:30129:19695 chr2 2185776 N chr2 2186182 N DEL 5
A00297:158:HT275DSXX:2:2126:20401:24831 chr2 2185723 N chr2 2185875 N DUP 5
A00404:155:HV27LDSXX:1:1521:15727:30076 chr2 2185839 N chr2 2186146 N DEL 5
A00297:158:HT275DSXX:1:1201:18728:14512 chr2 2185721 N chr2 2185821 N DEL 15
A00297:158:HT275DSXX:1:1201:20356:3176 chr2 2185637 N chr2 2185791 N DEL 5
A00404:155:HV27LDSXX:3:2605:16297:24455 chr2 2185874 N chr2 2186181 N DEL 5
A00404:155:HV27LDSXX:1:1521:15727:30076 chr2 2185839 N chr2 2186146 N DEL 15
A00404:156:HV37TDSXX:4:1446:22363:6245 chr2 2185741 N chr2 2185848 N DUP 5
A00404:155:HV27LDSXX:1:2242:11487:17284 chr2 2185990 N chr2 2186189 N DEL 12
A00297:158:HT275DSXX:3:1615:14407:4961 chr2 2185854 N chr2 2185963 N DEL 1
A00297:158:HT275DSXX:1:2624:19931:33567 chr2 2185710 N chr2 2186114 N DUP 2
A00297:158:HT275DSXX:3:1472:7907:3537 chr2 2185710 N chr2 2186114 N DUP 2
A00404:155:HV27LDSXX:3:1130:17309:27430 chr2 2185710 N chr2 2186114 N DUP 5
A00404:156:HV37TDSXX:2:2353:5159:32941 chr2 2185822 N chr2 2186129 N DEL 15
A00404:155:HV27LDSXX:1:2318:21287:10300 chr2 2185839 N chr2 2186146 N DEL 10
A00404:156:HV37TDSXX:1:2669:12102:9298 chr2 2185710 N chr2 2186114 N DUP 5
A00404:155:HV27LDSXX:2:2217:3694:13182 chr2 2185715 N chr2 2186119 N DUP 5
A00404:155:HV27LDSXX:4:1218:5819:7310 chr2 2186188 N chr2 2186288 N DEL 5
A00404:156:HV37TDSXX:1:1636:29830:22842 chr2 2185726 N chr2 2186132 N DEL 5
A00404:155:HV27LDSXX:2:2217:2899:14716 chr2 2186066 N chr2 2186166 N DEL 13
A00404:156:HV37TDSXX:2:2670:9019:36526 chr2 2186225 N chr2 2186379 N DEL 10
A00404:155:HV27LDSXX:3:2605:16297:24455 chr2 2185874 N chr2 2186181 N DEL 5
A00404:155:HV27LDSXX:1:2242:11487:17284 chr2 2185990 N chr2 2186189 N DEL 5
A00404:156:HV37TDSXX:2:1536:28673:6339 chr2 2186262 N chr2 2186362 N DEL 14
A00404:156:HV37TDSXX:3:2241:3034:21245 chr2 2185948 N chr2 2186244 N DUP 5
A00404:155:HV27LDSXX:3:1130:17309:27430 chr2 2185758 N chr2 2186263 N DEL 5
A00404:155:HV27LDSXX:2:2530:32145:8343 chr2 2185634 N chr2 2186292 N DEL 5
A00404:156:HV37TDSXX:1:1177:28094:1892 chr2 2186233 N chr2 2186333 N DEL 5
A00404:156:HV37TDSXX:2:2521:2889:11694 chr2 2186225 N chr2 2186325 N DEL 5
A00404:155:HV27LDSXX:2:1530:24379:13432 chr2 2185729 N chr2 2186387 N DEL 5
A00297:158:HT275DSXX:4:1109:28257:25379 chr2 2185745 N chr2 2186403 N DEL 1
A00297:158:HT275DSXX:1:2428:16025:32910 chr2 2185676 N chr2 2186433 N DEL 5
A00404:155:HV27LDSXX:4:1333:9959:16329 chr19 55266641 N chr19 55266803 N DEL 11
A00404:155:HV27LDSXX:1:1462:16016:12602 chr19 55266535 N chr19 55266645 N DUP 15
A00297:158:HT275DSXX:4:2378:31123:3818 chr19 55266535 N chr19 55266645 N DUP 28
A00404:156:HV37TDSXX:3:2418:8015:12211 chr19 55266535 N chr19 55266645 N DUP 28
A00404:156:HV37TDSXX:4:2609:16125:4554 chr19 55266535 N chr19 55266645 N DUP 19
A00404:155:HV27LDSXX:1:2348:4119:35274 chr19 55266609 N chr19 55266662 N DUP 7
A00297:158:HT275DSXX:4:1632:23945:27398 chr19 55266535 N chr19 55266645 N DUP 15
A00297:158:HT275DSXX:4:2632:18222:36119 chr19 55266535 N chr19 55266645 N DUP 15
A00404:155:HV27LDSXX:3:1232:17454:34945 chr19 55266634 N chr19 55266710 N DUP 27
A00297:158:HT275DSXX:4:1359:5466:22013 chr19 55266634 N chr19 55266710 N DUP 27
A00404:155:HV27LDSXX:4:1628:5782:16078 chr19 55266551 N chr19 55266627 N DEL 8
A00297:158:HT275DSXX:2:1332:31132:20901 chr19 55266637 N chr19 55266713 N DUP 10
A00404:155:HV27LDSXX:3:2339:18593:2910 chr19 55266704 N chr19 55266753 N DUP 16
A00297:158:HT275DSXX:1:2258:17969:8093 chr19 55266552 N chr19 55266646 N DEL 3
A00404:156:HV37TDSXX:3:1439:30933:21684 chr12 25199486 N chr12 25199546 N DEL 2
A00404:156:HV37TDSXX:3:1453:26838:18098 chr12 25199511 N chr12 25199570 N DUP 2
A00404:155:HV27LDSXX:2:1478:24080:20181 chr16 89017373 N chr16 89017673 N DEL 5
A00404:155:HV27LDSXX:3:1212:29568:2127 chr16 89017603 N chr16 89017674 N DEL 8
A00404:156:HV37TDSXX:2:1574:4463:23281 chr17 65500137 N chr17 65500242 N DUP 15
A00404:155:HV27LDSXX:4:1241:32913:3756 chr17 65500248 N chr17 65500383 N DEL 15
A00404:155:HV27LDSXX:4:2241:32407:1031 chr17 65500248 N chr17 65500383 N DEL 15
A00404:155:HV27LDSXX:1:1231:30318:34460 chr17 65500248 N chr17 65500383 N DEL 16
A00404:156:HV37TDSXX:3:2633:24297:14669 chr17 65500248 N chr17 65500383 N DEL 16
A00297:158:HT275DSXX:2:1470:2709:20776 chr17 65500105 N chr17 65500265 N DEL 2
A00404:155:HV27LDSXX:2:2534:1470:17816 chr17 65500123 N chr17 65500374 N DUP 12
A00404:155:HV27LDSXX:1:2311:5475:7842 chr17 65500109 N chr17 65500291 N DEL 5
A00297:158:HT275DSXX:2:2559:4490:6543 chr17 65500342 N chr17 65500415 N DEL 5
A00404:155:HV27LDSXX:4:2112:1344:11772 chr17 65500100 N chr17 65500540 N DEL 3
A00404:155:HV27LDSXX:3:1465:1814:12054 chr16 34658667 N chr16 34659356 N DEL 5
A00404:156:HV37TDSXX:4:2427:31539:6918 chr16 34659023 N chr16 34659168 N DEL 5
A00404:156:HV37TDSXX:3:2271:29649:10379 chr16 34658992 N chr16 34659578 N DEL 28
A00404:155:HV27LDSXX:2:1360:30553:26068 chr2 190365995 N chr2 190366440 N DEL 4
A00404:156:HV37TDSXX:2:2437:26295:34444 chr2 190366109 N chr2 190366736 N DEL 6
A00404:155:HV27LDSXX:4:2639:26458:31720 chr2 190366092 N chr2 190366183 N DEL 2
A00404:156:HV37TDSXX:2:1457:11921:34632 chr2 190366114 N chr2 190366717 N DEL 11
A00404:156:HV37TDSXX:2:2171:15302:34287 chr2 190365969 N chr2 190366174 N DEL 2
A00297:158:HT275DSXX:2:1116:14009:18928 chr2 190365993 N chr2 190366300 N DUP 1
A00404:155:HV27LDSXX:4:2249:2899:19820 chr2 190365993 N chr2 190366300 N DUP 2
A00297:158:HT275DSXX:1:1354:8865:12837 chr2 190366240 N chr2 190366765 N DUP 1
A00404:156:HV37TDSXX:3:1264:1886:29403 chr2 190366421 N chr2 190366732 N DEL 2
A00404:156:HV37TDSXX:3:1337:30020:32315 chr2 190366426 N chr2 190366735 N DEL 11
A00297:158:HT275DSXX:3:1416:10429:7091 chr2 190366289 N chr2 190366616 N DUP 2
A00297:158:HT275DSXX:4:1369:22724:19210 chr2 190366289 N chr2 190366616 N DUP 4
A00297:158:HT275DSXX:3:2243:15393:5885 chr2 190366026 N chr2 190366571 N DEL 13
A00404:156:HV37TDSXX:2:2672:28782:19711 chr2 190366290 N chr2 190366573 N DEL 11
A00297:158:HT275DSXX:2:2269:4933:26694 chr1 2348860 N chr1 2348951 N DEL 31
A00297:158:HT275DSXX:1:1218:27923:16720 chr1 2348877 N chr1 2348980 N DUP 23
A00297:158:HT275DSXX:4:1667:21305:29872 chr1 2348877 N chr1 2348980 N DUP 23
A00404:155:HV27LDSXX:2:2111:5990:1344 chr1 2348872 N chr1 2348975 N DUP 28
A00404:156:HV37TDSXX:3:1139:7600:20290 chr1 2348872 N chr1 2348975 N DUP 28
A00297:158:HT275DSXX:4:2270:1244:24189 chr1 2348817 N chr1 2348880 N DEL 5
A00404:155:HV27LDSXX:2:2612:20889:24205 chr1 2348818 N chr1 2348881 N DEL 4
A00404:156:HV37TDSXX:4:1317:31665:5353 chr5 181002525 N chr5 181002622 N DEL 8
A00404:156:HV37TDSXX:4:1153:5367:12790 chr5 181002529 N chr5 181002626 N DEL 10
A00297:158:HT275DSXX:2:1672:26720:31046 chr5 181002525 N chr5 181002624 N DEL 11
A00404:156:HV37TDSXX:1:1223:27263:27884 chr5 181002525 N chr5 181002622 N DEL 13
A00404:156:HV37TDSXX:2:1206:24921:34131 chr5 181002535 N chr5 181002624 N DUP 2
A00297:158:HT275DSXX:1:1219:32000:17989 chr9 40600971 N chr9 40601135 N DUP 9
A00404:155:HV27LDSXX:2:2370:3549:9925 chr11 2384573 N chr11 2384693 N DEL 5
A00297:158:HT275DSXX:4:2448:13847:11694 chr4 78623619 N chr4 78623676 N DUP 5
A00404:155:HV27LDSXX:1:1407:27986:8782 chr4 78623619 N chr4 78623676 N DUP 5
A00404:155:HV27LDSXX:1:1407:27995:8797 chr4 78623619 N chr4 78623676 N DUP 5
A00404:156:HV37TDSXX:2:2466:23927:17973 chr4 78623619 N chr4 78623676 N DUP 5
A00297:158:HT275DSXX:3:1316:31864:25958 chr4 78623619 N chr4 78623676 N DUP 5
A00404:155:HV27LDSXX:1:1542:8006:28322 chr4 78623619 N chr4 78623676 N DUP 5
A00404:155:HV27LDSXX:2:2676:26784:13088 chr4 78623619 N chr4 78623676 N DUP 5
A00404:156:HV37TDSXX:3:2371:20121:3364 chr4 78623619 N chr4 78623676 N DUP 5
A00404:156:HV37TDSXX:4:1225:32597:6621 chr4 78623619 N chr4 78623676 N DUP 5
A00404:156:HV37TDSXX:4:1225:32714:5760 chr4 78623619 N chr4 78623676 N DUP 5
A00404:155:HV27LDSXX:2:2507:26096:18662 chr8 1631062 N chr8 1631153 N DEL 5
A00404:156:HV37TDSXX:4:1138:30165:23954 chr10 113976807 N chr10 113976883 N DUP 2
A00404:156:HV37TDSXX:1:2638:18475:35274 chr19 20344154 N chr19 20344252 N DUP 3
A00297:158:HT275DSXX:2:1572:25192:16595 chr3 161369388 N chr3 161369461 N DEL 7
A00297:158:HT275DSXX:4:1115:7184:36918 chr3 161369410 N chr3 161369477 N DEL 2
A00404:156:HV37TDSXX:1:1647:1850:33442 chr13 26123040 N chr13 26123113 N DUP 10
A00404:156:HV37TDSXX:4:2535:16441:4382 chr10 3377298 N chr10 3377458 N DEL 5
A00404:156:HV37TDSXX:3:1340:16721:21245 chr7 154884642 N chr7 154884749 N DUP 2
A00404:155:HV27LDSXX:4:1102:8097:27164 chr4 1236669 N chr4 1236775 N DEL 2
A00297:158:HT275DSXX:3:1638:5141:20885 chr4 1236709 N chr4 1237060 N DEL 10
A00404:156:HV37TDSXX:4:1370:26512:21230 chr4 1236744 N chr4 1236850 N DEL 15
A00297:158:HT275DSXX:3:2432:24930:15953 chr4 1236744 N chr4 1236850 N DEL 15
A00404:155:HV27LDSXX:2:1601:4327:22106 chr4 1236781 N chr4 1236852 N DEL 5
A00404:155:HV27LDSXX:1:2651:5294:16955 chr4 1236783 N chr4 1236854 N DEL 5
A00297:158:HT275DSXX:2:1615:12192:35289 chr4 1236786 N chr4 1236857 N DEL 8
A00297:158:HT275DSXX:1:1638:5927:24095 chr4 1236763 N chr4 1236869 N DEL 4
A00297:158:HT275DSXX:1:2303:25030:20259 chr4 1236705 N chr4 1236881 N DEL 5
A00297:158:HT275DSXX:2:2247:27299:23281 chr4 1236717 N chr4 1236928 N DEL 10
A00404:156:HV37TDSXX:4:1370:26512:21230 chr4 1236705 N chr4 1236881 N DEL 5
A00297:158:HT275DSXX:1:1638:5927:24095 chr4 1236845 N chr4 1237054 N DUP 13
A00297:158:HT275DSXX:1:1130:25319:10113 chr4 1237066 N chr4 1237207 N DEL 32
A00404:155:HV27LDSXX:3:2251:12924:3020 chr4 1236827 N chr4 1237038 N DEL 13
A00297:158:HT275DSXX:3:1615:11062:7373 chr4 1236677 N chr4 1237098 N DEL 7
A00404:155:HV27LDSXX:1:2310:28574:28933 chr13 98663758 N chr13 98663822 N DEL 15
A00404:155:HV27LDSXX:2:1412:31485:14873 chr6 29719445 N chr6 29719746 N DUP 7
A00404:155:HV27LDSXX:4:2465:1796:13088 chr6 29719356 N chr6 29719481 N DUP 1
A00404:156:HV37TDSXX:4:1561:10357:11256 chr6 29719396 N chr6 29719476 N DUP 2
A00404:156:HV37TDSXX:4:1352:14687:4163 chr6 29719400 N chr6 29719829 N DEL 7
A00297:158:HT275DSXX:2:2660:13693:22514 chr11 116347377 N chr11 116347634 N DEL 24
A00297:158:HT275DSXX:3:1176:15528:6026 chr11 116347242 N chr11 116347442 N DUP 5
A00404:156:HV37TDSXX:2:2322:24894:27665 chr11 116347359 N chr11 116347440 N DEL 2
A00404:155:HV27LDSXX:4:2370:25220:19241 chr11 116347257 N chr11 116347459 N DEL 5
A00404:156:HV37TDSXX:4:2352:9742:13291 chr11 116347509 N chr11 116347601 N DUP 5
A00404:156:HV37TDSXX:4:2235:15447:7513 chr11 116347523 N chr11 116347617 N DEL 5
A00404:155:HV27LDSXX:1:2239:24695:18584 chr1 230038373 N chr1 230038504 N DUP 5
A00404:156:HV37TDSXX:2:2320:3595:35806 chr1 230038393 N chr1 230038510 N DEL 10
A00404:155:HV27LDSXX:4:1325:9598:16736 chr1 230038391 N chr1 230038512 N DEL 8
A00404:155:HV27LDSXX:1:2206:19831:8281 chr1 230038390 N chr1 230038519 N DEL 1
A00297:158:HT275DSXX:3:2109:25916:21543 chr2 6253357 N chr2 6253547 N DEL 24
A00297:158:HT275DSXX:3:1622:20112:10488 chr2 6253437 N chr2 6253596 N DEL 15
A00404:155:HV27LDSXX:4:2671:26738:29982 chr2 6253422 N chr2 6253677 N DEL 30
A00404:156:HV37TDSXX:3:2547:3586:12649 chr2 6253475 N chr2 6253664 N DEL 24
A00404:155:HV27LDSXX:3:1112:22028:25363 chr2 6253475 N chr2 6253664 N DEL 43
A00297:158:HT275DSXX:1:2653:18114:26193 chr2 6253475 N chr2 6253664 N DEL 42
A00404:156:HV37TDSXX:4:1460:1127:22733 chr2 6253475 N chr2 6253664 N DEL 36
A00404:155:HV27LDSXX:1:1339:10239:5071 chr2 6253475 N chr2 6253664 N DEL 33
A00297:158:HT275DSXX:2:2357:4164:15718 chr2 6253422 N chr2 6253677 N DEL 14
A00404:156:HV37TDSXX:2:1407:13268:12383 chr2 6253491 N chr2 6253666 N DEL 18
A00404:155:HV27LDSXX:3:2465:5412:7012 chr2 6253491 N chr2 6253666 N DEL 11
A00404:155:HV27LDSXX:3:2307:9489:2018 chr5 41312751 N chr5 41312846 N DEL 4
A00404:155:HV27LDSXX:1:1123:32940:14450 chr5 41312751 N chr5 41312846 N DEL 4
A00404:155:HV27LDSXX:3:2212:20916:15358 chr5 41312752 N chr5 41312847 N DEL 3
A00404:155:HV27LDSXX:3:2347:3577:7999 chr5 41312752 N chr5 41312847 N DEL 3
A00404:155:HV27LDSXX:4:2469:28917:24893 chr5 41312752 N chr5 41312847 N DEL 3
A00404:155:HV27LDSXX:3:1446:1298:34147 chr5 41312786 N chr5 41312889 N DEL 2
A00404:156:HV37TDSXX:3:1452:17002:5040 chr13 60978170 N chr13 60978235 N DEL 10
A00404:155:HV27LDSXX:1:2245:23448:22748 chr13 60978236 N chr13 60978315 N DEL 20
A00404:155:HV27LDSXX:2:2365:7808:27821 chr13 60978236 N chr13 60978315 N DEL 19
A00404:156:HV37TDSXX:2:1207:18792:29747 chr13 60978236 N chr13 60978315 N DEL 19
A00404:156:HV37TDSXX:2:1521:22661:15593 chr9 15455980 N chr9 15456157 N DEL 5
A00404:155:HV27LDSXX:3:1529:17400:6449 chr9 15455981 N chr9 15456158 N DEL 4
A00297:158:HT275DSXX:3:1153:17273:7482 chr19 2377686 N chr19 2377739 N DUP 10
A00404:155:HV27LDSXX:3:2463:9769:28776 chr18 13823314 N chr18 13823430 N DEL 17
A00404:156:HV37TDSXX:3:2577:10999:4319 chr18 13823173 N chr18 13823338 N DUP 1
A00297:158:HT275DSXX:2:2341:31485:28213 chr18 13823179 N chr18 13823336 N DUP 17
A00404:156:HV37TDSXX:1:1634:8395:26772 chr18 13823131 N chr18 13823294 N DEL 5
A00297:158:HT275DSXX:4:2164:8097:21277 chr18 13823131 N chr18 13823294 N DEL 5
A00404:155:HV27LDSXX:4:1415:31006:35023 chr18 13823131 N chr18 13823294 N DEL 5
A00404:155:HV27LDSXX:2:2340:31268:31594 chr18 13823131 N chr18 13823294 N DEL 5
A00297:158:HT275DSXX:2:2341:31485:28213 chr18 13823179 N chr18 13823294 N DEL 10
A00404:155:HV27LDSXX:2:1142:19009:14622 chr18 13823179 N chr18 13823294 N DEL 7
A00297:158:HT275DSXX:1:2434:23773:26944 chr18 13823179 N chr18 13823294 N DEL 6
A00404:155:HV27LDSXX:1:1403:20220:26115 chr18 13823179 N chr18 13823294 N DEL 6
A00404:155:HV27LDSXX:1:1403:21929:25786 chr18 13823179 N chr18 13823294 N DEL 6
A00297:158:HT275DSXX:4:2153:5737:36824 chr18 13823239 N chr18 13823406 N DUP 1
A00297:158:HT275DSXX:3:2278:18792:8954 chr18 13823303 N chr18 13823418 N DUP 5
A00404:156:HV37TDSXX:2:1234:30816:20697 chr18 13823099 N chr18 13823428 N DUP 5
A00297:158:HT275DSXX:2:1371:1289:14904 chr18 13823237 N chr18 13823404 N DUP 4
A00404:156:HV37TDSXX:1:2576:26151:30373 chr18 13823099 N chr18 13823428 N DUP 5
A00404:155:HV27LDSXX:2:1625:12337:11772 chr18 13823373 N chr18 13823428 N DUP 5
A00297:158:HT275DSXX:2:1444:24343:19507 chr18 13823373 N chr18 13823428 N DUP 5
A00297:158:HT275DSXX:2:1671:7654:3975 chr18 13823318 N chr18 13823482 N DEL 18
A00404:155:HV27LDSXX:4:1204:20048:2362 chr18 13823318 N chr18 13823482 N DEL 28
A00297:158:HT275DSXX:2:1303:11116:8531 chr18 13823214 N chr18 13823488 N DEL 11
A00404:155:HV27LDSXX:3:2553:10474:33974 chr18 13823209 N chr18 13823483 N DEL 16
A00297:158:HT275DSXX:2:1371:1289:14904 chr18 13823266 N chr18 13823482 N DEL 17
A00404:155:HV27LDSXX:1:1221:12156:7357 chr18 13823112 N chr18 13823490 N DEL 7
A00404:156:HV37TDSXX:2:1361:6641:36636 chr4 140810967 N chr4 140811064 N DEL 17
A00297:158:HT275DSXX:4:2128:19000:23500 chr1 24800093 N chr1 24800219 N DUP 5
A00404:155:HV27LDSXX:2:1443:15564:32330 chr1 24800212 N chr1 24800509 N DUP 5
A00404:155:HV27LDSXX:2:2363:22589:36761 chr1 24800206 N chr1 24800603 N DEL 5
A00404:156:HV37TDSXX:4:2105:16206:14967 chr1 24800232 N chr1 24800629 N DEL 10
A00297:158:HT275DSXX:1:1623:27832:29622 chr1 24799946 N chr1 24800641 N DEL 3
A00404:156:HV37TDSXX:4:2105:16206:14967 chr1 24799946 N chr1 24800641 N DEL 3
A00297:158:HT275DSXX:3:2518:28854:18646 chr2 32293869 N chr2 32293993 N DEL 5
A00297:158:HT275DSXX:1:1129:7211:29700 chr16 4479876 N chr16 4480193 N DUP 3
A00404:156:HV37TDSXX:1:1615:17345:23923 chr16 4479891 N chr16 4480496 N DUP 2
A00404:155:HV27LDSXX:1:1468:19696:33160 chr16 4480066 N chr16 4480982 N DEL 3
A00404:155:HV27LDSXX:1:1570:21947:6809 chr19 49427826 N chr19 49427899 N DUP 7
A00297:158:HT275DSXX:1:1230:26133:16658 chr19 49427796 N chr19 49427869 N DUP 13
A00297:158:HT275DSXX:2:1428:26576:4241 chr10 132362756 N chr10 132363076 N DEL 5
A00297:158:HT275DSXX:3:1202:21983:13823 chr10 132362756 N chr10 132363193 N DEL 10
A00297:158:HT275DSXX:2:1428:26576:4241 chr10 132362756 N chr10 132363076 N DEL 15
A00404:155:HV27LDSXX:4:2534:26033:32988 chr10 132362768 N chr10 132362850 N DEL 4
A00404:156:HV37TDSXX:4:2238:15944:22686 chr10 132362768 N chr10 132362850 N DEL 10
A00404:155:HV27LDSXX:2:2668:1533:24972 chr10 132362781 N chr10 132363257 N DEL 16
A00404:155:HV27LDSXX:3:2116:28827:34068 chr10 132362780 N chr10 132362862 N DEL 3
A00404:155:HV27LDSXX:1:1649:25138:36198 chr10 132362781 N chr10 132362863 N DEL 2
A00297:158:HT275DSXX:1:2232:3577:25222 chr10 132362773 N chr10 132362855 N DEL 10
A00404:155:HV27LDSXX:1:1225:26395:33364 chr10 132362771 N chr10 132362853 N DEL 12
A00404:156:HV37TDSXX:1:2408:13666:33833 chr10 132362802 N chr10 132363122 N DEL 3
A00297:158:HT275DSXX:4:1302:27416:13025 chr10 132363062 N chr10 132363178 N DUP 2
A00297:158:HT275DSXX:1:1640:4327:28620 chr10 132362774 N chr10 132363250 N DEL 2
A00404:155:HV27LDSXX:4:2528:1181:6543 chr10 132362820 N chr10 132363377 N DEL 25
A00404:156:HV37TDSXX:2:2507:17309:36354 chr3 130868397 N chr3 130868618 N DEL 13
A00297:158:HT275DSXX:4:2456:5493:13510 chr3 130868416 N chr3 130868544 N DEL 10
A00404:155:HV27LDSXX:1:1229:18701:32722 chr3 130868387 N chr3 130868688 N DUP 5
A00404:155:HV27LDSXX:3:2531:26051:15890 chr3 130868458 N chr3 130868632 N DUP 15
A00404:155:HV27LDSXX:4:1363:3613:15608 chr3 130868658 N chr3 130868784 N DEL 5
A00404:156:HV37TDSXX:3:1139:9173:9424 chr3 130868299 N chr3 130868601 N DEL 5
A00404:156:HV37TDSXX:2:1239:5737:8202 chr3 130868357 N chr3 130868659 N DEL 5
A00404:155:HV27LDSXX:4:2219:13205:24330 chr3 130868434 N chr3 130868736 N DEL 10
A00297:158:HT275DSXX:1:1149:9191:34444 chr3 130868364 N chr3 130868840 N DUP 4
A00297:158:HT275DSXX:3:1353:7491:28213 chr3 130868341 N chr3 130868769 N DEL 5
A00404:155:HV27LDSXX:2:1347:29993:30326 chr7 10162992 N chr7 10163053 N DUP 13
A00404:156:HV37TDSXX:4:1462:19750:1094 chr7 10162992 N chr7 10163053 N DUP 14
A00404:156:HV37TDSXX:1:2241:14362:6167 chr7 10162992 N chr7 10163053 N DUP 14
A00404:156:HV37TDSXX:1:2171:3179:14293 chr7 10162992 N chr7 10163205 N DUP 8
A00297:158:HT275DSXX:1:2204:2835:31610 chr7 10162992 N chr7 10163053 N DUP 7
A00297:158:HT275DSXX:4:1125:25446:18724 chr7 10163032 N chr7 10163093 N DEL 8
A00404:155:HV27LDSXX:2:2432:7292:27242 chr7 10162992 N chr7 10163053 N DUP 7
A00404:155:HV27LDSXX:3:2411:31105:35884 chr7 10162992 N chr7 10163205 N DUP 12
A00404:155:HV27LDSXX:1:2167:10791:35963 chr7 10163032 N chr7 10163093 N DEL 7
A00404:156:HV37TDSXX:4:2403:2772:12524 chr7 10163040 N chr7 10163101 N DEL 7
A00297:158:HT275DSXX:4:2306:23357:7435 chr7 10163031 N chr7 10163124 N DEL 6
A00297:158:HT275DSXX:2:1614:27941:24392 chr7 10163031 N chr7 10163124 N DEL 6
A00404:156:HV37TDSXX:3:2550:7310:30467 chr7 10163031 N chr7 10163124 N DEL 6
A00404:156:HV37TDSXX:3:2550:7636:30373 chr7 10163031 N chr7 10163124 N DEL 6
A00404:155:HV27LDSXX:3:1651:12138:13338 chr7 10163032 N chr7 10163154 N DEL 7
A00404:156:HV37TDSXX:1:2537:24795:18912 chr7 10163032 N chr7 10163154 N DEL 7
A00404:155:HV27LDSXX:1:1128:14443:5901 chr7 10163032 N chr7 10163154 N DEL 7
A00404:155:HV27LDSXX:1:1128:14461:5901 chr7 10163032 N chr7 10163154 N DEL 7
A00297:158:HT275DSXX:1:1474:15863:30749 chr7 10163032 N chr7 10163154 N DEL 7
A00297:158:HT275DSXX:1:1474:17038:11866 chr7 10163032 N chr7 10163154 N DEL 7
A00297:158:HT275DSXX:1:1509:26069:4085 chr7 10163032 N chr7 10163154 N DEL 7
A00297:158:HT275DSXX:1:2319:21884:31250 chr7 10163032 N chr7 10163154 N DEL 7
A00404:156:HV37TDSXX:1:1229:11469:9862 chr7 10163032 N chr7 10163154 N DEL 7
A00404:156:HV37TDSXX:1:2312:13367:3787 chr7 10163032 N chr7 10163154 N DEL 7
A00404:156:HV37TDSXX:2:1521:13792:7028 chr7 10163032 N chr7 10163154 N DEL 7
A00297:158:HT275DSXX:1:1116:10203:7733 chr7 10163032 N chr7 10163154 N DEL 7
A00404:156:HV37TDSXX:2:2443:17644:36871 chr7 10163032 N chr7 10163154 N DEL 7
A00297:158:HT275DSXX:1:2608:2908:6057 chr7 10163035 N chr7 10163157 N DEL 7
A00297:158:HT275DSXX:4:1435:27805:13228 chr7 10163015 N chr7 10163168 N DEL 1
A00404:155:HV27LDSXX:4:2349:26639:4163 chr7 10163014 N chr7 10163167 N DEL 2
A00404:156:HV37TDSXX:1:2322:12102:27148 chr1 13101560 N chr1 13101638 N DEL 6
A00297:158:HT275DSXX:3:1673:14091:23578 chr8 1344232 N chr8 1344287 N DEL 13
A00297:158:HT275DSXX:3:1216:32063:15186 chr8 1344233 N chr8 1344286 N DUP 5
A00404:156:HV37TDSXX:3:1572:11668:11271 chr8 1344233 N chr8 1344286 N DUP 5
A00297:158:HT275DSXX:1:1653:18430:12336 chr8 1344233 N chr8 1344286 N DUP 5
A00404:156:HV37TDSXX:1:1259:4209:26130 chr8 1344233 N chr8 1344286 N DUP 5
A00297:158:HT275DSXX:1:1330:24722:15342 chr8 1344233 N chr8 1344286 N DUP 12
A00404:156:HV37TDSXX:3:2240:8856:18740 chr8 1344233 N chr8 1344286 N DUP 13
A00404:156:HV37TDSXX:2:1502:26250:32017 chr8 1344240 N chr8 1344293 N DUP 8
A00404:156:HV37TDSXX:3:2669:8784:23281 chr8 1344240 N chr8 1344293 N DUP 8
A00404:156:HV37TDSXX:4:1431:24768:19335 chr8 1344239 N chr8 1344292 N DUP 9
A00404:156:HV37TDSXX:1:1165:14253:7576 chr8 1344264 N chr8 1344317 N DUP 5
A00404:155:HV27LDSXX:2:1535:5638:14888 chr8 1344271 N chr8 1344353 N DEL 5
A00404:155:HV27LDSXX:2:1535:5791:14747 chr8 1344271 N chr8 1344353 N DEL 5
A00297:158:HT275DSXX:4:2101:29812:19398 chr8 1344271 N chr8 1344353 N DEL 5
A00297:158:HT275DSXX:4:2101:29857:18850 chr8 1344271 N chr8 1344353 N DEL 5
A00297:158:HT275DSXX:4:2253:12689:21903 chr8 1344271 N chr8 1344353 N DEL 9
A00297:158:HT275DSXX:4:2253:12798:21872 chr8 1344271 N chr8 1344353 N DEL 9
A00297:158:HT275DSXX:1:1530:19651:18928 chr12 131779363 N chr12 131779418 N DUP 5
A00297:158:HT275DSXX:1:2265:22227:30154 chr12 131779366 N chr12 131779449 N DUP 10
A00297:158:HT275DSXX:2:2153:22390:23140 chr12 131779363 N chr12 131779418 N DUP 16
A00297:158:HT275DSXX:3:2642:14959:29653 chr12 131779346 N chr12 131779429 N DUP 26
A00297:158:HT275DSXX:2:1132:9724:19774 chr12 131779366 N chr12 131779449 N DUP 10
A00297:158:HT275DSXX:1:2501:25156:22263 chr12 131779346 N chr12 131779429 N DUP 26
A00404:156:HV37TDSXX:1:2476:10465:19210 chr12 131779363 N chr12 131779418 N DUP 17
A00297:158:HT275DSXX:2:2108:28022:19429 chr12 131779346 N chr12 131779429 N DUP 27
A00297:158:HT275DSXX:4:2352:24071:31908 chr12 131779363 N chr12 131779418 N DUP 33
A00404:156:HV37TDSXX:2:1619:10474:2378 chr12 131779323 N chr12 131779406 N DUP 23
A00297:158:HT275DSXX:1:2265:22227:30154 chr12 131779346 N chr12 131779401 N DUP 8
A00404:155:HV27LDSXX:2:1468:28456:15107 chr4 57173566 N chr4 57173617 N DEL 6
A00404:156:HV37TDSXX:2:2552:17924:31657 chr1 156170505 N chr1 156170796 N DEL 6
A00404:156:HV37TDSXX:2:2552:17924:31657 chr1 156170514 N chr1 156170805 N DEL 8
A00297:158:HT275DSXX:1:1627:31494:36338 chr2 113821627 N chr2 113821711 N DEL 18
A00297:158:HT275DSXX:1:1628:30382:16814 chr2 113821627 N chr2 113821711 N DEL 18
A00404:155:HV27LDSXX:1:2263:3947:33066 chr2 113821627 N chr2 113821711 N DEL 27
A00404:156:HV37TDSXX:2:1131:28067:31281 chr12 129549298 N chr12 129549561 N DEL 22
A00404:155:HV27LDSXX:3:2446:11984:27696 chr12 129549315 N chr12 129549579 N DEL 5
A00404:155:HV27LDSXX:3:2234:11089:19914 chr12 129549206 N chr12 129549470 N DEL 5
A00297:158:HT275DSXX:2:1505:18141:35352 chr12 129549248 N chr12 129549512 N DEL 5
A00404:155:HV27LDSXX:3:1166:16486:29042 chr12 129549315 N chr12 129549579 N DEL 15
A00404:155:HV27LDSXX:1:2376:15899:16971 chr5 137557089 N chr5 137557400 N DEL 3
A00404:156:HV37TDSXX:4:1303:5638:11819 chr5 137557089 N chr5 137557400 N DEL 3
A00404:156:HV37TDSXX:2:2278:10212:30044 chr5 137557089 N chr5 137557400 N DEL 4
A00404:156:HV37TDSXX:4:1276:5466:23703 chr4 52736361 N chr4 52736430 N DUP 2
A00404:156:HV37TDSXX:4:1617:29324:27915 chr4 52736380 N chr4 52736451 N DEL 5
A00404:156:HV37TDSXX:4:1617:29821:28056 chr4 52736380 N chr4 52736451 N DEL 5
A00404:156:HV37TDSXX:3:2533:22272:36965 chr8 141620188 N chr8 141620642 N DEL 1
A00404:155:HV27LDSXX:1:1507:31168:20838 chr8 141620235 N chr8 141620327 N DEL 10
A00404:156:HV37TDSXX:1:1330:5457:7247 chr8 141620244 N chr8 141620608 N DEL 5
A00404:156:HV37TDSXX:1:1330:5457:7247 chr8 141620244 N chr8 141620608 N DEL 11
A00404:155:HV27LDSXX:1:2113:31765:35180 chr8 141620206 N chr8 141620479 N DEL 3
A00404:156:HV37TDSXX:4:1239:14461:2863 chr8 141620335 N chr8 141620426 N DEL 7
A00404:155:HV27LDSXX:4:2530:4453:1282 chr12 132535915 N chr12 132535995 N DEL 13
A00297:158:HT275DSXX:2:2635:4327:29183 chr12 132535918 N chr12 132536047 N DEL 22
A00404:156:HV37TDSXX:3:2647:18548:34992 chrX 64680713 N chrX 64680818 N DUP 1
A00297:158:HT275DSXX:4:2327:1895:24095 chrX 1296674 N chrX 1296789 N DEL 4
A00404:155:HV27LDSXX:4:2210:13413:22373 chrX 1296677 N chrX 1296792 N DEL 5
A00404:156:HV37TDSXX:4:2445:16432:19930 chr5 148212697 N chr5 148212918 N DEL 5
A00404:156:HV37TDSXX:4:1349:10890:19758 chr1 143497448 N chr1 143497787 N DUP 5
A00404:156:HV37TDSXX:3:2367:8296:29481 chr1 143497359 N chr1 143497794 N DUP 13
A00404:155:HV27LDSXX:2:2302:6876:11459 chr2 3319833 N chr2 3319991 N DUP 8
A00404:155:HV27LDSXX:4:2144:30120:12195 chr2 3319833 N chr2 3319991 N DUP 8
A00404:155:HV27LDSXX:4:2144:30770:14043 chr2 3319833 N chr2 3319991 N DUP 8
A00404:155:HV27LDSXX:4:2144:30843:14293 chr2 3319828 N chr2 3319986 N DUP 8
A00404:155:HV27LDSXX:4:1519:21947:29199 chr2 3319976 N chr2 3320344 N DUP 1
A00404:155:HV27LDSXX:2:1224:23466:1485 chr2 3319972 N chr2 3320068 N DEL 20
A00404:155:HV27LDSXX:4:2411:20907:19476 chr2 3319972 N chr2 3320068 N DEL 20
A00404:156:HV37TDSXX:1:1112:8278:11350 chr2 3320032 N chr2 3320252 N DUP 12
A00297:158:HT275DSXX:4:2607:17734:21809 chr2 3319825 N chr2 3320176 N DUP 39
A00404:155:HV27LDSXX:2:1423:30662:13385 chr2 3319825 N chr2 3320176 N DUP 41
A00404:155:HV27LDSXX:1:1544:18719:30499 chr2 3319962 N chr2 3320197 N DEL 1
A00404:156:HV37TDSXX:4:2545:16758:16861 chr9 128507817 N chr9 128508110 N DEL 15
A00297:158:HT275DSXX:3:1203:15519:27868 chr8 143503733 N chr8 143503798 N DEL 15
A00404:155:HV27LDSXX:2:2512:15998:11350 chr8 143503738 N chr8 143503803 N DEL 10
A00404:156:HV37TDSXX:1:1345:7690:8453 chr8 143503744 N chr8 143503809 N DEL 4
A00404:156:HV37TDSXX:1:2211:20003:11021 chr8 143503745 N chr8 143503810 N DEL 3
A00404:156:HV37TDSXX:1:2328:26341:23876 chr8 143503742 N chr8 143503807 N DEL 6
A00404:156:HV37TDSXX:1:2625:10285:29199 chr8 143503745 N chr8 143503810 N DEL 3
A00404:156:HV37TDSXX:4:2363:17318:33238 chr8 143503744 N chr8 143503809 N DEL 4
A00297:158:HT275DSXX:4:1444:8775:28087 chr21 45484315 N chr21 45484448 N DEL 7
A00404:156:HV37TDSXX:4:1531:8874:20588 chr21 45484366 N chr21 45484623 N DEL 49
A00404:156:HV37TDSXX:3:2323:28881:16157 chr6 73791268 N chr6 73791347 N DUP 6
A00404:155:HV27LDSXX:2:1465:22968:30624 chr20 57962365 N chr20 57962428 N DEL 1
A00297:158:HT275DSXX:4:1262:4689:10081 chr4 126101007 N chr4 126101166 N DEL 7
A00404:155:HV27LDSXX:3:1429:13358:30264 chr4 126101056 N chr4 126101111 N DEL 24
A00404:155:HV27LDSXX:1:1406:5972:35822 chr4 126101005 N chr4 126101072 N DUP 14
A00297:158:HT275DSXX:2:2118:11930:4053 chr4 126101056 N chr4 126101111 N DEL 23
A00404:155:HV27LDSXX:3:2635:3206:34068 chr4 126101056 N chr4 126101111 N DEL 24
A00404:155:HV27LDSXX:3:2444:19452:15859 chr4 126101132 N chr4 126101189 N DEL 17
A00404:155:HV27LDSXX:1:1335:25708:2206 chr4 126101024 N chr4 126101093 N DEL 15
A00404:155:HV27LDSXX:3:2548:22345:32236 chr4 126101018 N chr4 126101264 N DUP 8
A00404:155:HV27LDSXX:4:2332:8169:31548 chr4 126101116 N chr4 126101264 N DUP 10
A00297:158:HT275DSXX:3:2414:30074:3787 chr4 126101116 N chr4 126101264 N DUP 10
A00297:158:HT275DSXX:3:1544:5999:7467 chr1 47322565 N chr1 47322735 N DEL 31
A00297:158:HT275DSXX:1:1256:27679:4147 chr1 47322547 N chr1 47322717 N DEL 20
A00404:155:HV27LDSXX:1:2176:25102:16313 chr17 82909595 N chr17 82909662 N DEL 5
A00404:156:HV37TDSXX:3:2625:29405:16313 chr17 82909595 N chr17 82909662 N DEL 5
A00297:158:HT275DSXX:3:2144:8811:35728 chr17 82909576 N chr17 82909779 N DEL 5
A00297:158:HT275DSXX:3:2506:6560:28166 chr17 82909595 N chr17 82909662 N DEL 5
A00404:155:HV27LDSXX:2:2219:18023:31704 chr17 82909595 N chr17 82909662 N DEL 5
A00404:155:HV27LDSXX:3:2505:26169:18505 chr17 82909595 N chr17 82909662 N DEL 5
A00297:158:HT275DSXX:3:1624:26124:8218 chr17 82909611 N chr17 82909814 N DEL 5
A00404:155:HV27LDSXX:3:1610:14082:22717 chr17 82909620 N chr17 82909685 N DUP 2
A00297:158:HT275DSXX:2:2452:5240:24878 chr11 112323985 N chr11 112324974 N DEL 5
A00404:155:HV27LDSXX:3:1126:9308:5368 chr11 112323987 N chr11 112324976 N DEL 5
A00404:155:HV27LDSXX:1:2309:10583:21543 chr9 136252481 N chr9 136252533 N DUP 5
A00404:156:HV37TDSXX:1:1355:29866:23124 chr10 31970667 N chr10 31970718 N DEL 5
A00404:155:HV27LDSXX:4:1326:20383:2597 chr10 31970661 N chr10 31970837 N DUP 7
A00404:156:HV37TDSXX:4:2169:32814:25128 chr10 31970661 N chr10 31970837 N DUP 7
A00404:155:HV27LDSXX:4:2350:2067:3537 chr10 31970843 N chr10 31971020 N DEL 5
A00297:158:HT275DSXX:1:1332:7862:3051 chr2 16649563 N chr2 16649708 N DUP 5
A00404:156:HV37TDSXX:3:2357:15248:26052 chr7 157867529 N chr7 157867664 N DEL 5
A00404:155:HV27LDSXX:4:2218:10945:3161 chr7 157867520 N chr7 157867689 N DEL 5
A00297:158:HT275DSXX:1:2274:10791:21652 chr5 82139691 N chr5 82139900 N DEL 5
A00404:155:HV27LDSXX:4:1343:12807:19288 chr5 82139520 N chr5 82139794 N DEL 5
A00404:155:HV27LDSXX:2:1147:25572:24048 chr5 82139472 N chr5 82139823 N DEL 5
A00297:158:HT275DSXX:3:2533:5132:31485 chr5 82139877 N chr5 82139954 N DUP 14
A00297:158:HT275DSXX:3:2125:5122:4163 chr5 82139957 N chr5 82140008 N DEL 5
A00297:158:HT275DSXX:1:2443:5511:4241 chr5 82139885 N chr5 82140061 N DUP 4
A00404:156:HV37TDSXX:1:2449:10257:36135 chr5 82139863 N chr5 82139993 N DEL 1
A00404:156:HV37TDSXX:2:2327:14118:20650 chr7 96816592 N chr7 96816673 N DUP 8
A00297:158:HT275DSXX:2:2611:24876:8187 chr7 96816553 N chr7 96816649 N DEL 5
A00297:158:HT275DSXX:1:1627:13910:4351 chr4 123498552 N chr4 123498655 N DUP 15
A00404:156:HV37TDSXX:4:1278:6949:27054 chr4 123498535 N chr4 123498723 N DUP 5
A00404:155:HV27LDSXX:3:2408:1642:4460 chr4 123498761 N chr4 123498826 N DUP 5
A00297:158:HT275DSXX:2:1315:8712:3991 chr19 38124426 N chr19 38124541 N DEL 19
A00297:158:HT275DSXX:1:1366:29514:24518 chr19 38124361 N chr19 38124440 N DUP 5
A00404:156:HV37TDSXX:1:2221:17743:8641 chr19 38124363 N chr19 38124442 N DUP 5
A00404:155:HV27LDSXX:4:2328:30779:20447 chr19 38124361 N chr19 38124440 N DUP 5
A00404:156:HV37TDSXX:4:2640:29921:5556 chr19 38124361 N chr19 38124440 N DUP 5
A00404:156:HV37TDSXX:3:1515:24053:21574 chr19 38124361 N chr19 38124440 N DUP 5
A00404:155:HV27LDSXX:4:1602:9932:9987 chr19 38124361 N chr19 38124440 N DUP 5
A00297:158:HT275DSXX:4:2628:24569:32831 chr19 38124587 N chr19 38124744 N DEL 11
A00404:155:HV27LDSXX:4:1407:30870:21042 chr21 42782092 N chr21 42782208 N DEL 5
A00404:155:HV27LDSXX:4:2563:17255:32409 chr5 167870704 N chr5 167870856 N DEL 3
A00404:156:HV37TDSXX:1:1312:24831:32659 chr4 40147886 N chr4 40148044 N DEL 9
A00404:156:HV37TDSXX:2:1158:22996:10128 chr4 40147962 N chr4 40148156 N DEL 24
A00404:155:HV27LDSXX:1:1363:29541:19742 chr4 40147965 N chr4 40148159 N DEL 10
A00404:155:HV27LDSXX:1:2568:18756:28119 chrX 1453341 N chrX 1453418 N DUP 7
A00404:155:HV27LDSXX:1:2568:18783:29136 chrX 1453341 N chrX 1453418 N DUP 7
A00404:156:HV37TDSXX:2:1554:8395:8735 chrX 1453341 N chrX 1453418 N DUP 7
A00404:155:HV27LDSXX:2:1221:26169:34726 chrX 1453173 N chrX 1453356 N DEL 9
A00404:155:HV27LDSXX:3:2378:11044:19836 chr17 49020082 N chr17 49020137 N DEL 6
A00404:156:HV37TDSXX:1:1307:4481:36370 chr17 49020082 N chr17 49020137 N DEL 13
A00404:155:HV27LDSXX:1:1169:21748:35869 chr3 162318974 N chr3 162319101 N DEL 3
A00404:155:HV27LDSXX:4:1210:7319:17487 chr3 162318974 N chr3 162319101 N DEL 3
A00404:155:HV27LDSXX:4:1671:32714:33599 chr3 162318974 N chr3 162319101 N DEL 3
A00297:158:HT275DSXX:2:1641:6903:14826 chr3 162318983 N chr3 162319110 N DEL 28
A00297:158:HT275DSXX:4:2205:23637:33755 chr3 162318983 N chr3 162319110 N DEL 29
A00297:158:HT275DSXX:1:1367:27742:17472 chr3 162318983 N chr3 162319110 N DEL 37
A00297:158:HT275DSXX:1:1367:28040:18145 chr3 162318983 N chr3 162319110 N DEL 37
A00404:156:HV37TDSXX:1:2367:31168:36245 chr3 162318983 N chr3 162319110 N DEL 45
A00297:158:HT275DSXX:2:2149:7690:5353 chr3 162318983 N chr3 162319110 N DEL 35
A00297:158:HT275DSXX:4:2556:14543:3912 chr3 162318983 N chr3 162319110 N DEL 29
A00297:158:HT275DSXX:2:2117:30635:32628 chr3 162318983 N chr3 162319110 N DEL 29
A00404:156:HV37TDSXX:1:2370:30924:21699 chr3 162318983 N chr3 162319110 N DEL 29
A00404:156:HV37TDSXX:2:1368:23303:34115 chr3 162318983 N chr3 162319110 N DEL 29
A00404:155:HV27LDSXX:4:2102:21947:34835 chr3 162318983 N chr3 162319110 N DEL 13
A00404:156:HV37TDSXX:1:2146:15393:15311 chr3 162318983 N chr3 162319110 N DEL 24
A00297:158:HT275DSXX:3:1339:19000:17550 chr3 162318983 N chr3 162319110 N DEL 22
A00404:155:HV27LDSXX:4:2642:28510:22310 chr3 162318983 N chr3 162319110 N DEL 5
A00404:155:HV27LDSXX:4:2642:28519:22294 chr3 162318983 N chr3 162319110 N DEL 10
A00404:155:HV27LDSXX:4:2642:28836:22905 chr3 162318983 N chr3 162319110 N DEL 10
A00297:158:HT275DSXX:4:1441:23791:28354 chr3 162318984 N chr3 162319111 N DEL 10
A00404:155:HV27LDSXX:3:1367:14398:31000 chr3 162319121 N chr3 162319528 N DUP 5
A00404:156:HV37TDSXX:1:2648:19886:4335 chr3 162318983 N chr3 162319110 N DEL 16
A00404:156:HV37TDSXX:1:1410:12536:33160 chr3 162318918 N chr3 162319227 N DUP 10
A00297:158:HT275DSXX:4:1501:32931:16752 chr3 162318918 N chr3 162319227 N DUP 5
A00404:156:HV37TDSXX:2:1116:32714:36198 chr3 162318918 N chr3 162319227 N DUP 5
A00404:156:HV37TDSXX:4:1126:26955:19617 chr3 162318918 N chr3 162319227 N DUP 10
A00404:155:HV27LDSXX:4:1210:7319:17487 chr3 162318918 N chr3 162319227 N DUP 14
A00297:158:HT275DSXX:2:1337:29848:6903 chr3 162318931 N chr3 162319338 N DEL 1
A00404:156:HV37TDSXX:2:2354:30635:21449 chr3 162319441 N chr3 162319532 N DEL 10
A00404:156:HV37TDSXX:2:2354:30906:21449 chr3 162319441 N chr3 162319532 N DEL 10
A00297:158:HT275DSXX:4:1462:5647:17472 chr3 162319441 N chr3 162319532 N DEL 10
A00404:155:HV27LDSXX:1:1169:21748:35869 chr3 162319219 N chr3 162319442 N DEL 10
A00404:155:HV27LDSXX:2:1452:1958:33786 chr3 162319471 N chr3 162319532 N DEL 3
A00404:156:HV37TDSXX:3:2245:5692:6402 chr3 162319441 N chr3 162319532 N DEL 10
A00404:155:HV27LDSXX:1:1350:11288:36511 chr3 162319441 N chr3 162319532 N DEL 10
A00404:155:HV27LDSXX:3:1469:7916:14888 chr3 162319474 N chr3 162319535 N DEL 10
A00404:155:HV27LDSXX:2:2315:15239:1736 chr3 162319474 N chr3 162319535 N DEL 10
A00297:158:HT275DSXX:1:2257:6677:32941 chr3 162319441 N chr3 162319532 N DEL 10
A00404:155:HV27LDSXX:1:1360:5891:5995 chr3 162319441 N chr3 162319532 N DEL 10
A00404:155:HV27LDSXX:1:1660:27715:20901 chr3 162319441 N chr3 162319532 N DEL 10
A00297:158:HT275DSXX:1:1258:24632:32784 chr3 162319441 N chr3 162319532 N DEL 10
A00404:155:HV27LDSXX:3:2214:2076:6809 chr3 162319431 N chr3 162319490 N DUP 24
A00404:156:HV37TDSXX:4:2638:30101:25379 chr3 162319456 N chr3 162319575 N DUP 15
A00404:156:HV37TDSXX:1:1244:13205:29684 chr3 162319456 N chr3 162319575 N DUP 14
A00404:156:HV37TDSXX:4:2251:10746:4539 chr3 162319456 N chr3 162319575 N DUP 14
A00404:156:HV37TDSXX:3:2132:29550:26522 chr3 162319419 N chr3 162319508 N DUP 42
A00404:156:HV37TDSXX:1:1447:15908:21997 chr3 162319419 N chr3 162319508 N DUP 43
A00297:158:HT275DSXX:2:2542:20898:9377 chr3 162319420 N chr3 162319509 N DUP 29
A00404:155:HV27LDSXX:1:1626:32108:31109 chr3 162319420 N chr3 162319509 N DUP 29
A00297:158:HT275DSXX:4:2577:9408:12806 chr3 162318967 N chr3 162319468 N DEL 3
A00404:155:HV27LDSXX:3:2336:29613:32925 chr3 162318967 N chr3 162319468 N DEL 3
A00297:158:HT275DSXX:1:2448:21441:22623 chr3 162319039 N chr3 162319536 N DEL 7
A00404:156:HV37TDSXX:2:1651:22507:25723 chr3 162319039 N chr3 162319536 N DEL 7
A00297:158:HT275DSXX:1:2638:31087:34976 chr3 162318938 N chr3 162319531 N DEL 12
A00404:156:HV37TDSXX:2:1446:23592:30514 chr3 162318938 N chr3 162319531 N DEL 12
A00404:155:HV27LDSXX:4:2674:23484:14794 chr3 162318938 N chr3 162319531 N DEL 12
A00404:155:HV27LDSXX:3:1417:4643:34710 chr3 162319040 N chr3 162319537 N DEL 7
A00404:156:HV37TDSXX:1:1229:16550:1939 chr8 62345511 N chr8 62345604 N DUP 9
A00404:155:HV27LDSXX:4:1157:31530:30608 chr8 62345464 N chr8 62345537 N DUP 7
A00404:156:HV37TDSXX:2:2469:7753:32800 chr8 62345498 N chr8 62345675 N DUP 22
A00404:156:HV37TDSXX:1:1220:32506:16360 chr8 62345457 N chr8 62345730 N DUP 1
A00297:158:HT275DSXX:3:1608:25382:31454 chr8 62345577 N chr8 62345662 N DEL 12
A00297:158:HT275DSXX:4:2547:2672:7059 chr8 62345577 N chr8 62345662 N DEL 9
A00404:156:HV37TDSXX:1:2124:3848:27414 chr8 62345577 N chr8 62345662 N DEL 9
A00297:158:HT275DSXX:2:2349:5710:23062 chr8 62345577 N chr8 62345662 N DEL 9
A00297:158:HT275DSXX:4:2128:20844:27258 chr8 62345478 N chr8 62345665 N DEL 9
A00404:156:HV37TDSXX:1:1658:30617:14090 chr8 62345470 N chr8 62345669 N DEL 7
A00297:158:HT275DSXX:3:1337:30346:6668 chr8 62345491 N chr8 62345766 N DEL 5
A00297:158:HT275DSXX:1:1654:24325:33379 chr8 62345491 N chr8 62345766 N DEL 5
A00404:156:HV37TDSXX:1:1363:21658:20306 chr8 62345491 N chr8 62345766 N DEL 5
A00297:158:HT275DSXX:1:2343:21450:22608 chr8 62345491 N chr8 62345766 N DEL 5
A00404:155:HV27LDSXX:2:1340:25473:26725 chr8 62345491 N chr8 62345766 N DEL 5
A00404:155:HV27LDSXX:2:1340:26738:26381 chr8 62345491 N chr8 62345766 N DEL 5
A00404:155:HV27LDSXX:3:1158:9471:20055 chr8 62345491 N chr8 62345766 N DEL 5
A00297:158:HT275DSXX:2:1620:13612:9314 chr8 62345525 N chr8 62345772 N DEL 5
A00404:156:HV37TDSXX:1:2508:11623:27258 chr3 129362618 N chr3 129362873 N DEL 5
A00404:156:HV37TDSXX:1:2508:11623:27258 chr3 129362618 N chr3 129362873 N DEL 5
A00404:156:HV37TDSXX:3:1672:3920:12164 chr3 129362570 N chr3 129363300 N DEL 5
A00297:158:HT275DSXX:1:2206:13485:28729 chr3 129362570 N chr3 129363300 N DEL 5
A00297:158:HT275DSXX:2:2429:25572:31908 chr3 129362502 N chr3 129362673 N DUP 9
A00404:156:HV37TDSXX:4:2615:6207:11490 chr3 129362518 N chr3 129363373 N DUP 5
A00404:155:HV27LDSXX:1:1521:12138:20917 chr3 129362594 N chr3 129362898 N DEL 10
A00297:158:HT275DSXX:1:2375:29071:10347 chr3 129362495 N chr3 129362926 N DEL 1
A00404:155:HV27LDSXX:3:2107:8350:1078 chr3 129363014 N chr3 129363318 N DEL 9
A00297:158:HT275DSXX:2:2359:17264:7968 chr3 129362564 N chr3 129363118 N DEL 5
A00297:158:HT275DSXX:4:2556:31250:33880 chr3 129362564 N chr3 129363118 N DEL 5
A00404:156:HV37TDSXX:1:2314:24397:26177 chr3 129362757 N chr3 129363135 N DEL 5
A00404:155:HV27LDSXX:2:1315:10538:31454 chr3 129362868 N chr3 129363244 N DUP 5
A00297:158:HT275DSXX:2:2316:10908:35978 chr3 129362518 N chr3 129363373 N DUP 5
A00297:158:HT275DSXX:1:1635:7175:15076 chr3 129362518 N chr3 129363373 N DUP 5
A00404:155:HV27LDSXX:3:2564:12454:8782 chr3 129362518 N chr3 129362644 N DUP 5
A00404:155:HV27LDSXX:4:1308:31864:15562 chr3 129362570 N chr3 129363300 N DEL 4
A00404:155:HV27LDSXX:4:1308:31864:15562 chr3 129362604 N chr3 129363334 N DEL 5
A00297:158:HT275DSXX:3:2236:20672:11804 chr3 129362604 N chr3 129363334 N DEL 5
A00297:158:HT275DSXX:1:1635:7175:15076 chr3 129362483 N chr3 129363388 N DUP 7
A00297:158:HT275DSXX:3:1205:1732:31015 chr3 129362483 N chr3 129363388 N DUP 9
A00404:155:HV27LDSXX:4:2673:2157:28964 chr3 129362655 N chr3 129363339 N DEL 8
A00297:158:HT275DSXX:1:2447:19859:9987 chr3 129362651 N chr3 129363283 N DEL 5
A00404:155:HV27LDSXX:3:2108:11876:1360 chr3 129362651 N chr3 129363283 N DEL 5
A00297:158:HT275DSXX:3:2406:29713:26584 chr3 129363310 N chr3 129363407 N DUP 5
A00297:158:HT275DSXX:3:1651:4842:33332 chr3 129362630 N chr3 129363407 N DUP 1
A00297:158:HT275DSXX:3:2451:28980:18051 chr3 129362630 N chr3 129363407 N DUP 2
A00404:155:HV27LDSXX:3:2639:12906:23531 chr3 129362630 N chr3 129363407 N DUP 5
A00404:155:HV27LDSXX:2:2222:18213:1752 chr3 129362472 N chr3 129363424 N DUP 6
A00297:158:HT275DSXX:2:1505:30671:36605 chr3 129362901 N chr3 129363279 N DEL 2
A00404:155:HV27LDSXX:1:1409:23439:17472 chr3 129363315 N chr3 129363412 N DUP 5
A00404:155:HV27LDSXX:4:1252:11125:1689 chr3 129362472 N chr3 129363424 N DUP 6
A00297:158:HT275DSXX:2:1332:22824:7858 chr19 36247185 N chr19 36247249 N DEL 1
A00404:156:HV37TDSXX:1:1470:14172:11350 chr15 95965534 N chr15 95965846 N DEL 16
A00297:158:HT275DSXX:3:2614:32072:23531 chr15 95965750 N chr15 95966061 N DEL 15
A00404:156:HV37TDSXX:2:1260:21612:22670 chr16 73173095 N chr16 73173167 N DEL 5
A00404:156:HV37TDSXX:1:1659:19804:17534 chr16 73173095 N chr16 73173169 N DEL 4
A00404:156:HV37TDSXX:4:1437:23990:11224 chr17 3656229 N chr17 3656342 N DUP 5
A00297:158:HT275DSXX:3:1256:32904:25441 chr17 3656355 N chr17 3656409 N DEL 16
A00404:155:HV27LDSXX:3:2652:21404:29951 chr3 54265749 N chr3 54265844 N DEL 5
A00404:156:HV37TDSXX:2:2662:19506:12070 chr3 54265749 N chr3 54265844 N DEL 5
A00404:156:HV37TDSXX:4:2554:20681:34397 chr3 54265749 N chr3 54265844 N DEL 5
A00404:156:HV37TDSXX:4:1419:8820:11945 chr3 54265749 N chr3 54265844 N DEL 5
A00404:155:HV27LDSXX:2:1314:3730:2409 chr3 54265749 N chr3 54265844 N DEL 5
A00297:158:HT275DSXX:4:1267:29414:19147 chr3 54265749 N chr3 54265844 N DEL 5
A00404:156:HV37TDSXX:2:2272:25861:21230 chr3 54265749 N chr3 54265844 N DEL 5
A00404:156:HV37TDSXX:4:1472:30870:17785 chr3 54265749 N chr3 54265844 N DEL 5
A00404:156:HV37TDSXX:4:2472:29035:24439 chr3 54265749 N chr3 54265844 N DEL 5
A00297:158:HT275DSXX:1:1529:23936:30389 chr4 189550597 N chr4 189550734 N DEL 5
A00297:158:HT275DSXX:2:2612:31150:31015 chr4 189550597 N chr4 189550734 N DEL 5
A00404:156:HV37TDSXX:2:1271:26449:19210 chr4 189550609 N chr4 189550678 N DEL 5
A00297:158:HT275DSXX:1:2145:14931:23844 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:2:1630:3314:25895 chr4 189550609 N chr4 189550678 N DEL 5
A00297:158:HT275DSXX:2:2645:25726:9659 chr4 189550609 N chr4 189550678 N DEL 5
A00297:158:HT275DSXX:2:1551:27163:30655 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:3:1636:22426:20666 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:3:2530:15492:21997 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:1:2659:10854:11459 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:1:2659:11288:10520 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:2:2127:10402:26741 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:2:1521:4616:2879 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:4:1673:28791:37043 chr4 189550609 N chr4 189550678 N DEL 5
A00404:156:HV37TDSXX:1:1334:30409:8876 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:2:1407:13096:8735 chr4 189550609 N chr4 189550678 N DEL 5
A00297:158:HT275DSXX:4:2506:4327:30185 chr4 189550609 N chr4 189550678 N DEL 5
A00297:158:HT275DSXX:1:2663:17598:6136 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:3:1318:24921:12618 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:2:2344:30101:14074 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:2:1476:13747:18004 chr4 189550609 N chr4 189550678 N DEL 5
A00404:156:HV37TDSXX:2:1535:19361:5462 chr4 189550609 N chr4 189550678 N DEL 5
A00404:156:HV37TDSXX:3:2332:14633:15718 chr4 189550609 N chr4 189550678 N DEL 5
A00404:156:HV37TDSXX:2:1322:22426:28682 chr4 189550609 N chr4 189550678 N DEL 5
A00404:156:HV37TDSXX:2:1322:22471:28635 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:3:1405:21594:5635 chr4 189550609 N chr4 189550678 N DEL 5
A00404:156:HV37TDSXX:4:2241:20699:30201 chr4 189550609 N chr4 189550678 N DEL 5
A00297:158:HT275DSXX:4:1165:13964:34851 chr4 189550609 N chr4 189550678 N DEL 5
A00404:155:HV27LDSXX:4:2127:23701:30170 chr4 189550597 N chr4 189550666 N DEL 11
A00297:158:HT275DSXX:1:1476:13512:30968 chr4 189550614 N chr4 189550749 N DUP 5
A00404:155:HV27LDSXX:1:1464:29134:32534 chr17 3746792 N chr17 3746926 N DEL 18
A00404:156:HV37TDSXX:3:2267:13123:20369 chr17 3746850 N chr17 3746984 N DEL 5
A00297:158:HT275DSXX:1:1547:6207:20259 chr6 143649046 N chr6 143649105 N DUP 8
A00404:155:HV27LDSXX:3:1503:30282:14293 chr13 41571427 N chr13 41571490 N DUP 5
A00297:158:HT275DSXX:1:1574:8938:1094 chr13 41571443 N chr13 41571502 N DEL 10
A00404:155:HV27LDSXX:3:1322:16794:20369 chr22 45092629 N chr22 45092693 N DEL 3
A00404:155:HV27LDSXX:4:2471:3079:22263 chr22 45092629 N chr22 45092693 N DEL 3
A00404:155:HV27LDSXX:4:2471:3088:22279 chr22 45092629 N chr22 45092693 N DEL 3
A00404:155:HV27LDSXX:2:2308:18964:9972 chr22 45092629 N chr22 45092693 N DEL 4
A00404:155:HV27LDSXX:2:2158:24053:24455 chr22 45092629 N chr22 45092693 N DEL 8
A00404:155:HV27LDSXX:4:1139:15872:1360 chr22 45092639 N chr22 45092703 N DEL 5
A00404:156:HV37TDSXX:4:1267:28944:27195 chr22 45092636 N chr22 45092700 N DEL 8
A00297:158:HT275DSXX:1:2271:18466:18349 chr22 45092640 N chr22 45092704 N DEL 4
A00297:158:HT275DSXX:1:2451:16577:18270 chr22 45092633 N chr22 45092697 N DEL 11
A00404:155:HV27LDSXX:3:2427:2908:33520 chr5 2280860 N chr5 2281249 N DUP 5
A00404:155:HV27LDSXX:1:2626:27507:27618 chr5 2280868 N chr5 2281429 N DUP 5
A00404:155:HV27LDSXX:1:2430:15691:3114 chr5 2281075 N chr5 2281465 N DUP 5
A00404:155:HV27LDSXX:4:2513:8006:16266 chr5 2281275 N chr5 2281476 N DEL 5
A00297:158:HT275DSXX:1:2576:19660:27555 chr5 2281270 N chr5 2281643 N DEL 31
A00404:155:HV27LDSXX:2:1359:14118:30452 chr5 2281266 N chr5 2281635 N DEL 15
A00404:156:HV37TDSXX:2:2627:10538:26381 chr5 2281266 N chr5 2281635 N DEL 13
A00404:155:HV27LDSXX:3:2624:26422:34976 chr5 2281278 N chr5 2281647 N DEL 3
A00404:156:HV37TDSXX:3:1255:22679:24236 chr6 20387066 N chr6 20387140 N DEL 2
A00297:158:HT275DSXX:4:1572:26395:27821 chr3 122868023 N chr3 122868158 N DEL 5
A00404:155:HV27LDSXX:3:1443:2519:27305 chr7 90744700 N chr7 90744828 N DEL 10
A00297:158:HT275DSXX:1:1577:29658:29152 chr7 90744783 N chr7 90744957 N DUP 11
A00404:155:HV27LDSXX:1:2410:20374:29074 chr7 90744784 N chr7 90744959 N DUP 5
A00404:156:HV37TDSXX:2:1307:23213:8093 chr7 90744784 N chr7 90744991 N DUP 7
A00404:156:HV37TDSXX:2:1307:23231:7936 chr7 90744784 N chr7 90744991 N DUP 7
A00404:156:HV37TDSXX:3:1138:32217:8375 chr7 90744784 N chr7 90744991 N DUP 7
A00404:156:HV37TDSXX:3:1264:25192:29966 chr7 90744784 N chr7 90744991 N DUP 7
A00404:155:HV27LDSXX:3:1244:14317:24377 chr7 90744784 N chr7 90744991 N DUP 7
A00404:156:HV37TDSXX:1:1259:14696:1986 chr7 90744784 N chr7 90744991 N DUP 7
A00404:156:HV37TDSXX:2:2340:24795:31845 chr7 90744784 N chr7 90744991 N DUP 7
A00404:155:HV27LDSXX:3:1436:10610:36401 chr7 90744784 N chr7 90744991 N DUP 7
A00404:156:HV37TDSXX:2:2178:21043:12759 chr7 90744784 N chr7 90744991 N DUP 7
A00297:158:HT275DSXX:4:1508:15709:4554 chr7 90744784 N chr7 90744991 N DUP 7
A00404:156:HV37TDSXX:2:2225:25437:14857 chr7 90744784 N chr7 90744991 N DUP 7
A00404:155:HV27LDSXX:4:1362:1344:18630 chr7 90744784 N chr7 90744991 N DUP 7
A00404:155:HV27LDSXX:1:1278:32425:8108 chr7 90744784 N chr7 90744991 N DUP 7
A00404:155:HV27LDSXX:2:2603:30454:32628 chr7 90744784 N chr7 90744991 N DUP 7
A00404:156:HV37TDSXX:1:1162:31792:5008 chr20 8570674 N chr20 8570761 N DEL 4
A00404:156:HV37TDSXX:3:2137:6994:24972 chr20 8570674 N chr20 8570761 N DEL 6
A00404:155:HV27LDSXX:3:2308:11116:7279 chr20 8570674 N chr20 8570761 N DEL 7
A00404:156:HV37TDSXX:4:2526:32371:15875 chr20 8570674 N chr20 8570761 N DEL 8
A00404:155:HV27LDSXX:4:1551:6605:11835 chr20 8570674 N chr20 8570761 N DEL 10
A00404:156:HV37TDSXX:4:1118:3857:4539 chr20 8570674 N chr20 8570761 N DEL 18
A00297:158:HT275DSXX:2:1155:7518:9502 chr20 8570684 N chr20 8570771 N DEL 5
A00297:158:HT275DSXX:2:1155:7898:9283 chr20 8570684 N chr20 8570771 N DEL 5
A00297:158:HT275DSXX:2:2506:27136:10535 chr9 34461262 N chr9 34461399 N DEL 15
A00297:158:HT275DSXX:3:2501:12084:17159 chr1 124835205 N chr1 124836049 N DUP 4
A00404:155:HV27LDSXX:4:1510:23402:36730 chr1 124835205 N chr1 124836049 N DUP 4
A00297:158:HT275DSXX:4:1176:21540:16063 chr1 43911727 N chr1 43911784 N DEL 1
A00404:156:HV37TDSXX:3:1239:4553:23218 chr1 43911684 N chr1 43911739 N DUP 20
A00404:155:HV27LDSXX:3:2676:1994:29340 chr1 43911684 N chr1 43911739 N DUP 20
A00297:158:HT275DSXX:2:2315:16468:8093 chr1 43911684 N chr1 43911739 N DUP 20
A00404:155:HV27LDSXX:3:2235:31430:31250 chr1 43911708 N chr1 43911793 N DEL 6
A00404:156:HV37TDSXX:3:1409:31204:25911 chr2 240226432 N chr2 240226591 N DUP 5
A00404:155:HV27LDSXX:3:2420:7591:20932 chr16 27294493 N chr16 27294849 N DEL 2
A00404:156:HV37TDSXX:4:1638:26051:30702 chr16 27294493 N chr16 27294659 N DEL 2
A00297:158:HT275DSXX:3:1105:5719:14998 chr16 27294493 N chr16 27294659 N DEL 5
A00404:155:HV27LDSXX:3:1367:12075:26944 chr16 27294526 N chr16 27294581 N DUP 3
A00404:155:HV27LDSXX:2:2154:14805:24251 chr16 27294526 N chr16 27294581 N DUP 5
A00297:158:HT275DSXX:4:2527:16351:27305 chr16 27294526 N chr16 27294746 N DUP 10
A00404:155:HV27LDSXX:3:1232:11641:25692 chr16 27294692 N chr16 27294771 N DUP 14
A00297:158:HT275DSXX:2:1542:14163:7545 chr16 27294615 N chr16 27294669 N DEL 11
A00297:158:HT275DSXX:4:1338:1515:22122 chr16 27294887 N chr16 27294953 N DEL 5
A00297:158:HT275DSXX:2:2134:10637:27868 chr16 27294856 N chr16 27294994 N DUP 17
A00404:155:HV27LDSXX:4:2167:9796:33771 chr16 27294849 N chr16 27294929 N DUP 13
A00297:158:HT275DSXX:3:1240:25319:8923 chr16 27294966 N chr16 27295032 N DUP 14
A00297:158:HT275DSXX:3:1237:15736:3223 chr16 27294855 N chr16 27295020 N DUP 12
A00404:155:HV27LDSXX:1:1623:10357:30953 chr16 27294856 N chr16 27294994 N DUP 16
A00404:156:HV37TDSXX:4:1123:2302:7733 chr16 27295017 N chr16 27295067 N DUP 26
A00404:155:HV27LDSXX:2:1662:22553:6762 chr16 27294967 N chr16 27295075 N DUP 18
A00297:158:HT275DSXX:4:2309:6479:13463 chr16 27294915 N chr16 27295018 N DEL 7
A00404:155:HV27LDSXX:3:1533:2474:17080 chr4 75884077 N chr4 75884379 N DEL 2
A00297:158:HT275DSXX:3:1248:19895:24987 chr4 75884095 N chr4 75884395 N DUP 5
A00404:156:HV37TDSXX:2:1363:6813:10848 chr4 75884095 N chr4 75884395 N DUP 5
A00297:158:HT275DSXX:3:1330:22272:9251 chr4 75884101 N chr4 75884401 N DUP 4
A00404:156:HV37TDSXX:3:2670:10908:25426 chr4 75883808 N chr4 75884121 N DEL 5
A00404:156:HV37TDSXX:4:2257:22941:2613 chr6 82589298 N chr6 82589379 N DUP 1
A00297:158:HT275DSXX:3:2662:9064:36010 chr6 82589298 N chr6 82589379 N DUP 15
A00404:156:HV37TDSXX:4:1103:27236:9674 chrX 972040 N chrX 972317 N DUP 1
A00404:156:HV37TDSXX:3:2437:11143:9893 chr13 103471555 N chr13 103471628 N DUP 5
A00404:156:HV37TDSXX:3:2437:11180:9893 chr13 103471555 N chr13 103471628 N DUP 5
A00404:155:HV27LDSXX:4:2202:2383:27383 chr13 103471555 N chr13 103471628 N DUP 5
A00297:158:HT275DSXX:4:1574:15103:30436 chr18 78693481 N chr18 78693533 N DEL 6
A00404:156:HV37TDSXX:4:2332:1841:4085 chr18 78693482 N chr18 78693534 N DEL 6
A00404:156:HV37TDSXX:1:1351:27977:4914 chr4 186252603 N chr4 186252736 N DUP 5
A00404:155:HV27LDSXX:1:2204:28257:28917 chr4 186252595 N chr4 186252759 N DUP 9
A00297:158:HT275DSXX:3:2266:16830:4335 chr4 186252707 N chr4 186252797 N DUP 22
A00404:156:HV37TDSXX:1:2352:22878:15562 chr4 186252707 N chr4 186252797 N DUP 26
A00297:158:HT275DSXX:2:1129:10954:26193 chr4 186252643 N chr4 186252874 N DUP 5
A00297:158:HT275DSXX:1:2505:17680:32330 chr4 186252711 N chr4 186252801 N DUP 29
A00297:158:HT275DSXX:1:1119:20437:17127 chr4 186252749 N chr4 186252903 N DEL 30
A00297:158:HT275DSXX:3:2634:10691:23140 chr20 61971684 N chr20 61971869 N DUP 8
A00404:156:HV37TDSXX:3:1563:29984:24486 chr20 61971669 N chr20 61971730 N DUP 5
A00404:155:HV27LDSXX:1:1664:11831:20666 chr20 61971672 N chr20 61971733 N DUP 5
A00404:155:HV27LDSXX:3:2315:19271:25473 chr20 61971697 N chr20 61971758 N DUP 3
A00404:155:HV27LDSXX:1:2272:23213:7404 chr20 61971700 N chr20 61971761 N DUP 1
A00404:156:HV37TDSXX:4:1541:20157:30420 chr20 61971639 N chr20 61971824 N DUP 5
A00404:155:HV27LDSXX:3:2656:10041:10833 chr20 61971639 N chr20 61971824 N DUP 10
A00404:155:HV27LDSXX:3:2363:28167:15264 chr20 61971743 N chr20 61971806 N DEL 5
A00297:158:HT275DSXX:4:2304:14796:4257 chr20 61971775 N chr20 61971836 N DUP 5
A00297:158:HT275DSXX:2:2402:24740:2691 chr20 61971668 N chr20 61971793 N DEL 5
A00297:158:HT275DSXX:2:2402:24740:2691 chr20 61971806 N chr20 61971867 N DUP 10
A00297:158:HT275DSXX:1:1535:28248:29590 chr20 61971757 N chr20 61971820 N DEL 1
A00404:156:HV37TDSXX:4:1665:20546:16783 chr9 84526482 N chr9 84526824 N DEL 34
A00404:156:HV37TDSXX:3:2420:25129:10379 chr9 84526575 N chr9 84526804 N DEL 5
A00297:158:HT275DSXX:2:1135:6406:29935 chr9 84526587 N chr9 84527637 N DUP 3
A00404:155:HV27LDSXX:2:1568:16649:28103 chr9 84526638 N chr9 84526715 N DEL 6
A00404:156:HV37TDSXX:3:1678:19180:13886 chr9 84526510 N chr9 84526700 N DEL 11
A00297:158:HT275DSXX:2:2230:14136:34334 chr9 84526829 N chr9 84527348 N DEL 5
A00297:158:HT275DSXX:3:1276:7491:12555 chr9 84526698 N chr9 84526777 N DEL 5
A00404:155:HV27LDSXX:4:1310:17942:5822 chr9 84526698 N chr9 84526777 N DEL 5
A00404:155:HV27LDSXX:3:2145:11216:34569 chr9 84526698 N chr9 84526777 N DEL 5
A00404:156:HV37TDSXX:3:2443:14064:4178 chr9 84526830 N chr9 84526905 N DUP 5
A00404:155:HV27LDSXX:2:2167:6171:15843 chr9 84526516 N chr9 84526932 N DUP 10
A00404:155:HV27LDSXX:4:1347:16694:6480 chr9 84526941 N chr9 84527234 N DEL 14
A00297:158:HT275DSXX:4:2120:27597:20415 chr9 84526986 N chr9 84527097 N DEL 5
A00404:156:HV37TDSXX:1:1466:28528:17080 chr9 84526633 N chr9 84527010 N DUP 5
A00404:155:HV27LDSXX:3:2119:16848:2456 chr9 84526508 N chr9 84526963 N DEL 5
A00297:158:HT275DSXX:1:2307:2700:32283 chr9 84526511 N chr9 84526966 N DEL 5
A00297:158:HT275DSXX:3:1276:7491:12555 chr9 84526895 N chr9 84526970 N DEL 1
A00404:155:HV27LDSXX:3:1343:12924:10692 chr9 84527060 N chr9 84527318 N DEL 26
A00404:155:HV27LDSXX:2:2167:6171:15843 chr9 84526535 N chr9 84526990 N DEL 5
A00404:155:HV27LDSXX:3:1343:12924:10692 chr9 84527064 N chr9 84527439 N DEL 39
A00297:158:HT275DSXX:2:1650:21215:24987 chr9 84527078 N chr9 84527189 N DEL 10
A00404:156:HV37TDSXX:2:1402:18991:36918 chr9 84527093 N chr9 84527350 N DUP 5
A00297:158:HT275DSXX:1:1523:9679:26710 chr9 84526614 N chr9 84527478 N DEL 25
A00404:156:HV37TDSXX:4:2325:27977:16626 chr9 84527589 N chr9 84527825 N DEL 31
A00404:156:HV37TDSXX:3:1455:24487:29496 chr9 84526566 N chr9 84527771 N DUP 5
A00297:158:HT275DSXX:3:1411:4915:33176 chr9 84527350 N chr9 84527772 N DUP 10
A00404:155:HV27LDSXX:3:2563:2103:22420 chr9 84527676 N chr9 84527834 N DUP 4
A00404:156:HV37TDSXX:2:1229:8205:32456 chr9 84527676 N chr9 84527834 N DUP 5
A00404:155:HV27LDSXX:2:1335:14371:25661 chr9 84527676 N chr9 84527834 N DUP 5
A00404:156:HV37TDSXX:4:1239:28519:12837 chr9 84527573 N chr9 84527849 N DEL 1
A00404:156:HV37TDSXX:4:1605:7636:8234 chr9 84527694 N chr9 84527854 N DEL 5
A00404:155:HV27LDSXX:3:1235:24433:21198 chr9 84527696 N chr9 84527856 N DEL 5
A00404:155:HV27LDSXX:2:1301:20419:23735 chr9 84527699 N chr9 84527859 N DEL 5
A00297:158:HT275DSXX:2:2208:13232:27070 chr9 84527437 N chr9 84527864 N DEL 5
A00297:158:HT275DSXX:4:2610:25807:30217 chr12 73107992 N chr12 73108162 N DEL 5
A00404:155:HV27LDSXX:3:2155:2772:5321 chrX 148704366 N chrX 148704421 N DUP 15
A00404:156:HV37TDSXX:4:1431:20862:24471 chrX 148704366 N chrX 148704421 N DUP 18
A00404:156:HV37TDSXX:4:1431:21703:24330 chrX 148704366 N chrX 148704421 N DUP 18
A00404:155:HV27LDSXX:2:1504:13485:12915 chrX 148704366 N chrX 148704421 N DUP 18
A00404:155:HV27LDSXX:1:1153:9408:17409 chrX 148704366 N chrX 148704421 N DUP 14
A00297:158:HT275DSXX:1:1375:27290:10551 chrX 148704370 N chrX 148704425 N DUP 15
A00297:158:HT275DSXX:2:2254:28709:23406 chrX 148704366 N chrX 148704421 N DUP 18
A00404:156:HV37TDSXX:3:2524:22562:12821 chrX 148704366 N chrX 148704449 N DUP 18
A00404:156:HV37TDSXX:4:2360:14552:18834 chrX 148704366 N chrX 148704449 N DUP 18
A00404:156:HV37TDSXX:3:1361:11062:26757 chrX 148704385 N chrX 148704504 N DUP 11
A00404:156:HV37TDSXX:4:1633:25346:22936 chrX 148704385 N chrX 148704504 N DUP 11
A00297:158:HT275DSXX:1:1125:12816:27602 chrX 148704396 N chrX 148704449 N DUP 16
A00404:155:HV27LDSXX:2:1256:27661:2300 chrX 148704408 N chrX 148704461 N DUP 3
A00404:156:HV37TDSXX:1:1132:21151:24345 chrX 148704396 N chrX 148704449 N DUP 10
A00297:158:HT275DSXX:2:1408:1533:6057 chrX 148704396 N chrX 148704449 N DUP 15
A00404:155:HV27LDSXX:2:1129:29414:16705 chrX 148704396 N chrX 148704449 N DUP 16
A00404:155:HV27LDSXX:3:2155:2772:5321 chrX 148704477 N chrX 148704530 N DEL 16
A00404:155:HV27LDSXX:2:1264:29604:28369 chrX 148704395 N chrX 148704530 N DEL 9
A00297:158:HT275DSXX:1:2543:25644:25207 chrX 148704401 N chrX 148704536 N DEL 9
A00297:158:HT275DSXX:1:2269:12048:6699 chrX 148704402 N chrX 148704537 N DEL 8
A00297:158:HT275DSXX:1:2269:13123:6026 chrX 148704402 N chrX 148704537 N DEL 8
A00297:158:HT275DSXX:1:2269:14407:11757 chrX 148704402 N chrX 148704537 N DEL 8
A00404:155:HV27LDSXX:2:1129:29414:16705 chrX 148704404 N chrX 148704539 N DEL 6
A00297:158:HT275DSXX:3:1438:18105:18818 chrX 148704405 N chrX 148704540 N DEL 5
A00297:158:HT275DSXX:2:1134:31638:7905 chr5 45207043 N chr5 45207157 N DEL 36
A00404:156:HV37TDSXX:2:2324:26503:1736 chr5 45207031 N chr5 45207145 N DEL 1
A00404:155:HV27LDSXX:3:1170:14922:1031 chrX 50447518 N chrX 50447571 N DUP 4
A00404:155:HV27LDSXX:1:1577:22634:2550 chr13 80981393 N chr13 80981464 N DUP 8
A00404:155:HV27LDSXX:4:2324:32669:32863 chr13 80981342 N chr13 80981395 N DEL 13
A00404:156:HV37TDSXX:2:1131:5303:9361 chr11 57025923 N chr11 57026010 N DUP 40
A00404:155:HV27LDSXX:1:1312:10429:7153 chr11 57025903 N chr11 57026035 N DEL 6
A00404:155:HV27LDSXX:3:2404:17517:25128 chr11 57025962 N chr11 57026037 N DEL 4
A00404:155:HV27LDSXX:3:2454:24885:14810 chr11 57025982 N chr11 57026051 N DEL 6
A00297:158:HT275DSXX:1:1621:16631:27477 chr11 57025982 N chr11 57026051 N DEL 6
A00404:156:HV37TDSXX:3:2367:8205:28698 chr11 57026061 N chr11 57026122 N DUP 5
A00404:155:HV27LDSXX:3:2321:29948:17691 chr12 114830922 N chr12 114831026 N DEL 6
A00404:155:HV27LDSXX:2:2224:12328:25786 chr21 44417099 N chr21 44417176 N DUP 5
A00297:158:HT275DSXX:1:2119:23818:36479 chr21 44417127 N chr21 44417242 N DUP 12
A00404:156:HV37TDSXX:2:2440:25952:28119 chr21 44417063 N chr21 44417218 N DUP 1
A00404:156:HV37TDSXX:2:1509:32624:33880 chr21 44417087 N chr21 44417166 N DEL 1
A00297:158:HT275DSXX:1:1403:15573:33849 chr21 44417074 N chr21 44417269 N DUP 5
A00404:156:HV37TDSXX:3:1218:30942:6449 chr21 44417241 N chr21 44417318 N DUP 5
A00404:156:HV37TDSXX:2:2166:30535:20212 chr1 125069391 N chr1 125069627 N DEL 5
A00404:156:HV37TDSXX:1:1169:12274:27132 chr1 125069284 N chr1 125069572 N DEL 2
A00404:155:HV27LDSXX:1:1524:26503:4586 chr1 125069483 N chr1 125069717 N DUP 10
A00297:158:HT275DSXX:3:2565:22923:1297 chr1 125069607 N chr1 125069776 N DUP 11
A00404:156:HV37TDSXX:1:1415:6958:1924 chr10 112594042 N chr10 112594216 N DEL 22
A00404:156:HV37TDSXX:3:1522:6569:35822 chr4 181151457 N chr4 181151557 N DEL 1
A00404:155:HV27LDSXX:1:2640:24460:22279 chr4 181151457 N chr4 181151557 N DEL 5
A00404:156:HV37TDSXX:4:2631:30029:24471 chr4 181151541 N chr4 181151632 N DUP 5
A00297:158:HT275DSXX:1:1170:4472:27117 chr16 67712862 N chr16 67713019 N DEL 30
A00297:158:HT275DSXX:2:1261:26440:6292 chr17 9471194 N chr17 9471309 N DEL 7
A00297:158:HT275DSXX:3:2574:3287:7310 chr20 26205917 N chr20 26205966 N DUP 12
A00297:158:HT275DSXX:2:2106:14290:10802 chr21 41829569 N chr21 41830037 N DEL 14
A00404:155:HV27LDSXX:4:1437:15727:34428 chr5 17773455 N chr5 17773533 N DEL 7
A00404:156:HV37TDSXX:1:2537:10872:8108 chr19 8611349 N chr19 8611429 N DEL 6
A00404:156:HV37TDSXX:1:2348:28519:24674 chr19 8611280 N chr19 8611478 N DEL 11
A00297:158:HT275DSXX:4:1642:25048:11835 chr16 59893097 N chr16 59893194 N DEL 4
A00404:156:HV37TDSXX:2:2652:21206:16297 chr5 78448006 N chr5 78448117 N DEL 12
A00404:155:HV27LDSXX:2:1152:21513:16485 chr1 95538565 N chr1 95538721 N DUP 5
A00297:158:HT275DSXX:1:2540:3287:30076 chr1 95538565 N chr1 95538721 N DUP 5
A00404:156:HV37TDSXX:4:1176:7184:31125 chr1 95538631 N chr1 95538721 N DUP 5
A00297:158:HT275DSXX:3:2663:2483:7733 chr1 95538558 N chr1 95538741 N DEL 2
A00297:158:HT275DSXX:1:1408:30861:2049 chr7 155934840 N chr7 155934899 N DEL 6
A00297:158:HT275DSXX:4:1139:8043:14199 chr7 155934840 N chr7 155934934 N DEL 12
A00297:158:HT275DSXX:2:1525:10945:9831 chr7 155934840 N chr7 155934934 N DEL 28
A00404:155:HV27LDSXX:1:1162:17852:25488 chrX 54630863 N chrX 54630924 N DUP 7
A00404:155:HV27LDSXX:4:1333:9959:16329 chr19 55266641 N chr19 55266803 N DEL 11
A00404:155:HV27LDSXX:1:1462:16016:12602 chr19 55266535 N chr19 55266645 N DUP 15
A00297:158:HT275DSXX:4:2378:31123:3818 chr19 55266535 N chr19 55266645 N DUP 28
A00404:156:HV37TDSXX:3:2418:8015:12211 chr19 55266535 N chr19 55266645 N DUP 28
A00404:156:HV37TDSXX:4:2609:16125:4554 chr19 55266535 N chr19 55266645 N DUP 19
A00404:155:HV27LDSXX:1:2348:4119:35274 chr19 55266609 N chr19 55266662 N DUP 7
A00297:158:HT275DSXX:4:1632:23945:27398 chr19 55266535 N chr19 55266645 N DUP 15
A00297:158:HT275DSXX:4:2632:18222:36119 chr19 55266535 N chr19 55266645 N DUP 15
A00404:155:HV27LDSXX:3:1232:17454:34945 chr19 55266634 N chr19 55266710 N DUP 27
A00297:158:HT275DSXX:4:1359:5466:22013 chr19 55266634 N chr19 55266710 N DUP 27
A00404:155:HV27LDSXX:4:1628:5782:16078 chr19 55266551 N chr19 55266627 N DEL 8
A00297:158:HT275DSXX:2:1332:31132:20901 chr19 55266637 N chr19 55266713 N DUP 10
A00404:155:HV27LDSXX:3:2339:18593:2910 chr19 55266704 N chr19 55266753 N DUP 16
A00297:158:HT275DSXX:1:2258:17969:8093 chr19 55266552 N chr19 55266646 N DEL 3
A00404:156:HV37TDSXX:4:1263:2636:21089 chr12 90223765 N chr12 90223876 N DEL 18
A00404:156:HV37TDSXX:2:1559:11053:34757 chr12 90223765 N chr12 90223876 N DEL 27
A00404:155:HV27LDSXX:3:1351:8522:4038 chr12 90223741 N chr12 90223887 N DEL 4
A00404:155:HV27LDSXX:1:2644:16604:32252 chr8 144125849 N chr8 144125909 N DEL 16
A00404:156:HV37TDSXX:2:2177:30969:16235 chr8 144126075 N chr8 144126195 N DEL 5
A00297:158:HT275DSXX:4:2246:22173:8077 chr8 144125791 N chr8 144126028 N DUP 1
A00404:156:HV37TDSXX:2:1238:23827:35055 chr8 144125796 N chr8 144125914 N DUP 2
A00297:158:HT275DSXX:4:2545:17110:33379 chr8 144125956 N chr8 144126045 N DUP 9
A00404:156:HV37TDSXX:4:2254:4906:23985 chr8 144126059 N chr8 144126120 N DEL 16
A00404:155:HV27LDSXX:3:1277:7066:4961 chr8 144125932 N chr8 144125992 N DEL 12
A00297:158:HT275DSXX:1:1365:9182:6997 chr8 144125783 N chr8 144126140 N DUP 13
A00404:156:HV37TDSXX:3:2269:30960:7263 chr8 144125767 N chr8 144126213 N DUP 29
A00297:158:HT275DSXX:3:1421:21368:7529 chr8 144125858 N chr8 144125917 N DUP 24
A00297:158:HT275DSXX:2:2204:6108:23187 chr8 144125846 N chr8 144125995 N DEL 22
A00404:156:HV37TDSXX:2:2457:30563:9862 chr8 144125792 N chr8 144126059 N DUP 30
A00404:155:HV27LDSXX:3:2229:28971:3098 chr8 144126059 N chr8 144126120 N DEL 20
A00404:155:HV27LDSXX:1:1678:10872:20415 chr8 144126059 N chr8 144126120 N DEL 21
A00297:158:HT275DSXX:1:2207:22616:23249 chr8 144125919 N chr8 144126069 N DEL 10
A00404:156:HV37TDSXX:1:2455:16767:16971 chr8 144125965 N chr8 144126054 N DUP 22
A00404:156:HV37TDSXX:1:2308:18331:1705 chr8 144125875 N chr8 144125995 N DEL 15
A00297:158:HT275DSXX:4:2124:4047:24815 chr8 144125890 N chr8 144126008 N DUP 5
A00404:156:HV37TDSXX:3:2269:30960:7263 chr8 144125851 N chr8 144125970 N DEL 22
A00404:156:HV37TDSXX:4:1110:13666:29543 chr8 144125921 N chr8 144126011 N DEL 8
A00404:156:HV37TDSXX:1:2661:16134:30561 chr8 144125861 N chr8 144126011 N DEL 6
A00404:155:HV27LDSXX:4:2625:24731:25003 chr8 144125777 N chr8 144126016 N DEL 6
A00404:155:HV27LDSXX:4:1335:5746:12540 chr8 144125995 N chr8 144126054 N DUP 24
A00297:158:HT275DSXX:2:2607:12943:35681 chr8 144125911 N chr8 144126059 N DUP 14
A00404:155:HV27LDSXX:1:1623:15881:19382 chr8 144126007 N chr8 144126155 N DUP 10
A00297:158:HT275DSXX:3:1266:8657:27696 chr8 144125908 N chr8 144126205 N DUP 3
A00404:155:HV27LDSXX:3:1665:11731:12132 chr8 144125918 N chr8 144126038 N DEL 5
A00404:155:HV27LDSXX:2:2140:10926:29935 chr8 144125803 N chr8 144126189 N DUP 5
A00404:156:HV37TDSXX:2:1313:4399:29403 chr8 144125764 N chr8 144125912 N DUP 42
A00404:156:HV37TDSXX:2:2362:21739:17660 chr8 144125783 N chr8 144126199 N DUP 32
A00404:156:HV37TDSXX:2:1625:32488:36119 chr8 144125775 N chr8 144126072 N DUP 16
A00404:155:HV27LDSXX:1:1543:25229:14810 chr8 144125995 N chr8 144126054 N DUP 25
A00297:158:HT275DSXX:4:1650:18665:9048 chr8 144125783 N chr8 144126050 N DUP 10
A00297:158:HT275DSXX:4:1267:27290:6511 chr8 144125792 N chr8 144126059 N DUP 14
A00404:156:HV37TDSXX:2:1604:2094:28855 chr8 144125862 N chr8 144126012 N DEL 10
A00404:155:HV27LDSXX:3:1113:16342:35587 chr8 144125803 N chr8 144125861 N DUP 20
A00404:155:HV27LDSXX:1:1429:17056:6480 chr8 144125827 N chr8 144125915 N DUP 5
A00404:155:HV27LDSXX:3:1173:7346:30248 chr8 144125887 N chr8 144126035 N DUP 27
A00404:156:HV37TDSXX:2:2265:18385:21778 chr8 144125991 N chr8 144126050 N DUP 20
A00404:156:HV37TDSXX:4:2365:14045:7654 chr8 144125788 N chr8 144125965 N DUP 25
A00404:155:HV27LDSXX:1:1654:23430:29919 chr8 144125797 N chr8 144125915 N DUP 1
A00404:156:HV37TDSXX:1:2308:18331:1705 chr8 144126059 N chr8 144126120 N DEL 29
A00404:156:HV37TDSXX:1:2155:23981:35164 chr8 144125851 N chr8 144126120 N DEL 15
A00404:155:HV27LDSXX:2:2110:19813:33489 chr8 144125927 N chr8 144125985 N DUP 5
A00297:158:HT275DSXX:4:2609:18267:8015 chr8 144125902 N chr8 144125960 N DUP 7
A00404:156:HV37TDSXX:3:1437:29487:29262 chr8 144125927 N chr8 144126194 N DUP 10
A00297:158:HT275DSXX:2:2105:12798:25347 chr8 144125753 N chr8 144125960 N DUP 15
A00404:155:HV27LDSXX:2:1263:25726:25817 chr8 144125995 N chr8 144126203 N DUP 33
A00404:156:HV37TDSXX:4:1344:3577:26349 chr8 144126025 N chr8 144126116 N DEL 6
A00404:155:HV27LDSXX:2:2528:11849:7200 chr8 144125866 N chr8 144126136 N DEL 23
A00404:155:HV27LDSXX:3:2436:28284:2347 chr8 144126000 N chr8 144126059 N DUP 22
A00404:156:HV37TDSXX:2:1625:32488:36119 chr8 144125906 N chr8 144125964 N DUP 40
A00404:155:HV27LDSXX:1:2330:15402:9345 chr8 144125761 N chr8 144125879 N DUP 12
A00297:158:HT275DSXX:1:1314:27181:16282 chr8 144126025 N chr8 144126146 N DEL 6
A00404:155:HV27LDSXX:2:1372:17463:14700 chr8 144125834 N chr8 144126101 N DUP 20
A00404:156:HV37TDSXX:3:1542:27181:31438 chr8 144125887 N chr8 144125975 N DUP 18
A00404:156:HV37TDSXX:1:1663:25174:5196 chr8 144125866 N chr8 144126016 N DEL 10
A00404:155:HV27LDSXX:3:2229:28971:3098 chr8 144125764 N chr8 144126061 N DUP 25
A00297:158:HT275DSXX:4:1347:25238:18176 chr8 144125882 N chr8 144126032 N DEL 14
A00297:158:HT275DSXX:3:1333:32533:5791 chr8 144125887 N chr8 144126095 N DUP 28
A00297:158:HT275DSXX:2:2403:19316:23954 chr8 144126059 N chr8 144126120 N DEL 23
A00404:155:HV27LDSXX:3:1375:24731:35775 chr8 144125858 N chr8 144125917 N DUP 28
A00297:158:HT275DSXX:1:1463:30852:6480 chr8 144125783 N chr8 144125960 N DUP 22
A00404:155:HV27LDSXX:3:2314:32588:21386 chr8 144125930 N chr8 144126048 N DUP 7
A00404:155:HV27LDSXX:3:2247:16785:3850 chr8 144125991 N chr8 144126050 N DUP 12
A00297:158:HT275DSXX:3:2370:7581:32315 chr8 144125927 N chr8 144126045 N DUP 5
A00404:156:HV37TDSXX:3:1302:13404:34225 chr8 144125902 N chr8 144126050 N DUP 2
A00297:158:HT275DSXX:2:2608:17155:4836 chr8 144125995 N chr8 144126203 N DUP 14
A00404:155:HV27LDSXX:1:1503:7618:31281 chr8 144125764 N chr8 144126061 N DUP 25
A00404:155:HV27LDSXX:4:1343:31222:22341 chr8 144125783 N chr8 144126199 N DUP 18
A00404:156:HV37TDSXX:3:1473:3278:13651 chr8 144125947 N chr8 144126036 N DUP 12
A00404:155:HV27LDSXX:1:1401:21703:25363 chr8 144126125 N chr8 144126213 N DUP 39
A00404:155:HV27LDSXX:1:1543:25229:14810 chr8 144125995 N chr8 144126054 N DUP 35
A00297:158:HT275DSXX:4:2629:19723:4022 chr8 144125927 N chr8 144126045 N DUP 12
A00404:156:HV37TDSXX:4:1536:27923:19633 chr8 144125910 N chr8 144126120 N DEL 16
A00404:155:HV27LDSXX:1:2534:12454:23062 chr8 144125816 N chr8 144125995 N DEL 17
A00297:158:HT275DSXX:2:1552:26793:22310 chr8 144125764 N chr8 144126061 N DUP 25
A00297:158:HT275DSXX:1:2270:30924:23109 chr8 144125918 N chr8 144126038 N DEL 5
A00404:155:HV27LDSXX:2:1464:20238:27336 chr8 144125947 N chr8 144126036 N DUP 16
A00297:158:HT275DSXX:2:2656:5565:36558 chr8 144125995 N chr8 144126203 N DUP 28
A00297:158:HT275DSXX:1:1248:16179:35587 chr8 144125792 N chr8 144126059 N DUP 30
A00297:158:HT275DSXX:4:1654:15646:20917 chr8 144126059 N chr8 144126120 N DEL 32
A00404:156:HV37TDSXX:4:2365:14045:7654 chr8 144125916 N chr8 144126094 N DUP 6
A00404:156:HV37TDSXX:2:1227:9281:2973 chr8 144125908 N chr8 144125998 N DEL 15
A00297:158:HT275DSXX:3:1421:21947:7404 chr8 144125858 N chr8 144125917 N DUP 24
A00404:155:HV27LDSXX:4:2663:19732:1658 chr8 144125834 N chr8 144125981 N DUP 7
A00404:155:HV27LDSXX:4:1162:3965:28494 chr8 144125996 N chr8 144126174 N DUP 21
A00404:156:HV37TDSXX:4:2251:2076:17832 chr8 144125765 N chr8 144126092 N DUP 3
A00404:156:HV37TDSXX:3:2667:16712:1501 chr8 144125906 N chr8 144125964 N DUP 40
A00404:156:HV37TDSXX:2:1241:25201:20870 chr8 144125970 N chr8 144126059 N DUP 5
A00297:158:HT275DSXX:3:2216:6741:30358 chr8 144125764 N chr8 144126061 N DUP 30
A00297:158:HT275DSXX:4:1347:25238:18176 chr8 144125995 N chr8 144126203 N DUP 32
A00404:156:HV37TDSXX:1:2655:17083:28197 chr8 144125853 N chr8 144126002 N DEL 20
A00404:156:HV37TDSXX:3:1570:30029:28573 chr8 144126097 N chr8 144126215 N DUP 30
A00404:155:HV27LDSXX:1:1375:13602:7138 chr8 144125995 N chr8 144126054 N DUP 21
A00297:158:HT275DSXX:3:1267:32524:31454 chr8 144126003 N chr8 144126122 N DUP 5
A00297:158:HT275DSXX:2:2203:20302:5807 chr8 144125962 N chr8 144126051 N DUP 12
A00404:155:HV27LDSXX:1:1327:14751:30013 chr8 144125792 N chr8 144125940 N DUP 15
A00297:158:HT275DSXX:4:1351:25979:23844 chr8 144126055 N chr8 144126116 N DEL 27
A00404:156:HV37TDSXX:2:2656:32651:21903 chr8 144125963 N chr8 144126024 N DEL 10
A00404:156:HV37TDSXX:1:2503:28845:8077 chr8 144125950 N chr8 144126039 N DUP 15
A00297:158:HT275DSXX:3:1266:8657:27696 chr8 144126059 N chr8 144126120 N DEL 31
A00404:155:HV27LDSXX:4:2449:31882:29622 chr8 144125995 N chr8 144126203 N DUP 30
A00404:155:HV27LDSXX:2:2529:16550:25394 chr8 144125866 N chr8 144126136 N DEL 14
A00404:155:HV27LDSXX:3:2509:27055:15781 chr8 144125858 N chr8 144125917 N DUP 17
A00404:155:HV27LDSXX:3:1522:16658:12148 chr8 144125995 N chr8 144126054 N DUP 20
A00404:156:HV37TDSXX:2:2550:25681:8703 chr8 144125896 N chr8 144126014 N DUP 5
A00404:156:HV37TDSXX:4:2409:27814:26177 chr8 144125898 N chr8 144125986 N DUP 5
A00297:158:HT275DSXX:2:2612:30789:17018 chr8 144125776 N chr8 144126221 N DUP 10
A00404:156:HV37TDSXX:1:1256:26485:15327 chr8 144125783 N chr8 144126140 N DUP 12
A00297:158:HT275DSXX:4:1640:28167:34929 chr8 144125842 N chr8 144125961 N DEL 1
A00404:155:HV27LDSXX:3:1257:22887:15233 chr8 144125789 N chr8 144126056 N DUP 17
A00404:156:HV37TDSXX:2:2550:26539:9189 chr8 144125910 N chr8 144126120 N DEL 12
A00297:158:HT275DSXX:4:2506:10791:13385 chr8 144125888 N chr8 144126036 N DUP 6
A00404:155:HV27LDSXX:2:2135:14335:30358 chr8 144125955 N chr8 144126016 N DEL 12
A00297:158:HT275DSXX:2:1632:24731:20588 chr8 144125995 N chr8 144126203 N DUP 25
A00297:158:HT275DSXX:1:2233:21540:14779 chr8 144125887 N chr8 144125975 N DUP 1
A00404:155:HV27LDSXX:2:1362:22968:30060 chr8 144125824 N chr8 144126003 N DEL 5
A00297:158:HT275DSXX:2:2619:21875:33426 chr8 144125823 N chr8 144126092 N DEL 8
A00404:155:HV27LDSXX:4:1362:24894:8688 chr8 144125826 N chr8 144126033 N DUP 5
A00404:156:HV37TDSXX:4:1344:3577:26349 chr8 144125899 N chr8 144126137 N DUP 6
A00404:156:HV37TDSXX:2:2550:26539:9189 chr8 144125896 N chr8 144126014 N DUP 5
A00297:158:HT275DSXX:4:2266:21106:16783 chr8 144125910 N chr8 144126120 N DEL 12
A00404:155:HV27LDSXX:3:2638:32090:10880 chr8 144125995 N chr8 144126203 N DUP 25
A00404:156:HV37TDSXX:1:2435:3233:14575 chr8 144125887 N chr8 144126035 N DUP 6
A00404:155:HV27LDSXX:1:1558:16595:9001 chr8 144125764 N chr8 144125853 N DUP 36
A00297:158:HT275DSXX:1:2615:4526:22545 chr8 144125875 N chr8 144125995 N DEL 15
A00404:155:HV27LDSXX:1:2639:9046:33160 chr8 144125881 N chr8 144126001 N DEL 20
A00404:156:HV37TDSXX:1:2144:30165:13933 chr8 144125917 N chr8 144126067 N DEL 10
A00404:156:HV37TDSXX:1:1256:26738:17801 chr8 144125771 N chr8 144126098 N DUP 16
A00297:158:HT275DSXX:2:2546:24668:21919 chr8 144125995 N chr8 144126173 N DUP 32
A00404:155:HV27LDSXX:3:1401:25599:1329 chr8 144125907 N chr8 144126204 N DUP 7
A00404:155:HV27LDSXX:4:2604:21513:2581 chr8 144125778 N chr8 144125898 N DEL 4
A00297:158:HT275DSXX:4:2418:32190:11835 chr8 144125838 N chr8 144126194 N DUP 10
A00404:155:HV27LDSXX:2:1370:28492:31203 chr8 144125999 N chr8 144126058 N DUP 15
A00404:155:HV27LDSXX:2:2146:25536:20196 chr8 144125764 N chr8 144126210 N DUP 23
A00404:155:HV27LDSXX:1:2542:21576:21136 chr8 144125991 N chr8 144126050 N DUP 7
A00297:158:HT275DSXX:4:1676:17381:3192 chr8 144125842 N chr8 144126081 N DEL 6
A00297:158:HT275DSXX:3:1144:18258:11318 chr8 144125887 N chr8 144126035 N DUP 29
A00297:158:HT275DSXX:4:2369:9824:17347 chr8 144125858 N chr8 144125917 N DUP 37
A00297:158:HT275DSXX:3:1416:1696:29450 chr8 144125769 N chr8 144125976 N DUP 11
A00404:156:HV37TDSXX:1:1574:25283:32972 chr8 144125784 N chr8 144126200 N DUP 14
A00297:158:HT275DSXX:4:2107:6614:31360 chr8 144125927 N chr8 144126045 N DUP 5
A00404:155:HV27LDSXX:1:2540:27163:18912 chr8 144125947 N chr8 144126036 N DUP 13
A00404:156:HV37TDSXX:1:1343:16631:5024 chr8 144125995 N chr8 144126173 N DUP 22
A00404:155:HV27LDSXX:2:2503:3658:36448 chr8 144125941 N chr8 144126178 N DUP 21
A00404:156:HV37TDSXX:2:2645:31494:5118 chr8 144125995 N chr8 144126173 N DUP 28
A00404:155:HV27LDSXX:4:1125:28212:18411 chr8 144125995 N chr8 144126173 N DUP 23
A00404:155:HV27LDSXX:4:1336:28818:31046 chr8 144125779 N chr8 144126018 N DEL 5
A00404:156:HV37TDSXX:3:2276:1452:18787 chr6 25137369 N chr6 25137478 N DEL 4
A00404:156:HV37TDSXX:2:2257:11053:16814 chr3 70211432 N chr3 70211721 N DEL 25
A00297:158:HT275DSXX:1:1178:18828:32127 chr3 70211440 N chr3 70211596 N DEL 23
A00404:156:HV37TDSXX:3:1378:28718:33692 chr3 70211414 N chr3 70211597 N DEL 44
A00404:155:HV27LDSXX:3:2103:30743:5478 chr3 70211492 N chr3 70211611 N DEL 10
A00404:155:HV27LDSXX:3:2103:32470:6120 chr3 70211492 N chr3 70211611 N DEL 10
A00404:155:HV27LDSXX:3:2103:32479:6136 chr3 70211492 N chr3 70211611 N DEL 10
A00404:156:HV37TDSXX:3:1263:13006:3161 chr3 70211492 N chr3 70211611 N DEL 19
A00404:156:HV37TDSXX:3:1263:13322:2895 chr3 70211492 N chr3 70211611 N DEL 19
A00404:155:HV27LDSXX:4:1438:31412:32283 chr3 70211492 N chr3 70211611 N DEL 31
A00404:156:HV37TDSXX:2:2106:27416:32534 chr3 70211568 N chr3 70211651 N DUP 22
A00404:155:HV27LDSXX:4:1348:8278:23249 chr3 70211556 N chr3 70211639 N DUP 27
A00404:155:HV27LDSXX:2:2155:19741:7185 chr3 70211596 N chr3 70211664 N DUP 2
A00404:156:HV37TDSXX:3:2151:23439:26710 chr3 70211496 N chr3 70211667 N DEL 24
A00404:155:HV27LDSXX:1:2607:26368:25457 chr3 70211556 N chr3 70211639 N DUP 27
A00404:155:HV27LDSXX:3:2271:31458:2675 chr3 70211670 N chr3 70211730 N DEL 9
A00297:158:HT275DSXX:2:2314:11243:29450 chr3 70211522 N chr3 70211725 N DEL 10
A00404:156:HV37TDSXX:3:1421:26982:30154 chr3 70211634 N chr3 70211736 N DEL 10
A00404:155:HV27LDSXX:4:2438:28592:17378 chr3 70211466 N chr3 70211728 N DEL 2
A00404:156:HV37TDSXX:1:1213:18891:21746 chr3 70211679 N chr3 70211834 N DEL 27
A00404:155:HV27LDSXX:2:2337:27923:23703 chr3 70211616 N chr3 70211855 N DEL 5
A00404:156:HV37TDSXX:1:2247:4960:20290 chr2 31805882 N chr2 31805971 N DEL 14
A00404:156:HV37TDSXX:1:2566:30662:9784 chr2 31805984 N chr2 31806163 N DUP 1
A00404:155:HV27LDSXX:2:2678:27471:30248 chr2 31805917 N chr2 31806094 N DEL 2
A00404:156:HV37TDSXX:1:2552:18475:2112 chr2 31805890 N chr2 31806109 N DEL 5
A00297:158:HT275DSXX:2:1646:31448:15060 chr2 31805940 N chr2 31806185 N DEL 19
A00404:155:HV27LDSXX:2:2477:25346:11976 chr7 155410040 N chr7 155410105 N DEL 5
A00404:155:HV27LDSXX:2:2243:30852:36198 chr7 155410061 N chr7 155410120 N DUP 6
A00297:158:HT275DSXX:1:1330:12481:25739 chr7 155410061 N chr7 155410120 N DUP 6
A00297:158:HT275DSXX:1:1330:12988:23923 chr7 155410061 N chr7 155410120 N DUP 6
A00404:155:HV27LDSXX:2:1359:1823:20275 chr7 155410061 N chr7 155410120 N DUP 6
A00404:156:HV37TDSXX:4:2566:5122:1783 chr17 670288 N chr17 670415 N DUP 5
A00297:158:HT275DSXX:1:1555:3604:32847 chr21 18690314 N chr21 18690899 N DEL 5
A00404:155:HV27LDSXX:3:2656:30544:31814 chr21 18690314 N chr21 18690388 N DEL 10
A00297:158:HT275DSXX:2:1141:16098:26021 chr21 18690396 N chr21 18690762 N DEL 15
A00404:156:HV37TDSXX:2:1413:22209:24674 chr21 18690387 N chr21 18690459 N DUP 5
A00404:155:HV27LDSXX:1:1230:29306:7842 chr21 18690334 N chr21 18690698 N DUP 5
A00404:155:HV27LDSXX:4:2654:1380:10457 chr21 18690543 N chr21 18690617 N DEL 5
A00404:156:HV37TDSXX:2:1438:26747:30091 chr21 18690550 N chr21 18690697 N DEL 5
A00404:156:HV37TDSXX:4:2476:27724:31782 chr21 18690437 N chr21 18690730 N DEL 5
A00297:158:HT275DSXX:3:2421:20582:2159 chr21 18690391 N chr21 18690757 N DEL 23
A00404:155:HV27LDSXX:1:2502:31557:36135 chr21 18690625 N chr21 18690772 N DEL 20
A00297:158:HT275DSXX:2:1141:16098:26021 chr21 18690396 N chr21 18690762 N DEL 15
A00297:158:HT275DSXX:3:2650:12563:20494 chr21 18690514 N chr21 18690877 N DUP 6
A00404:155:HV27LDSXX:4:1506:22281:4633 chr21 18690514 N chr21 18690807 N DEL 4
A00404:155:HV27LDSXX:4:2654:1380:10457 chr21 18690742 N chr21 18690962 N DEL 15
A00404:156:HV37TDSXX:4:1333:23845:7028 chr1 23504431 N chr1 23504557 N DUP 2
A00404:155:HV27LDSXX:4:2678:7907:30592 chr1 23504431 N chr1 23504557 N DUP 3
A00404:155:HV27LDSXX:4:1306:21142:1564 chr1 23504431 N chr1 23504557 N DUP 4
A00297:158:HT275DSXX:4:2601:12653:34272 chr1 23504447 N chr1 23504573 N DUP 13
A00297:158:HT275DSXX:3:1611:3305:14074 chr1 23504447 N chr1 23504573 N DUP 15
A00297:158:HT275DSXX:1:1153:19244:25895 chr1 23504447 N chr1 23504573 N DUP 15
A00404:155:HV27LDSXX:1:1129:6135:29810 chr1 23504447 N chr1 23504573 N DUP 13
A00404:156:HV37TDSXX:2:1501:27199:3724 chrX 71741215 N chrX 71741272 N DEL 6
A00404:156:HV37TDSXX:2:1501:27272:3724 chrX 71741215 N chrX 71741272 N DEL 6
A00404:155:HV27LDSXX:3:1343:2844:1564 chrX 71741215 N chrX 71741272 N DEL 6
A00404:156:HV37TDSXX:3:1621:17734:1861 chrX 71741209 N chrX 71741318 N DUP 4
A00297:158:HT275DSXX:4:2419:32850:34554 chrX 71741209 N chrX 71741318 N DUP 5
A00404:156:HV37TDSXX:3:2245:7934:35806 chrX 71741209 N chrX 71741318 N DUP 8
A00404:156:HV37TDSXX:3:2245:8513:34147 chrX 71741209 N chrX 71741318 N DUP 8
A00297:158:HT275DSXX:4:1524:12463:27148 chrX 71741339 N chrX 71742012 N DEL 15
A00297:158:HT275DSXX:2:1135:10926:9361 chrX 71741160 N chrX 71741351 N DEL 5
A00404:155:HV27LDSXX:3:2307:13476:12430 chrX 71741374 N chrX 71742045 N DUP 10
A00404:156:HV37TDSXX:4:1365:4698:11882 chrX 71741366 N chrX 71741953 N DUP 7
A00297:158:HT275DSXX:4:1438:15420:4805 chrX 71741363 N chrX 71741948 N DUP 17
A00404:156:HV37TDSXX:1:2137:11234:15311 chrX 71741374 N chrX 71742017 N DUP 9
A00404:155:HV27LDSXX:2:2429:26702:17550 chrX 71741374 N chrX 71742017 N DUP 10
A00404:155:HV27LDSXX:3:1550:29514:4194 chrX 71741362 N chrX 71741949 N DUP 6
A00404:155:HV27LDSXX:1:1109:19524:24940 chrX 71741379 N chrX 71741966 N DUP 5
A00297:158:HT275DSXX:1:2270:2112:3615 chrX 71741967 N chrX 71742022 N DUP 5
A00297:158:HT275DSXX:1:1447:22010:29997 chr3 177271601 N chr3 177271762 N DEL 5
A00297:158:HT275DSXX:2:1603:6985:1438 chrX 122710639 N chrX 122710848 N DUP 10
A00297:158:HT275DSXX:2:1632:3812:31454 chr9 36482197 N chr9 36482501 N DUP 1
A00404:156:HV37TDSXX:4:1340:31584:12571 chr9 36482202 N chr9 36482502 N DUP 5
A00297:158:HT275DSXX:2:2340:31964:28573 chr9 36482211 N chr9 36482516 N DEL 2
A00404:156:HV37TDSXX:4:2455:31901:22701 chr9 36482211 N chr9 36482516 N DEL 2
A00404:156:HV37TDSXX:1:1278:6451:3208 chr9 36482211 N chr9 36482516 N DEL 2
A00404:156:HV37TDSXX:3:1378:12680:17190 chr20 57629519 N chr20 57629636 N DUP 6
A00404:156:HV37TDSXX:2:2423:23954:30796 chr20 57629492 N chr20 57629610 N DUP 5
A00404:156:HV37TDSXX:1:2410:31982:32174 chr20 57629492 N chr20 57629610 N DUP 5
A00297:158:HT275DSXX:1:1444:25500:20071 chr20 57629492 N chr20 57629610 N DUP 5
A00297:158:HT275DSXX:1:1445:25174:5791 chr20 57629492 N chr20 57629610 N DUP 5
A00297:158:HT275DSXX:3:2358:5819:35149 chr20 57629519 N chr20 57629636 N DUP 6
A00404:155:HV27LDSXX:4:1248:28791:14779 chr20 57629492 N chr20 57629610 N DUP 5
A00404:155:HV27LDSXX:1:2502:31421:1611 chr20 57629492 N chr20 57629610 N DUP 10
A00297:158:HT275DSXX:4:2521:16694:12774 chr20 57629492 N chr20 57629610 N DUP 10
A00297:158:HT275DSXX:4:2521:17707:13683 chr20 57629492 N chr20 57629610 N DUP 10
A00404:155:HV27LDSXX:2:2418:1307:5259 chr1 121875927 N chr1 121876262 N DUP 5
A00404:155:HV27LDSXX:2:1560:28284:5916 chr1 121875930 N chr1 121876265 N DUP 4
A00297:158:HT275DSXX:2:2262:13548:31156 chr1 121876030 N chr1 121876696 N DEL 5
A00297:158:HT275DSXX:3:1465:12337:22983 chr1 121876030 N chr1 121876696 N DEL 5
A00404:155:HV27LDSXX:2:2327:15736:23610 chr1 121875968 N chr1 121876803 N DUP 3
A00297:158:HT275DSXX:2:2443:17065:13667 chr1 121876030 N chr1 121876696 N DEL 5
A00404:155:HV27LDSXX:3:2421:19135:36855 chr4 68870559 N chr4 68870628 N DEL 8
A00404:156:HV37TDSXX:3:1406:30463:32111 chr4 68870522 N chr4 68870592 N DEL 10
A00404:155:HV27LDSXX:2:2243:31919:13307 chr4 53256009 N chr4 53256183 N DUP 5
A00404:155:HV27LDSXX:3:1144:17074:33724 chr4 53256009 N chr4 53256183 N DUP 5
A00404:155:HV27LDSXX:2:1550:7753:19930 chr4 53256062 N chr4 53256283 N DEL 27
A00404:156:HV37TDSXX:2:2238:19343:34741 chr2 41747894 N chr2 41748122 N DUP 2
A00404:156:HV37TDSXX:1:2345:6470:11381 chr2 41747816 N chr2 41747994 N DEL 7
A00297:158:HT275DSXX:1:2337:24930:11130 chr2 41747833 N chr2 41748064 N DEL 6
A00404:156:HV37TDSXX:2:2330:5882:20228 chr4 21247740 N chr4 21247900 N DUP 3
A00297:158:HT275DSXX:2:2447:10547:17691 chr4 21247738 N chr4 21247900 N DUP 5
A00404:155:HV27LDSXX:4:1307:32117:20040 chr4 21247754 N chr4 21247948 N DUP 5
A00404:155:HV27LDSXX:4:2307:29261:13119 chr4 21247754 N chr4 21247948 N DUP 5
A00297:158:HT275DSXX:2:2534:31801:34084 chr8 67461762 N chr8 67461890 N DEL 5
A00404:155:HV27LDSXX:4:1435:10710:31594 chr8 67461798 N chr8 67461926 N DEL 5
A00297:158:HT275DSXX:2:1644:9362:14982 chr3 112430487 N chr3 112430551 N DUP 5
A00297:158:HT275DSXX:4:1626:17300:14920 chr3 112430487 N chr3 112430551 N DUP 5
A00297:158:HT275DSXX:1:2271:8061:15546 chr10 36789766 N chr10 36789897 N DEL 2
A00404:155:HV27LDSXX:4:1659:30156:27790 chr10 124598906 N chr10 124598963 N DEL 10
A00404:155:HV27LDSXX:2:1474:4508:21981 chr8 142185888 N chr8 142186044 N DUP 13
A00404:155:HV27LDSXX:2:2163:29478:26897 chr12 9197926 N chr12 9197989 N DEL 12
A00297:158:HT275DSXX:4:1301:1199:15718 chr12 9197926 N chr12 9197989 N DEL 5
A00404:156:HV37TDSXX:4:1629:9317:32377 chr12 9197926 N chr12 9197989 N DEL 8
A00404:155:HV27LDSXX:2:2619:31566:8469 chr12 9197895 N chr12 9197989 N DEL 5
A00297:158:HT275DSXX:1:2114:7527:1157 chr12 9197864 N chr12 9197989 N DEL 5
A00297:158:HT275DSXX:3:2642:24813:35759 chr12 9197864 N chr12 9197989 N DEL 5
A00404:155:HV27LDSXX:3:1304:18864:8390 chr12 9197842 N chr12 9197998 N DEL 5
A00404:156:HV37TDSXX:1:2463:9896:19038 chr7 76172220 N chr7 76172529 N DEL 30
A00297:158:HT275DSXX:3:1175:12988:9267 chr3 91261061 N chr3 91261911 N DEL 2
A00404:155:HV27LDSXX:3:1266:24406:19648 chr3 91261061 N chr3 91261911 N DEL 2
A00404:156:HV37TDSXX:1:1121:8006:9001 chr3 91261227 N chr3 91262244 N DUP 13
A00404:155:HV27LDSXX:3:2215:28167:35055 chr3 91261285 N chr3 91261793 N DUP 5
A00404:155:HV27LDSXX:1:1641:12038:36432 chr3 91261162 N chr3 91261503 N DEL 5
A00404:156:HV37TDSXX:3:2271:21712:5525 chr3 91261162 N chr3 91261503 N DEL 5
A00297:158:HT275DSXX:3:1332:30065:13228 chr3 91261185 N chr3 91261693 N DUP 5
A00297:158:HT275DSXX:3:2160:24822:36996 chr3 91261208 N chr3 91261718 N DEL 2
A00404:156:HV37TDSXX:3:2437:2510:32049 chr3 91261009 N chr3 91261857 N DUP 8
A00404:156:HV37TDSXX:4:2129:6777:11224 chr3 91261112 N chr3 91261961 N DUP 8
A00297:158:HT275DSXX:1:2619:20283:28761 chr3 91261112 N chr3 91261961 N DUP 10
A00297:158:HT275DSXX:1:2619:20392:28260 chr3 91261112 N chr3 91261961 N DUP 10
A00404:155:HV27LDSXX:1:1641:12038:36432 chr3 91261198 N chr3 91262047 N DUP 5
A00404:156:HV37TDSXX:3:2271:21712:5525 chr3 91261198 N chr3 91262047 N DUP 5
A00404:155:HV27LDSXX:4:1662:23854:25676 chr3 91261779 N chr3 91262118 N DUP 5
A00297:158:HT275DSXX:3:1626:20518:9408 chr3 91261067 N chr3 91262087 N DEL 15
A00404:156:HV37TDSXX:4:2656:3341:20995 chr3 91261786 N chr3 91262127 N DEL 10
A00404:156:HV37TDSXX:1:1442:19705:4867 chr3 91261100 N chr3 91262121 N DEL 5
A00297:158:HT275DSXX:3:2178:27181:36573 chr3 91261806 N chr3 91262147 N DEL 5
A00404:156:HV37TDSXX:3:2562:27841:17613 chr3 91261809 N chr3 91262150 N DEL 5
A00404:156:HV37TDSXX:2:1535:19904:30264 chr3 91261318 N chr3 91262168 N DEL 6
A00404:156:HV37TDSXX:3:1166:27760:9706 chr3 91261318 N chr3 91262168 N DEL 5
A00404:155:HV27LDSXX:4:2247:11858:7122 chr16 34736501 N chr16 34736882 N DUP 10
A00404:155:HV27LDSXX:3:2510:22507:34522 chr8 143342250 N chr8 143342341 N DUP 3
A00404:156:HV37TDSXX:4:2642:6361:33927 chr8 143342227 N chr8 143342321 N DEL 11
A00404:155:HV27LDSXX:3:1332:15763:8406 chr11 41304194 N chr11 41304322 N DEL 2
A00404:156:HV37TDSXX:1:1510:32027:22169 chr11 41304120 N chr11 41304201 N DUP 2
A00297:158:HT275DSXX:1:1125:16125:31986 chr11 41304194 N chr11 41304371 N DEL 8
A00297:158:HT275DSXX:1:1125:16125:31986 chr11 41304194 N chr11 41304371 N DEL 10
A00404:156:HV37TDSXX:4:1656:32136:29215 chr11 41304231 N chr11 41304408 N DEL 1
A00404:156:HV37TDSXX:1:2676:3531:35853 chr11 41304303 N chr11 41304478 N DUP 1
A00297:158:HT275DSXX:1:2659:9426:31657 chr11 41304215 N chr11 41304343 N DEL 21
A00404:156:HV37TDSXX:4:2131:5294:32612 chr11 41304159 N chr11 41304335 N DEL 1
A00297:158:HT275DSXX:1:2477:11369:9659 chr11 41304215 N chr11 41304343 N DEL 10
A00404:156:HV37TDSXX:2:1668:3558:4586 chr11 41304163 N chr11 41304464 N DUP 5
A00297:158:HT275DSXX:3:1404:2600:17926 chr11 41304292 N chr11 41304516 N DUP 5
A00404:155:HV27LDSXX:1:2214:25102:32158 chr2 118973423 N chr2 118973491 N DUP 5
A00297:158:HT275DSXX:1:1418:21043:28823 chr18 13673855 N chr18 13674031 N DUP 2
A00404:155:HV27LDSXX:2:2504:16676:34538 chr18 13673901 N chr18 13674036 N DEL 9
A00404:155:HV27LDSXX:2:2619:16143:30514 chr18 13673967 N chr18 13674105 N DEL 11
A00297:158:HT275DSXX:4:1516:7545:13620 chr18 13673901 N chr18 13674036 N DEL 10
A00404:155:HV27LDSXX:3:2219:30590:24533 chr18 13673897 N chr18 13674122 N DUP 14
A00404:155:HV27LDSXX:1:2241:12852:21089 chr18 13673929 N chr18 13674020 N DUP 7
A00297:158:HT275DSXX:3:1438:5276:8688 chr18 13673929 N chr18 13674020 N DUP 7
A00297:158:HT275DSXX:3:2438:1244:16078 chr18 13673929 N chr18 13674020 N DUP 7
A00404:156:HV37TDSXX:2:2248:26829:11036 chr18 13674013 N chr18 13674105 N DEL 12
A00297:158:HT275DSXX:3:2218:7970:4711 chr5 99426191 N chr5 99426267 N DEL 5
A00404:156:HV37TDSXX:1:2451:17635:22545 chr5 99426191 N chr5 99426267 N DEL 7
A00297:158:HT275DSXX:1:2144:23854:35571 chr5 99426191 N chr5 99426267 N DEL 10
A00404:156:HV37TDSXX:3:1469:6451:2080 chr5 99426191 N chr5 99426267 N DEL 10
A00404:156:HV37TDSXX:2:2678:10963:5541 chr5 99426191 N chr5 99426267 N DEL 10
A00404:155:HV27LDSXX:3:2505:12355:7451 chr5 99426191 N chr5 99426267 N DEL 10
A00297:158:HT275DSXX:3:1229:19325:6558 chr5 99426191 N chr5 99426267 N DEL 10
A00297:158:HT275DSXX:3:1229:19407:6543 chr5 99426191 N chr5 99426267 N DEL 10
A00297:158:HT275DSXX:1:1636:6542:17581 chr5 99426191 N chr5 99426267 N DEL 10
A00297:158:HT275DSXX:4:2240:29939:8406 chr5 99426194 N chr5 99426270 N DEL 9
A00297:158:HT275DSXX:4:2240:30418:7921 chr5 99426192 N chr5 99426268 N DEL 10
A00297:158:HT275DSXX:2:2439:31295:3552 chr5 99426194 N chr5 99426270 N DEL 10
A00404:156:HV37TDSXX:1:1376:29758:15389 chr5 99426214 N chr5 99426386 N DUP 7
A00297:158:HT275DSXX:1:2144:23854:35571 chr5 99426214 N chr5 99426386 N DUP 7
A00404:156:HV37TDSXX:4:1528:2157:19727 chr5 99426201 N chr5 99426277 N DEL 5
A00297:158:HT275DSXX:3:2144:21486:11741 chr5 99426197 N chr5 99426273 N DEL 9
A00404:156:HV37TDSXX:1:2216:9905:4742 chr5 99426407 N chr5 99426889 N DEL 7
A00404:155:HV27LDSXX:1:1519:27905:22232 chr5 99426411 N chr5 99426464 N DEL 12
A00404:155:HV27LDSXX:1:2509:19741:30326 chr5 99426411 N chr5 99426464 N DEL 12
A00297:158:HT275DSXX:3:1602:24288:29622 chr5 99426208 N chr5 99426457 N DUP 5
A00404:156:HV37TDSXX:4:2447:5466:28870 chr5 99426210 N chr5 99426482 N DUP 5
A00297:158:HT275DSXX:2:1158:16884:20337 chr5 99426435 N chr5 99426486 N DUP 9
A00297:158:HT275DSXX:4:2465:22978:11287 chr5 99426332 N chr5 99426585 N DEL 16
A00404:155:HV27LDSXX:1:2622:8024:25880 chr5 99426488 N chr5 99426666 N DEL 15
A00404:156:HV37TDSXX:1:1561:8178:7733 chr5 99426488 N chr5 99426666 N DEL 17
A00404:156:HV37TDSXX:1:2676:17083:12446 chr5 99426488 N chr5 99426666 N DEL 17
A00297:158:HT275DSXX:4:1272:10664:4554 chr5 99426488 N chr5 99426666 N DEL 19
A00404:155:HV27LDSXX:1:1256:12409:29559 chr5 99426232 N chr5 99426585 N DEL 14
A00404:156:HV37TDSXX:2:1350:11876:23312 chr5 99426488 N chr5 99426666 N DEL 32
A00404:155:HV27LDSXX:4:1318:8847:30655 chr5 99426517 N chr5 99426668 N DEL 23
A00297:158:HT275DSXX:2:2171:15971:24236 chr5 99426488 N chr5 99426641 N DEL 24
A00404:155:HV27LDSXX:3:1147:31105:6136 chr5 99426537 N chr5 99426769 N DUP 19
A00404:156:HV37TDSXX:2:2131:26277:9925 chr5 99426537 N chr5 99426769 N DUP 14
A00404:156:HV37TDSXX:2:1572:27588:3709 chr5 99426459 N chr5 99426566 N DEL 9
A00404:156:HV37TDSXX:3:1437:7880:1955 chr5 99426465 N chr5 99426566 N DEL 13
A00297:158:HT275DSXX:2:2650:23303:20870 chr5 99426524 N chr5 99426577 N DEL 2
A00297:158:HT275DSXX:1:1124:8169:1861 chr5 99426525 N chr5 99426578 N DEL 1
A00297:158:HT275DSXX:1:1124:8359:2033 chr5 99426525 N chr5 99426578 N DEL 1
A00297:158:HT275DSXX:4:1272:10664:4554 chr5 99426670 N chr5 99426954 N DEL 2
A00404:155:HV27LDSXX:3:1147:31105:6136 chr5 99426684 N chr5 99426862 N DEL 4
A00297:158:HT275DSXX:1:2351:29713:30436 chr5 99426520 N chr5 99426719 N DUP 11
A00297:158:HT275DSXX:3:2574:3857:23328 chr5 99426520 N chr5 99426719 N DUP 11
A00404:155:HV27LDSXX:1:2509:19741:30326 chr5 99426711 N chr5 99426862 N DEL 5
A00404:155:HV27LDSXX:4:2676:12753:25113 chr5 99426907 N chr5 99426962 N DEL 9
A00404:155:HV27LDSXX:3:1201:16667:29324 chr5 99426448 N chr5 99426628 N DEL 3
A00404:155:HV27LDSXX:3:1201:16857:28714 chr5 99426448 N chr5 99426628 N DEL 3
A00404:155:HV27LDSXX:2:1534:24117:17613 chr5 99426517 N chr5 99426668 N DEL 23
A00297:158:HT275DSXX:2:2650:23303:20870 chr5 99426488 N chr5 99426641 N DEL 24
A00404:156:HV37TDSXX:2:1350:11876:23312 chr5 99426896 N chr5 99426951 N DEL 14
A00404:155:HV27LDSXX:3:1201:16667:29324 chr5 99426565 N chr5 99426951 N DEL 9
A00404:155:HV27LDSXX:3:1201:16857:28714 chr5 99426565 N chr5 99426951 N DEL 9
A00297:158:HT275DSXX:4:1220:11677:22623 chr5 99426572 N chr5 99426719 N DUP 11
A00404:155:HV27LDSXX:2:1419:23791:5055 chr5 99426738 N chr5 99426862 N DEL 14
A00404:155:HV27LDSXX:3:2505:12355:7451 chr5 99426572 N chr5 99426719 N DUP 11
A00297:158:HT275DSXX:1:2129:32172:14121 chr5 99426542 N chr5 99426668 N DEL 12
A00404:156:HV37TDSXX:2:1676:16369:33692 chr5 99426572 N chr5 99426719 N DUP 11
A00404:156:HV37TDSXX:1:2149:8278:25817 chr5 99426572 N chr5 99426719 N DUP 11
A00404:155:HV27LDSXX:3:2374:9019:25379 chr5 99426542 N chr5 99426668 N DEL 15
A00404:155:HV27LDSXX:4:1124:32000:33270 chr5 99426658 N chr5 99426711 N DUP 12
A00297:158:HT275DSXX:3:1469:28257:19836 chr5 99426572 N chr5 99426719 N DUP 11
A00297:158:HT275DSXX:3:2468:27471:28902 chr5 99426572 N chr5 99426719 N DUP 11
A00404:156:HV37TDSXX:2:1409:32687:13448 chr5 99426572 N chr5 99426719 N DUP 11
A00404:155:HV27LDSXX:3:2302:31684:12117 chr5 99426465 N chr5 99426566 N DEL 14
A00404:156:HV37TDSXX:4:2140:13512:32189 chr5 99426537 N chr5 99426769 N DUP 18
A00297:158:HT275DSXX:3:1101:22923:16423 chr5 99426537 N chr5 99426769 N DUP 18
A00404:156:HV37TDSXX:2:1244:27028:14074 chr5 99426572 N chr5 99426719 N DUP 11
A00404:155:HV27LDSXX:2:2177:7970:20494 chr5 99426537 N chr5 99426769 N DUP 18
A00404:155:HV27LDSXX:3:1423:4291:31626 chr5 99426537 N chr5 99426769 N DUP 18
A00404:155:HV27LDSXX:3:2423:2754:31313 chr5 99426537 N chr5 99426769 N DUP 18
A00404:156:HV37TDSXX:1:1502:15374:18098 chr5 99426572 N chr5 99426719 N DUP 14
A00404:155:HV27LDSXX:3:2642:32425:4977 chr5 99426572 N chr5 99426719 N DUP 12
A00297:158:HT275DSXX:1:2173:9372:11459 chr5 99426459 N chr5 99426564 N DEL 9
A00404:155:HV27LDSXX:4:1276:22137:12524 chr5 99426459 N chr5 99426564 N DEL 8
A00297:158:HT275DSXX:3:1229:19325:6558 chr5 99426459 N chr5 99426564 N DEL 5
A00404:155:HV27LDSXX:1:1429:2917:10207 chr5 99426459 N chr5 99426564 N DEL 5
A00404:155:HV27LDSXX:2:1472:2880:12023 chr5 99426656 N chr5 99426836 N DEL 5
A00404:156:HV37TDSXX:2:1327:10981:6230 chr5 99426459 N chr5 99426564 N DEL 5
A00297:158:HT275DSXX:1:1321:32127:26725 chr5 99426459 N chr5 99426564 N DEL 5
A00404:156:HV37TDSXX:4:1257:21097:18615 chr5 99426459 N chr5 99426564 N DEL 5
A00404:155:HV27LDSXX:2:1617:27606:18333 chr5 99426460 N chr5 99426565 N DEL 5
A00404:156:HV37TDSXX:3:2206:3839:21198 chr5 99426656 N chr5 99426836 N DEL 5
A00297:158:HT275DSXX:3:1560:22571:36793 chr5 99426656 N chr5 99426836 N DEL 5
A00404:156:HV37TDSXX:4:2211:22299:27774 chr5 99426656 N chr5 99426836 N DEL 5
A00404:155:HV27LDSXX:2:2203:18674:18082 chr5 99426896 N chr5 99426951 N DEL 14
A00404:155:HV27LDSXX:4:1351:7048:32800 chr5 99426738 N chr5 99426862 N DEL 4
A00404:156:HV37TDSXX:1:1163:18493:32550 chr5 99426896 N chr5 99426951 N DEL 14
A00404:156:HV37TDSXX:1:1163:18683:32628 chr5 99426896 N chr5 99426951 N DEL 9
A00404:156:HV37TDSXX:1:2149:8278:25817 chr5 99426897 N chr5 99426950 N DEL 15
A00404:155:HV27LDSXX:2:2203:19054:17394 chr5 99426896 N chr5 99426951 N DEL 14
A00404:155:HV27LDSXX:4:1537:14986:14168 chr5 99426897 N chr5 99426950 N DEL 18
A00404:156:HV37TDSXX:2:1647:14244:21809 chr5 99426897 N chr5 99426950 N DEL 17
A00404:156:HV37TDSXX:2:1647:14687:21762 chr5 99426897 N chr5 99426950 N DEL 17
A00297:158:HT275DSXX:2:2316:28194:24236 chr5 99426897 N chr5 99426950 N DEL 17
A00404:155:HV27LDSXX:3:2417:29071:4304 chr5 99426904 N chr5 99426957 N DEL 5
A00297:158:HT275DSXX:3:2468:27471:28902 chr5 99426705 N chr5 99426962 N DEL 3
A00404:156:HV37TDSXX:4:1630:16179:25410 chr5 99426464 N chr5 99426950 N DEL 6
A00297:158:HT275DSXX:3:2102:3613:8594 chr5 99426464 N chr5 99426950 N DEL 6
A00297:158:HT275DSXX:3:2102:3739:7717 chr5 99426464 N chr5 99426950 N DEL 6
A00404:156:HV37TDSXX:2:1113:27181:5102 chr5 99426464 N chr5 99426950 N DEL 7
A00404:156:HV37TDSXX:1:2421:29369:12649 chr5 99426464 N chr5 99426950 N DEL 5
A00297:158:HT275DSXX:1:1124:16071:28917 chr5 99426691 N chr5 99427027 N DUP 4
A00404:156:HV37TDSXX:4:2140:13512:32189 chr5 99426691 N chr5 99427027 N DUP 5
A00297:158:HT275DSXX:1:1275:21856:13510 chr5 99426904 N chr5 99426957 N DEL 5
A00297:158:HT275DSXX:3:1469:28257:19836 chr5 99426705 N chr5 99426962 N DEL 3
A00404:155:HV27LDSXX:1:1519:27905:22232 chr5 99426464 N chr5 99426950 N DEL 5
A00404:155:HV27LDSXX:3:1423:4291:31626 chr5 99426862 N chr5 99427075 N DUP 2
A00404:155:HV27LDSXX:3:2423:2754:31313 chr5 99426862 N chr5 99427075 N DUP 2
A00404:155:HV27LDSXX:2:2209:19994:25473 chr5 99426862 N chr5 99427075 N DUP 2
A00297:158:HT275DSXX:2:2430:28637:31548 chr5 99426902 N chr5 99426955 N DEL 5
A00404:156:HV37TDSXX:4:1614:20012:19899 chr5 99426464 N chr5 99427031 N DEL 5
A00404:156:HV37TDSXX:4:1257:21097:18615 chr5 99426902 N chr5 99427036 N DEL 5
A00297:158:HT275DSXX:1:1264:23095:3004 chr5 99426903 N chr5 99427064 N DEL 5
A00404:156:HV37TDSXX:1:1502:15374:18098 chr5 99426705 N chr5 99427070 N DEL 3
A00404:156:HV37TDSXX:3:1167:17264:8719 chr5 99426706 N chr5 99427071 N DEL 2
A00404:156:HV37TDSXX:2:1244:27028:14074 chr5 99426464 N chr5 99427085 N DEL 5
A00404:156:HV37TDSXX:4:2421:22064:15029 chr5 99426707 N chr5 99427099 N DEL 1
A00297:158:HT275DSXX:3:1101:22923:16423 chr5 99426464 N chr5 99427112 N DEL 5
A00404:155:HV27LDSXX:3:1466:9001:21089 chr5 99426904 N chr5 99427119 N DEL 5
A00404:155:HV27LDSXX:4:1508:7139:1235 chr5 99426897 N chr5 99427139 N DEL 5
A00404:156:HV37TDSXX:3:1232:31720:5666 chr5 99426464 N chr5 99427139 N DEL 5
A00404:155:HV27LDSXX:2:1217:5900:2378 chr5 99426466 N chr5 99427141 N DEL 5
A00404:156:HV37TDSXX:2:2407:26449:21089 chr5 99426900 N chr5 99427142 N DEL 5
A00404:155:HV27LDSXX:2:1617:27606:18333 chr5 99426904 N chr5 99427146 N DEL 5
A00297:158:HT275DSXX:3:2157:29351:15937 chr14 20506571 N chr14 20506747 N DUP 5
A00404:156:HV37TDSXX:4:2415:31765:27539 chr14 20506427 N chr14 20506603 N DUP 5
A00404:155:HV27LDSXX:4:1469:9191:17848 chr14 20506571 N chr14 20506747 N DUP 5
A00297:158:HT275DSXX:4:1669:1895:22122 chr14 20506570 N chr14 20507071 N DEL 5
A00297:158:HT275DSXX:4:1669:1895:22122 chr14 20506683 N chr14 20507007 N DEL 5
A00297:158:HT275DSXX:4:1307:1805:6089 chr14 20506500 N chr14 20506805 N DEL 4
A00297:158:HT275DSXX:2:2669:15727:12038 chr14 20506461 N chr14 20506816 N DEL 3
A00297:158:HT275DSXX:4:1227:5077:1767 chr14 20506463 N chr14 20506817 N DEL 9
A00297:158:HT275DSXX:4:2217:30255:5854 chr14 20506468 N chr14 20506870 N DEL 7
A00297:158:HT275DSXX:4:2465:32723:15233 chr14 20506815 N chr14 20506913 N DUP 7
A00297:158:HT275DSXX:1:2424:24026:10128 chr14 20506978 N chr14 20507057 N DEL 2
A00297:158:HT275DSXX:3:2119:1380:12148 chr14 20506456 N chr14 20506811 N DEL 6
A00297:158:HT275DSXX:2:2233:3848:10723 chr14 20506586 N chr14 20506861 N DEL 5
A00297:158:HT275DSXX:3:2539:1551:17801 chr14 20506462 N chr14 20506961 N DUP 5
A00404:155:HV27LDSXX:2:2549:7844:20369 chr14 20506567 N chr14 20506891 N DEL 4
A00404:156:HV37TDSXX:2:2528:6126:4867 chr14 20506570 N chr14 20506894 N DEL 13
A00404:156:HV37TDSXX:4:2445:30789:19742 chr14 20506669 N chr14 20506992 N DUP 17
A00404:155:HV27LDSXX:4:1563:18909:3020 chr14 20506982 N chr14 20507160 N DEL 9
A00297:158:HT275DSXX:4:2409:15013:29872 chr14 20506496 N chr14 20506995 N DUP 4
A00404:155:HV27LDSXX:4:1511:9543:10880 chr14 20506442 N chr14 20507069 N DUP 4
A00404:156:HV37TDSXX:4:2550:4797:27680 chr14 20506491 N chr14 20506992 N DEL 5
A00297:158:HT275DSXX:3:1616:4589:25222 chr14 20506835 N chr14 20507060 N DUP 5
A00297:158:HT275DSXX:4:1177:2781:25316 chr14 20506459 N chr14 20507135 N DUP 10
A00297:158:HT275DSXX:2:1639:31611:33285 chr14 20506560 N chr14 20507061 N DEL 5
A00297:158:HT275DSXX:3:1616:4589:25222 chr14 20506983 N chr14 20507159 N DUP 5
A00404:155:HV27LDSXX:4:2171:18313:21151 chr14 20506467 N chr14 20507096 N DEL 8
A00297:158:HT275DSXX:3:1456:1045:30984 chr14 20506873 N chr14 20507100 N DEL 4
A00404:156:HV37TDSXX:2:1353:10113:30968 chr14 20506446 N chr14 20507174 N DEL 5
A00404:156:HV37TDSXX:4:2468:19732:22451 chr6 18565684 N chr6 18566294 N DEL 5
A00297:158:HT275DSXX:4:1375:8269:13119 chr6 18565684 N chr6 18566294 N DEL 5
A00404:155:HV27LDSXX:1:1462:25852:7529 chr6 18565722 N chr6 18566187 N DEL 5
A00404:155:HV27LDSXX:3:1374:31620:2832 chr6 18565796 N chr6 18565849 N DEL 1
A00297:158:HT275DSXX:2:1430:30418:18129 chr6 18566081 N chr6 18566189 N DEL 2
A00404:155:HV27LDSXX:1:1453:29252:10661 chr6 18566277 N chr6 18566385 N DUP 5
A00404:155:HV27LDSXX:1:1259:8097:30890 chr5 80361387 N chr5 80361454 N DEL 9
A00297:158:HT275DSXX:3:2608:10312:29089 chr10 477632 N chr10 477775 N DEL 4
A00297:158:HT275DSXX:3:2608:9751:29465 chr10 477632 N chr10 477775 N DEL 4
A00404:155:HV27LDSXX:2:1310:19967:2409 chr1 8851229 N chr1 8851327 N DEL 1
A00404:156:HV37TDSXX:4:2248:19633:37027 chr18 77343514 N chr18 77343605 N DEL 5
A00404:156:HV37TDSXX:4:1452:23122:30890 chr18 77343514 N chr18 77343605 N DEL 16
A00404:156:HV37TDSXX:4:1127:8838:11851 chrX 2225372 N chrX 2225570 N DEL 13
A00297:158:HT275DSXX:3:2436:8006:29042 chrX 2225226 N chrX 2225322 N DEL 7
A00404:155:HV27LDSXX:4:1124:12156:2910 chrX 2225226 N chrX 2225322 N DEL 7
A00297:158:HT275DSXX:3:2409:23845:9659 chr6 169376868 N chr6 169377149 N DEL 1
A00297:158:HT275DSXX:3:2409:24731:9659 chr6 169376868 N chr6 169377149 N DEL 1
A00404:155:HV27LDSXX:1:2609:12888:8531 chr6 169376868 N chr6 169377149 N DEL 5
A00297:158:HT275DSXX:1:2656:22028:5916 chr6 169376868 N chr6 169377149 N DEL 5
A00297:158:HT275DSXX:1:1432:2519:6574 chr6 169376840 N chr6 169376933 N DEL 35
A00404:156:HV37TDSXX:2:2244:12572:19225 chr6 169376868 N chr6 169377149 N DEL 5
A00404:155:HV27LDSXX:2:2628:32850:10629 chr6 169376856 N chr6 169377137 N DEL 5
A00297:158:HT275DSXX:1:1202:28203:18270 chr6 169376868 N chr6 169377149 N DEL 5
A00297:158:HT275DSXX:1:1209:19795:21339 chr6 169376868 N chr6 169377149 N DEL 5
A00297:158:HT275DSXX:1:2201:24469:16376 chr6 169376868 N chr6 169377149 N DEL 5
A00404:155:HV27LDSXX:1:2617:27489:22106 chr6 169376868 N chr6 169377149 N DEL 5
A00404:156:HV37TDSXX:1:2218:10502:24721 chr6 169376868 N chr6 169377149 N DEL 5
A00297:158:HT275DSXX:1:2309:20320:14231 chr6 169376868 N chr6 169377149 N DEL 2
A00404:156:HV37TDSXX:4:1315:2003:32612 chr6 169376878 N chr6 169377110 N DUP 15
A00297:158:HT275DSXX:3:2166:20464:5838 chr6 169377063 N chr6 169377765 N DEL 5
A00297:158:HT275DSXX:4:2636:23213:16830 chr6 169376868 N chr6 169377149 N DEL 10
A00404:155:HV27LDSXX:2:1610:28203:31892 chr6 169376868 N chr6 169377149 N DEL 10
A00404:155:HV27LDSXX:1:1332:5358:9956 chr6 169376868 N chr6 169377149 N DEL 10
A00404:155:HV27LDSXX:1:2552:9344:34710 chr6 169376868 N chr6 169377149 N DEL 10
A00404:155:HV27LDSXX:2:2468:12825:11960 chr6 169376868 N chr6 169377149 N DEL 10
A00404:156:HV37TDSXX:1:2238:31955:23578 chr6 169376868 N chr6 169377149 N DEL 10
A00404:156:HV37TDSXX:2:1522:26142:15483 chr6 169376868 N chr6 169377149 N DEL 10
A00404:155:HV27LDSXX:4:1629:6126:35869 chr6 169376871 N chr6 169377152 N DEL 5
A00404:155:HV27LDSXX:4:1630:6054:1485 chr6 169376871 N chr6 169377152 N DEL 5
A00297:158:HT275DSXX:3:1166:10655:27993 chr6 169376879 N chr6 169377160 N DEL 2
A00404:156:HV37TDSXX:4:1105:3622:11052 chr6 169376875 N chr6 169377203 N DEL 10
A00404:156:HV37TDSXX:1:2450:28058:1830 chr6 169376878 N chr6 169377251 N DUP 10
A00404:155:HV27LDSXX:2:1340:7292:12179 chr6 169376878 N chr6 169377251 N DUP 10
A00297:158:HT275DSXX:3:1629:1099:18928 chr6 169376903 N chr6 169377231 N DEL 10
A00404:155:HV27LDSXX:1:1575:16559:31829 chr6 169376903 N chr6 169377231 N DEL 6
A00404:155:HV27LDSXX:3:2521:18728:35775 chr6 169376903 N chr6 169377231 N DEL 6
A00297:158:HT275DSXX:1:2457:18756:15937 chr6 169376878 N chr6 169377251 N DUP 10
A00297:158:HT275DSXX:2:1139:32316:2284 chr6 169376878 N chr6 169377251 N DUP 10
A00404:156:HV37TDSXX:3:1175:29812:21966 chr6 169376878 N chr6 169377251 N DUP 10
A00297:158:HT275DSXX:3:1246:9200:5838 chr6 169377347 N chr6 169377769 N DEL 4
A00404:155:HV27LDSXX:2:1507:31268:19288 chr6 169376926 N chr6 169377301 N DEL 5
A00297:158:HT275DSXX:4:2571:4363:22545 chr6 169377031 N chr6 169377171 N DUP 5
A00404:155:HV27LDSXX:1:1612:6424:10958 chr6 169377065 N chr6 169377160 N DEL 10
A00297:158:HT275DSXX:3:2328:31367:13354 chr6 169376831 N chr6 169377159 N DEL 14
A00297:158:HT275DSXX:3:1246:9200:5838 chr6 169376878 N chr6 169377251 N DUP 10
A00404:156:HV37TDSXX:2:1211:4734:25598 chr6 169377002 N chr6 169377751 N DEL 5
A00297:158:HT275DSXX:3:1223:28176:29371 chr6 169376869 N chr6 169377804 N DEL 30
A00297:158:HT275DSXX:3:2511:7319:32299 chr6 169377129 N chr6 169377831 N DEL 23
A00404:156:HV37TDSXX:3:2647:22959:17738 chr4 46265562 N chr4 46265640 N DEL 9
A00404:155:HV27LDSXX:4:2174:24768:16611 chr4 46265562 N chr4 46265640 N DEL 9
A00404:156:HV37TDSXX:4:2141:31006:3333 chr4 46265562 N chr4 46265640 N DEL 9
A00404:155:HV27LDSXX:4:1352:4435:25927 chr3 94930354 N chr3 94930405 N DEL 5
A00404:155:HV27LDSXX:1:2257:4860:3458 chr3 94930354 N chr3 94930405 N DEL 5
A00404:155:HV27LDSXX:1:1552:14579:28620 chr3 94930354 N chr3 94930405 N DEL 5
A00404:156:HV37TDSXX:1:1508:14199:32628 chr3 94930329 N chr3 94930405 N DEL 5
A00404:156:HV37TDSXX:4:1171:22299:5791 chr3 94930329 N chr3 94930405 N DEL 5
A00297:158:HT275DSXX:2:1206:26087:29731 chr3 94930308 N chr3 94930409 N DEL 5
A00297:158:HT275DSXX:2:1526:12644:26303 chr1 195722690 N chr1 195722851 N DEL 5
A00404:155:HV27LDSXX:2:1365:16233:13260 chr1 160134223 N chr1 160134378 N DEL 8
A00297:158:HT275DSXX:3:1130:26657:31000 chr1 160134235 N chr1 160134438 N DEL 5
A00297:158:HT275DSXX:4:1326:29993:3991 chr5 176558486 N chr5 176558656 N DEL 34
A00404:156:HV37TDSXX:1:1559:19596:26443 chr5 176558514 N chr5 176558681 N DUP 5
A00404:156:HV37TDSXX:4:1452:15447:27054 chr5 176558528 N chr5 176558697 N DEL 5
A00297:158:HT275DSXX:4:1326:29993:3991 chr5 176558534 N chr5 176558703 N DEL 2
A00297:158:HT275DSXX:4:2168:27932:35869 chr7 61062974 N chr7 61063091 N DUP 3
A00297:158:HT275DSXX:1:1127:2184:30608 chr7 61062972 N chr7 61063089 N DUP 5
A00297:158:HT275DSXX:3:2324:29288:17394 chr7 61062905 N chr7 61062975 N DEL 2
A00404:155:HV27LDSXX:2:1421:20654:1971 chr7 61062974 N chr7 61063091 N DUP 3
A00404:155:HV27LDSXX:2:1173:15302:27148 chr7 61062984 N chr7 61063101 N DUP 5
A00404:156:HV37TDSXX:4:2252:30400:32377 chr7 61062984 N chr7 61063101 N DUP 5
A00404:156:HV37TDSXX:4:2607:20573:3364 chr17 32521822 N chr17 32521957 N DEL 13
A00404:156:HV37TDSXX:4:2607:20573:3364 chr17 32521823 N chr17 32521958 N DEL 8
A00404:156:HV37TDSXX:2:2536:29640:2848 chr1 1596583 N chr1 1596780 N DEL 3
A00404:155:HV27LDSXX:2:2169:29098:18098 chr1 1596583 N chr1 1596780 N DEL 4
A00404:155:HV27LDSXX:1:1409:1823:20556 chr1 1596583 N chr1 1596780 N DEL 5
A00404:155:HV27LDSXX:2:2403:12798:24377 chr1 1596583 N chr1 1596780 N DEL 5
A00404:155:HV27LDSXX:4:1234:27986:5274 chr1 1596605 N chr1 1596800 N DUP 5
A00404:155:HV27LDSXX:3:2143:12066:11866 chr1 1596606 N chr1 1596801 N DUP 5
A00404:155:HV27LDSXX:4:1172:28944:13135 chr1 1596495 N chr1 1596608 N DEL 5
A00297:158:HT275DSXX:3:2216:25048:8202 chr1 1596530 N chr1 1596737 N DUP 7
A00404:155:HV27LDSXX:2:2169:29098:18098 chr1 1596497 N chr1 1596744 N DEL 7
A00297:158:HT275DSXX:2:1634:10375:16924 chr1 1596501 N chr1 1596748 N DEL 7
A00297:158:HT275DSXX:1:2625:2853:18302 chr13 113371540 N chr13 113371957 N DEL 1
A00297:158:HT275DSXX:1:2625:3323:18615 chr13 113371540 N chr13 113371957 N DEL 1
A00404:156:HV37TDSXX:2:2326:17318:28447 chr13 113371540 N chr13 113371957 N DEL 1
A00297:158:HT275DSXX:4:1342:28718:34538 chr13 113371600 N chr13 113371840 N DEL 1
A00297:158:HT275DSXX:1:2153:22381:19272 chr13 113371540 N chr13 113371957 N DEL 5
A00297:158:HT275DSXX:1:1669:14778:36918 chr13 113371540 N chr13 113371957 N DEL 5
A00297:158:HT275DSXX:1:1605:10339:35806 chr13 113371570 N chr13 113371630 N DEL 7
A00404:156:HV37TDSXX:2:2175:16224:31093 chr13 113371570 N chr13 113371810 N DEL 10
A00404:155:HV27LDSXX:3:2123:12563:2926 chr13 113371570 N chr13 113371790 N DEL 27
A00297:158:HT275DSXX:4:2110:14425:27946 chr13 113371570 N chr13 113371790 N DEL 33
A00404:155:HV27LDSXX:3:1627:19587:5979 chr13 113371578 N chr13 113371798 N DEL 33
A00404:155:HV27LDSXX:1:1211:13792:1673 chr13 113371570 N chr13 113371790 N DEL 30
A00404:155:HV27LDSXX:1:2149:32208:19038 chr13 113371987 N chr13 113372046 N DUP 22
A00404:156:HV37TDSXX:2:2144:1244:31767 chr13 113371542 N chr13 113371660 N DUP 18
A00297:158:HT275DSXX:2:2223:6741:16141 chr13 113371649 N chr13 113372063 N DUP 16
A00297:158:HT275DSXX:2:2221:18566:28698 chr13 113371542 N chr13 113371660 N DUP 23
A00297:158:HT275DSXX:1:1204:30092:23703 chr13 113371615 N chr13 113371950 N DUP 14
A00404:156:HV37TDSXX:1:2359:30960:12148 chr13 113371668 N chr13 113371965 N DEL 15
A00404:156:HV37TDSXX:4:1548:19985:23265 chr13 113371541 N chr13 113371898 N DUP 23
A00297:158:HT275DSXX:3:2609:5746:34366 chr13 113371648 N chr13 113372063 N DUP 5
A00404:155:HV27LDSXX:1:2672:3522:29105 chr13 113371614 N chr13 113371691 N DUP 11
A00404:156:HV37TDSXX:2:2551:20681:27915 chr13 113371808 N chr13 113371945 N DUP 11
A00404:155:HV27LDSXX:2:2517:3477:11898 chr13 113371542 N chr13 113371660 N DUP 24
A00404:156:HV37TDSXX:1:2265:16613:11976 chr13 113371831 N chr13 113371951 N DUP 17
A00297:158:HT275DSXX:2:2451:12924:6840 chr13 113371890 N chr13 113371970 N DUP 17
A00297:158:HT275DSXX:2:1309:24180:28307 chr13 113371542 N chr13 113371899 N DUP 23
A00404:155:HV27LDSXX:2:1339:25409:31031 chr13 113371651 N chr13 113371729 N DUP 4
A00404:156:HV37TDSXX:2:2122:25012:7044 chr13 113371542 N chr13 113371899 N DUP 23
A00404:155:HV27LDSXX:1:2622:24243:37059 chr13 113371542 N chr13 113371601 N DUP 18
A00404:155:HV27LDSXX:1:1575:9805:17566 chr13 113371604 N chr13 113371980 N DEL 16
A00404:156:HV37TDSXX:3:1574:19623:19100 chr13 113371604 N chr13 113371980 N DEL 16
A00404:156:HV37TDSXX:3:2670:30355:5932 chr13 113371580 N chr13 113371976 N DEL 5
A00404:155:HV27LDSXX:2:1425:14335:23782 chr13 113371567 N chr13 113372005 N DEL 5
A00404:156:HV37TDSXX:4:2177:19235:2738 chr13 113371676 N chr13 113372014 N DEL 5
A00297:158:HT275DSXX:3:1650:8992:10958 chr13 113371677 N chr13 113372015 N DEL 5
A00404:155:HV27LDSXX:4:1158:6198:18458 chr13 113371965 N chr13 113372046 N DEL 3
A00297:158:HT275DSXX:2:1549:2672:22936 chr10 30677445 N chr10 30677578 N DUP 7
A00404:155:HV27LDSXX:2:1222:5674:32049 chr10 30677555 N chr10 30677932 N DUP 14
A00297:158:HT275DSXX:1:1425:30861:16141 chr10 30677624 N chr10 30677826 N DEL 27
A00297:158:HT275DSXX:3:2648:14823:32487 chr10 30677624 N chr10 30677826 N DEL 22
A00404:155:HV27LDSXX:1:2168:31286:13714 chr10 30677555 N chr10 30677932 N DUP 14
A00297:158:HT275DSXX:4:2146:23204:10927 chr10 30677685 N chr10 30677930 N DUP 13
A00404:155:HV27LDSXX:4:1111:3875:36605 chr10 30677674 N chr10 30677919 N DUP 8
A00297:158:HT275DSXX:3:1426:18168:33332 chr10 30677553 N chr10 30677930 N DUP 14
A00404:155:HV27LDSXX:2:2344:28519:16595 chr10 30677710 N chr10 30677867 N DUP 5
A00297:158:HT275DSXX:4:1411:4273:17910 chr10 30677447 N chr10 30677870 N DUP 1
A00404:156:HV37TDSXX:4:2335:30816:7169 chr10 30677779 N chr10 30677871 N DEL 14
A00297:158:HT275DSXX:2:2309:32479:17754 chr10 30677841 N chr10 30677909 N DEL 9
A00404:156:HV37TDSXX:1:2577:8838:18834 chr10 30677470 N chr10 30677917 N DEL 5
A00404:155:HV27LDSXX:4:2517:16902:15796 chr10 30677466 N chr10 30677913 N DEL 5
A00404:156:HV37TDSXX:2:1133:14353:8406 chr10 30677429 N chr10 30677921 N DEL 3
A00404:156:HV37TDSXX:2:1133:14407:9032 chr10 30677429 N chr10 30677921 N DEL 3
A00404:156:HV37TDSXX:2:1341:24596:13777 chr10 30677469 N chr10 30677938 N DEL 5
A00404:155:HV27LDSXX:2:1134:14696:22561 chr10 30677469 N chr10 30677938 N DEL 5
A00404:155:HV27LDSXX:1:1256:7645:21966 chr10 30677428 N chr10 30677942 N DEL 1
A00297:158:HT275DSXX:3:2212:15347:11819 chr14 104527031 N chr14 104527204 N DUP 9
A00297:158:HT275DSXX:3:2538:19623:36479 chr14 104527031 N chr14 104527204 N DUP 9
A00404:156:HV37TDSXX:4:2617:11867:9173 chr14 104527047 N chr14 104527226 N DEL 1
A00297:158:HT275DSXX:4:1142:16360:16266 chr14 104527086 N chr14 104527251 N DEL 9
A00404:155:HV27LDSXX:3:2634:3604:6010 chr14 104527254 N chr14 104527351 N DUP 8
A00404:155:HV27LDSXX:4:2304:14678:28291 chr19 4163852 N chr19 4164313 N DUP 1
A00297:158:HT275DSXX:2:1203:28619:14325 chr19 4163852 N chr19 4164313 N DUP 1
A00297:158:HT275DSXX:3:1302:15826:1939 chr15 74968159 N chr15 74968341 N DEL 5
A00404:156:HV37TDSXX:2:1515:11632:8484 chr15 74968148 N chr15 74968330 N DEL 18
A00404:156:HV37TDSXX:1:2322:17372:1830 chr15 74968194 N chr15 74968376 N DEL 45
A00404:156:HV37TDSXX:1:2322:17372:1830 chr15 74968194 N chr15 74968376 N DEL 58
A00297:158:HT275DSXX:1:2535:5032:8015 chr5 144865642 N chr5 144865989 N DUP 5
A00404:156:HV37TDSXX:1:2214:16568:34976 chr5 144865642 N chr5 144865989 N DUP 5
A00404:155:HV27LDSXX:4:1371:15564:13479 chr5 144865642 N chr5 144865989 N DUP 5
A00404:156:HV37TDSXX:4:2253:12445:12242 chr5 144865642 N chr5 144865989 N DUP 5
A00404:155:HV27LDSXX:1:2405:20039:22013 chr5 144865642 N chr5 144865989 N DUP 5
A00404:155:HV27LDSXX:4:2678:13386:36667 chr5 144865661 N chr5 144866010 N DEL 5
A00404:156:HV37TDSXX:4:1174:1398:27242 chr5 144865666 N chr5 144866015 N DEL 4
A00404:156:HV37TDSXX:2:2154:16993:2550 chr2 241472296 N chr2 241473193 N DEL 1
A00404:155:HV27LDSXX:3:2405:6162:4022 chr2 241472372 N chr2 241472664 N DEL 12
A00404:155:HV27LDSXX:2:2674:20374:11945 chr2 241472305 N chr2 241472712 N DEL 5
A00404:156:HV37TDSXX:3:1574:31711:35430 chr16 86884201 N chr16 86884284 N DUP 1
A00404:156:HV37TDSXX:1:2138:25102:32503 chr16 86884201 N chr16 86884284 N DUP 2
A00297:158:HT275DSXX:1:1209:4246:26475 chr16 86884284 N chr16 86884384 N DEL 10
A00404:156:HV37TDSXX:1:1411:18674:5462 chr16 86884284 N chr16 86884384 N DEL 12
A00404:156:HV37TDSXX:3:2563:9507:10629 chr16 86884334 N chr16 86884417 N DEL 12
A00404:155:HV27LDSXX:1:1568:9986:13714 chr16 86884334 N chr16 86884417 N DEL 43
A00297:158:HT275DSXX:1:2152:22290:7874 chr16 86884334 N chr16 86884417 N DEL 25
A00297:158:HT275DSXX:2:2365:19714:17378 chr16 86884334 N chr16 86884417 N DEL 30
A00297:158:HT275DSXX:3:1429:27028:21590 chr16 86884334 N chr16 86884417 N DEL 26
A00297:158:HT275DSXX:1:2152:22299:7545 chr16 86884334 N chr16 86884417 N DEL 34
A00404:155:HV27LDSXX:3:1514:30996:28714 chr16 86884334 N chr16 86884417 N DEL 24
A00404:155:HV27LDSXX:3:2544:24623:14794 chr16 86884279 N chr16 86884363 N DEL 3
A00404:156:HV37TDSXX:1:1266:20410:30545 chr16 86884334 N chr16 86884417 N DEL 18
A00404:156:HV37TDSXX:3:2307:15980:4335 chr16 86884238 N chr16 86884422 N DEL 5
A00404:156:HV37TDSXX:1:1470:26133:32847 chr16 86884239 N chr16 86884423 N DEL 5
A00404:156:HV37TDSXX:1:1470:28772:33755 chr16 86884239 N chr16 86884423 N DEL 5
A00404:155:HV27LDSXX:4:1334:7039:7200 chr16 86884240 N chr16 86884424 N DEL 5
A00404:156:HV37TDSXX:4:2244:17083:13886 chr16 86884193 N chr16 86884427 N DEL 5
A00404:155:HV27LDSXX:3:2526:16315:26396 chr17 80274755 N chr17 80274886 N DEL 10
A00404:155:HV27LDSXX:2:1557:31937:23077 chr7 82999628 N chr7 82999757 N DEL 5
A00297:158:HT275DSXX:2:1538:11523:29935 chr7 82999628 N chr7 82999757 N DEL 9
A00404:156:HV37TDSXX:2:1160:8287:13495 chr7 82999628 N chr7 82999757 N DEL 12
A00404:155:HV27LDSXX:1:1154:9453:33270 chr7 82999628 N chr7 82999757 N DEL 12
A00404:155:HV27LDSXX:2:1219:12518:19727 chr7 82999640 N chr7 82999693 N DEL 5
A00297:158:HT275DSXX:4:2207:28149:11130 chr7 82999771 N chr7 82999837 N DEL 25
A00404:156:HV37TDSXX:1:1510:27037:28463 chr7 82999771 N chr7 82999837 N DEL 25
A00404:156:HV37TDSXX:1:1510:27199:33254 chr7 82999771 N chr7 82999837 N DEL 25
A00297:158:HT275DSXX:4:2449:13422:17221 chr7 82999769 N chr7 82999861 N DEL 24
A00404:156:HV37TDSXX:4:1167:23529:9142 chr7 82999771 N chr7 82999837 N DEL 19
A00297:158:HT275DSXX:2:1443:26747:30029 chr7 82999837 N chr7 82999992 N DUP 14
A00404:156:HV37TDSXX:4:1505:32127:23782 chr7 82999772 N chr7 82999838 N DEL 9
A00404:156:HV37TDSXX:3:2141:5873:13855 chr7 82999880 N chr7 82999957 N DUP 15
A00404:155:HV27LDSXX:2:1346:8350:36808 chr7 82999880 N chr7 82999957 N DUP 14
A00404:155:HV27LDSXX:3:2546:32633:3145 chr7 82999769 N chr7 82999861 N DEL 7
A00404:155:HV27LDSXX:3:2203:6569:18724 chr7 82999880 N chr7 82999931 N DUP 10
A00404:156:HV37TDSXX:4:2468:14850:29559 chr7 82999880 N chr7 82999957 N DUP 10
A00404:155:HV27LDSXX:3:1110:4535:36808 chr7 82999880 N chr7 82999957 N DUP 12
A00404:156:HV37TDSXX:2:1564:6126:24815 chr7 82999880 N chr7 82999957 N DUP 12
A00297:158:HT275DSXX:2:1277:16966:24079 chr7 82999880 N chr7 82999957 N DUP 15
A00404:156:HV37TDSXX:2:1253:3902:24251 chr7 82999956 N chr7 83000007 N DEL 14
A00297:158:HT275DSXX:4:2314:9715:28494 chr7 82999938 N chr7 83000041 N DEL 14
A00404:155:HV27LDSXX:2:2345:19108:9846 chr7 82999938 N chr7 83000041 N DEL 14
A00404:155:HV27LDSXX:3:1461:1298:2738 chr7 82999938 N chr7 83000041 N DEL 14
A00404:155:HV27LDSXX:2:1630:28366:20650 chr7 82999938 N chr7 83000041 N DEL 14
A00297:158:HT275DSXX:2:2237:9127:12915 chr7 82999912 N chr7 83000041 N DEL 5
A00297:158:HT275DSXX:2:1207:2663:32878 chr7 82999912 N chr7 83000041 N DEL 5
A00404:155:HV27LDSXX:2:1454:27552:35900 chr7 82999912 N chr7 83000041 N DEL 5
A00404:156:HV37TDSXX:2:1253:3902:24251 chr7 82999912 N chr7 83000041 N DEL 5
A00404:155:HV27LDSXX:1:1215:19877:14779 chr7 82999763 N chr7 83000042 N DEL 5
A00404:155:HV27LDSXX:1:1603:29288:22373 chr7 82999614 N chr7 83000049 N DEL 5
A00404:156:HV37TDSXX:4:1457:18873:25254 chr7 82999614 N chr7 83000049 N DEL 5
A00404:155:HV27LDSXX:1:2160:13458:9267 chr19 7229122 N chr19 7229478 N DEL 4
A00404:156:HV37TDSXX:4:2330:29496:21605 chr19 7229122 N chr19 7229478 N DEL 5
A00404:155:HV27LDSXX:1:1353:17183:15812 chr19 7229130 N chr19 7229482 N DEL 6
A00404:155:HV27LDSXX:1:2353:16884:2581 chr19 7229130 N chr19 7229482 N DEL 6
A00404:156:HV37TDSXX:2:2644:29125:2738 chr19 7229130 N chr19 7229482 N DEL 13
A00297:158:HT275DSXX:3:1518:2058:17895 chr19 7229345 N chr19 7229451 N DEL 4
A00297:158:HT275DSXX:2:1650:2365:34240 chr19 7229144 N chr19 7229452 N DEL 12
A00297:158:HT275DSXX:3:1611:25644:26897 chr19 7229418 N chr19 7229486 N DEL 8
A00404:155:HV27LDSXX:1:2547:24849:17848 chr19 7229145 N chr19 7229493 N DEL 4
A00297:158:HT275DSXX:1:1547:6207:20259 chr6 143649046 N chr6 143649105 N DUP 8
A00404:156:HV37TDSXX:2:1505:29695:13119 chr3 95784086 N chr3 95784237 N DEL 16
A00297:158:HT275DSXX:4:2665:6361:7247 chr3 95784086 N chr3 95784237 N DEL 16
A00297:158:HT275DSXX:1:1531:18674:1517 chr3 95784110 N chr3 95784193 N DUP 24
A00404:156:HV37TDSXX:4:2671:24876:14512 chr3 95784110 N chr3 95784193 N DUP 29
A00404:156:HV37TDSXX:2:1214:14172:27602 chr3 95784110 N chr3 95784262 N DUP 18
A00404:155:HV27LDSXX:2:1213:24668:18944 chr3 95784138 N chr3 95784193 N DUP 16
A00297:158:HT275DSXX:1:1238:13602:3067 chr3 95784110 N chr3 95784262 N DUP 27
A00404:156:HV37TDSXX:1:2621:29197:13228 chr3 95784138 N chr3 95784193 N DUP 16
A00297:158:HT275DSXX:4:1341:26711:25113 chr3 95784110 N chr3 95784193 N DUP 21
A00297:158:HT275DSXX:1:1531:18674:1517 chr3 95784110 N chr3 95784193 N DUP 21
A00297:158:HT275DSXX:4:2645:28583:19711 chr3 95784136 N chr3 95784232 N DUP 11
A00297:158:HT275DSXX:3:1135:18629:9079 chr3 95784136 N chr3 95784232 N DUP 11
A00404:156:HV37TDSXX:4:1547:30960:11021 chr3 95784136 N chr3 95784232 N DUP 16
A00297:158:HT275DSXX:1:1251:29423:22169 chr3 95784138 N chr3 95784262 N DUP 25
A00404:156:HV37TDSXX:4:1222:18132:20400 chr3 95784087 N chr3 95784311 N DUP 4
A00297:158:HT275DSXX:1:2364:16495:21981 chr3 95784087 N chr3 95784136 N DUP 25
A00297:158:HT275DSXX:1:2364:16694:22138 chr3 95784087 N chr3 95784136 N DUP 25
A00404:155:HV27LDSXX:3:2405:20871:30812 chr3 95784135 N chr3 95784238 N DEL 7
A00404:155:HV27LDSXX:2:2572:5168:7435 chr3 95784088 N chr3 95784360 N DUP 7
A00297:158:HT275DSXX:2:1514:19931:14810 chr3 95784086 N chr3 95784335 N DUP 5
A00404:155:HV27LDSXX:2:1125:28718:32784 chr3 95784134 N chr3 95784355 N DUP 5
A00404:156:HV37TDSXX:1:2670:1570:27414 chr3 95784087 N chr3 95784311 N DUP 11
A00404:155:HV27LDSXX:1:2403:7581:35008 chr3 95784094 N chr3 95784220 N DEL 7
A00404:156:HV37TDSXX:4:1222:17770:20400 chr3 95784087 N chr3 95784311 N DUP 4
A00404:155:HV27LDSXX:4:1174:4155:7028 chr3 95784087 N chr3 95784286 N DUP 12
A00404:155:HV27LDSXX:4:1461:3821:20478 chr3 95784135 N chr3 95784238 N DEL 7
A00297:158:HT275DSXX:1:1237:25201:16329 chr3 95784238 N chr3 95784310 N DUP 7
A00404:156:HV37TDSXX:4:1522:11876:21465 chr3 95784088 N chr3 95784335 N DUP 7
A00404:155:HV27LDSXX:1:2404:10131:7545 chr3 95784097 N chr3 95784223 N DEL 7
A00297:158:HT275DSXX:2:1127:4065:26036 chr3 95784087 N chr3 95784311 N DUP 11
A00297:158:HT275DSXX:1:2448:6958:15828 chr3 95784296 N chr3 95784349 N DEL 7
A00297:158:HT275DSXX:3:1135:18629:9079 chr3 95784352 N chr3 95784424 N DUP 7
A00404:156:HV37TDSXX:3:2355:6352:33849 chr3 95784357 N chr3 95784429 N DUP 7
A00404:155:HV27LDSXX:4:1224:7410:10974 chr3 95784447 N chr3 95784496 N DUP 31
A00297:158:HT275DSXX:4:1341:26711:25113 chr3 95784399 N chr3 95784521 N DUP 14
A00297:158:HT275DSXX:1:1238:13602:3067 chr3 95784447 N chr3 95784496 N DUP 29
A00404:156:HV37TDSXX:4:1561:13621:18317 chr3 95784447 N chr3 95784496 N DUP 21
A00404:156:HV37TDSXX:1:2177:30861:27007 chr9 20973087 N chr9 20973402 N DEL 5
A00404:155:HV27LDSXX:4:2476:15718:36605 chr9 20973087 N chr9 20973402 N DEL 5
A00404:156:HV37TDSXX:1:1355:19804:14559 chr9 20973087 N chr9 20973402 N DEL 5
A00404:155:HV27LDSXX:3:1369:27525:5729 chr9 20973087 N chr9 20973402 N DEL 5
A00404:155:HV27LDSXX:4:2513:14895:12038 chr9 20973087 N chr9 20973402 N DEL 5
A00297:158:HT275DSXX:2:2336:9607:36605 chr9 20973087 N chr9 20973402 N DEL 5
A00404:156:HV37TDSXX:4:1450:4851:17534 chr9 20973087 N chr9 20973402 N DEL 5
A00404:155:HV27LDSXX:2:2364:9796:17832 chr9 20973105 N chr9 20973312 N DUP 5
A00404:155:HV27LDSXX:4:2574:31539:17910 chr9 20973108 N chr9 20973315 N DUP 5
A00297:158:HT275DSXX:1:1620:32117:7513 chr9 20973200 N chr9 20973410 N DEL 5
A00297:158:HT275DSXX:1:1503:9977:18959 chr9 77761943 N chr9 77762169 N DEL 6
A00404:155:HV27LDSXX:2:2368:4110:12868 chr9 77762081 N chr9 77762384 N DEL 4
A00404:156:HV37TDSXX:2:1375:19135:31219 chr9 77761980 N chr9 77762301 N DUP 1
A00297:158:HT275DSXX:1:1503:9977:18959 chr9 77762012 N chr9 77762235 N DUP 3
A00404:155:HV27LDSXX:3:2607:20039:35509 chr9 77762011 N chr9 77762234 N DUP 3
A00404:155:HV27LDSXX:3:2203:13783:2597 chr9 77761906 N chr9 77762035 N DEL 5
A00404:155:HV27LDSXX:2:1515:1298:2112 chr9 77762184 N chr9 77762282 N DEL 5
A00297:158:HT275DSXX:1:1661:18566:23500 chr9 77761999 N chr9 77762098 N DEL 5
A00404:155:HV27LDSXX:4:1578:17870:13432 chr9 77762118 N chr9 77762468 N DUP 1
A00404:155:HV27LDSXX:1:2255:4345:15123 chr9 77761998 N chr9 77762221 N DUP 5
A00404:156:HV37TDSXX:1:1518:5385:35900 chr9 77761933 N chr9 77762159 N DEL 5
A00297:158:HT275DSXX:1:2361:1976:26083 chr9 77762243 N chr9 77762370 N DEL 4
A00404:155:HV27LDSXX:1:1544:5159:27179 chr9 77762049 N chr9 77762224 N DUP 9
A00404:155:HV27LDSXX:3:2653:26232:6183 chr9 77761999 N chr9 77762222 N DUP 5
A00297:158:HT275DSXX:3:2221:19361:28604 chr9 77762271 N chr9 77762448 N DEL 15
A00404:155:HV27LDSXX:4:2664:24162:27993 chr9 77762063 N chr9 77762288 N DEL 5
A00404:155:HV27LDSXX:4:1110:23140:1830 chr9 77762271 N chr9 77762397 N DUP 10
A00404:156:HV37TDSXX:3:1609:19226:35070 chr9 77762045 N chr9 77762395 N DUP 5
A00404:156:HV37TDSXX:4:2628:29523:9064 chr9 77761902 N chr9 77762303 N DEL 5
A00297:158:HT275DSXX:3:2221:19361:28604 chr9 77762271 N chr9 77762448 N DEL 21
A00404:155:HV27LDSXX:3:2577:9977:22310 chr9 77761993 N chr9 77762394 N DEL 5
A00297:158:HT275DSXX:2:2630:32108:32769 chr9 77762070 N chr9 77762422 N DEL 6
A00297:158:HT275DSXX:4:1555:27552:19053 chr9 77762433 N chr9 77762608 N DUP 5
A00297:158:HT275DSXX:3:1402:12472:34710 chr9 77761973 N chr9 77762550 N DEL 5
A00404:156:HV37TDSXX:3:2372:2456:24283 chr9 77762134 N chr9 77762660 N DUP 5
A00297:158:HT275DSXX:2:2623:7591:34898 chr9 77762287 N chr9 77762415 N DEL 11
A00404:156:HV37TDSXX:2:2451:25726:20181 chr9 77762324 N chr9 77762536 N DUP 2
A00404:155:HV27LDSXX:1:1311:7374:4116 chr9 77761902 N chr9 77762655 N DEL 4
A00404:155:HV27LDSXX:1:1578:26060:24017 chr19 55147494 N chr19 55147568 N DEL 10
A00404:156:HV37TDSXX:2:2427:27163:3975 chr19 55147494 N chr19 55147568 N DEL 21
A00297:158:HT275DSXX:4:2173:17806:31986 chr19 55147494 N chr19 55147568 N DEL 21
A00404:156:HV37TDSXX:2:1405:6659:28651 chr19 55147494 N chr19 55147568 N DEL 22
A00404:156:HV37TDSXX:2:1405:6858:27993 chr19 55147494 N chr19 55147568 N DEL 22
A00404:156:HV37TDSXX:3:2547:11198:5509 chr19 55147494 N chr19 55147568 N DEL 26
A00404:155:HV27LDSXX:4:2103:25997:33051 chr19 55147494 N chr19 55147568 N DEL 31
A00297:158:HT275DSXX:2:1657:29080:15718 chr19 55147494 N chr19 55147568 N DEL 26
A00404:156:HV37TDSXX:2:2649:16134:19100 chr19 55147494 N chr19 55147568 N DEL 26
A00404:156:HV37TDSXX:4:1474:24704:7044 chr19 55147494 N chr19 55147568 N DEL 22
A00297:158:HT275DSXX:1:2140:27263:25911 chr19 55147494 N chr19 55147568 N DEL 20
A00297:158:HT275DSXX:1:1662:24704:7357 chr19 55147494 N chr19 55147568 N DEL 20
A00404:156:HV37TDSXX:4:1314:22643:28181 chr19 55147404 N chr19 55147565 N DEL 4
A00404:156:HV37TDSXX:4:1421:7961:36761 chr19 55147494 N chr19 55147568 N DEL 8
A00404:155:HV27LDSXX:1:1413:30843:25723 chr19 55147802 N chr19 55147876 N DEL 5
A00297:158:HT275DSXX:3:2472:19741:35243 chr19 55147802 N chr19 55147876 N DEL 20
A00404:155:HV27LDSXX:3:2163:22182:25567 chr19 55147680 N chr19 55147836 N DEL 21
A00404:156:HV37TDSXX:4:2437:8766:28134 chr19 55147415 N chr19 55147839 N DEL 7
A00404:155:HV27LDSXX:4:2131:15185:19867 chr19 55147532 N chr19 55148015 N DUP 3
A00404:155:HV27LDSXX:1:1538:27046:3865 chr19 55380417 N chr19 55380555 N DEL 13
A00404:155:HV27LDSXX:1:2369:25644:10645 chr22 47810008 N chr22 47810310 N DUP 15
A00297:158:HT275DSXX:2:1259:10004:36260 chr22 47810156 N chr22 47810237 N DEL 5
A00404:155:HV27LDSXX:4:2159:19732:21480 chr22 47810156 N chr22 47810237 N DEL 5
A00404:156:HV37TDSXX:1:1157:30382:13620 chr22 47810156 N chr22 47810237 N DEL 5
A00297:158:HT275DSXX:2:2352:3170:8985 chr22 47810156 N chr22 47810237 N DEL 5
A00404:156:HV37TDSXX:4:1628:5918:3818 chr22 47810141 N chr22 47810298 N DEL 25
A00404:156:HV37TDSXX:2:1134:21115:20776 chr22 47810122 N chr22 47810177 N DUP 24
A00404:156:HV37TDSXX:2:1245:26802:20384 chr22 47810157 N chr22 47810251 N DUP 22
A00404:155:HV27LDSXX:1:2469:13792:1830 chr22 47810176 N chr22 47810268 N DUP 12
A00297:158:HT275DSXX:2:1570:31232:7106 chr22 47810024 N chr22 47810193 N DUP 2
A00404:155:HV27LDSXX:3:1420:4978:21292 chr22 47810040 N chr22 47810110 N DEL 12
A00404:155:HV27LDSXX:3:1420:6840:22013 chr22 47810040 N chr22 47810110 N DEL 12
A00404:155:HV27LDSXX:4:2367:26883:6433 chr22 47810043 N chr22 47810215 N DUP 5
A00404:155:HV27LDSXX:4:1341:7600:33943 chr22 47810044 N chr22 47810216 N DUP 23
A00297:158:HT275DSXX:3:1151:10438:4820 chr22 47810043 N chr22 47810215 N DUP 22
A00404:155:HV27LDSXX:3:2419:23258:19225 chr22 47810043 N chr22 47810215 N DUP 23
A00404:155:HV27LDSXX:1:2409:31557:18255 chr22 47810157 N chr22 47810251 N DUP 18
A00404:156:HV37TDSXX:4:2217:25346:20525 chr22 47810157 N chr22 47810251 N DUP 17
A00404:155:HV27LDSXX:3:1368:16604:30592 chr22 47810160 N chr22 47810254 N DUP 12
A00297:158:HT275DSXX:1:2671:23140:2300 chr22 47810097 N chr22 47810324 N DEL 9
A00404:156:HV37TDSXX:2:2437:7437:23453 chr22 47810103 N chr22 47810330 N DEL 9
A00404:156:HV37TDSXX:4:2262:5999:31391 chr15 98162836 N chr15 98162891 N DEL 5
A00404:155:HV27LDSXX:2:1652:8784:6464 chr15 98162836 N chr15 98162891 N DEL 5
A00297:158:HT275DSXX:3:2217:10899:33082 chr15 98162836 N chr15 98162891 N DEL 5
A00404:155:HV27LDSXX:3:1340:26214:3020 chr15 98162836 N chr15 98162891 N DEL 5
A00404:155:HV27LDSXX:4:1114:12626:22106 chr15 98162836 N chr15 98162891 N DEL 5
A00404:156:HV37TDSXX:3:2211:28031:9580 chr15 98162836 N chr15 98162891 N DEL 5
A00404:156:HV37TDSXX:4:1506:22453:30044 chr15 98162836 N chr15 98162891 N DEL 5
A00297:158:HT275DSXX:2:2471:25400:3615 chr15 98162836 N chr15 98162891 N DEL 5
A00404:156:HV37TDSXX:4:1237:23927:3599 chr15 98162875 N chr15 98162928 N DUP 5
A00404:156:HV37TDSXX:3:2268:27127:28307 chr15 98162875 N chr15 98162928 N DUP 5
A00297:158:HT275DSXX:2:1413:28637:30044 chr15 98162875 N chr15 98162928 N DUP 5
A00404:155:HV27LDSXX:4:2317:6668:25441 chr15 98162875 N chr15 98162928 N DUP 5
A00404:155:HV27LDSXX:4:1537:25735:11021 chr15 98162875 N chr15 98162928 N DUP 5
A00297:158:HT275DSXX:3:2363:12825:13307 chr15 98162889 N chr15 98162942 N DUP 1
A00404:155:HV27LDSXX:4:1161:17002:11021 chr4 179604351 N chr4 179604483 N DUP 1
A00404:156:HV37TDSXX:3:2612:21875:29418 chr16 81413027 N chr16 81413164 N DEL 18
A00297:158:HT275DSXX:1:1261:17870:13902 chr4 2955124 N chr4 2955407 N DEL 7
A00297:158:HT275DSXX:1:1261:17870:13902 chr4 2955124 N chr4 2955407 N DEL 7
A00297:158:HT275DSXX:1:1440:6741:17080 chr4 2955386 N chr4 2955605 N DEL 9
A00404:155:HV27LDSXX:2:1413:24966:12383 chr4 2955152 N chr4 2955628 N DEL 7
A00404:156:HV37TDSXX:2:1354:23484:6934 chr4 2955437 N chr4 2955718 N DEL 14
A00297:158:HT275DSXX:1:1608:5448:35728 chr4 2955442 N chr4 2955723 N DEL 10
A00297:158:HT275DSXX:4:2213:30110:22138 chr2 60250412 N chr2 60250462 N DUP 3
A00297:158:HT275DSXX:4:1274:15176:7169 chr12 132470921 N chr12 132471072 N DUP 7
A00404:156:HV37TDSXX:1:1405:22770:35509 chr12 132471106 N chr12 132471161 N DEL 4
A00297:158:HT275DSXX:3:2323:28791:6198 chr20 24431066 N chr20 24431189 N DUP 5
A00404:156:HV37TDSXX:2:2565:22471:18208 chr21 34016644 N chr21 34016941 N DEL 30
A00404:156:HV37TDSXX:4:1526:2266:12837 chr21 34016732 N chr21 34017029 N DEL 20
A00297:158:HT275DSXX:4:1111:11632:32722 chr21 34016713 N chr21 34017010 N DEL 19
A00404:156:HV37TDSXX:3:2271:23656:30780 chr21 34016764 N chr21 34017061 N DEL 2
A00297:158:HT275DSXX:3:2407:11478:32643 chr11 429278 N chr11 429502 N DEL 8
A00297:158:HT275DSXX:1:2532:32136:32503 chr11 429301 N chr11 429460 N DUP 5
A00297:158:HT275DSXX:3:2260:20202:11303 chr11 429116 N chr11 429466 N DEL 2
A00404:156:HV37TDSXX:3:1419:29830:29418 chr11 429178 N chr11 429528 N DEL 11
A00404:155:HV27LDSXX:1:2137:30581:1125 chr2 543942 N chr2 544035 N DEL 20
A00404:155:HV27LDSXX:1:1330:21685:10582 chr2 543924 N chr2 544055 N DEL 7
A00404:155:HV27LDSXX:1:1330:21703:10582 chr2 543924 N chr2 544055 N DEL 7
A00297:158:HT275DSXX:1:2109:2320:27148 chr2 86942615 N chr2 86942672 N DEL 5
A00297:158:HT275DSXX:1:1161:17580:14559 chr2 86942615 N chr2 86942672 N DEL 2
A00404:155:HV27LDSXX:4:2647:1371:30859 chr2 86942615 N chr2 86942672 N DEL 13
A00404:155:HV27LDSXX:2:2434:18900:32471 chr2 86942520 N chr2 86942717 N DEL 5
A00404:155:HV27LDSXX:2:1258:19651:36996 chr2 86942501 N chr2 86942720 N DEL 7
A00404:156:HV37TDSXX:4:1671:17390:28072 chr2 86942611 N chr2 86942694 N DUP 22
A00297:158:HT275DSXX:3:1312:27353:14011 chr2 86942513 N chr2 86942626 N DEL 5
A00297:158:HT275DSXX:4:2172:16396:29888 chr2 86942514 N chr2 86942627 N DEL 4
A00404:156:HV37TDSXX:4:2373:12355:15186 chr2 86942516 N chr2 86942629 N DEL 2
A00404:155:HV27LDSXX:2:2316:30228:32925 chr2 86942628 N chr2 86942685 N DEL 2
A00297:158:HT275DSXX:1:1233:15465:15123 chr2 86942498 N chr2 86942692 N DEL 8
A00297:158:HT275DSXX:4:1215:9290:32737 chr2 86942504 N chr2 86942723 N DEL 8
A00297:158:HT275DSXX:3:2274:14118:31861 chr2 86942643 N chr2 86942728 N DEL 14
A00404:156:HV37TDSXX:2:2261:8006:32737 chr2 86942615 N chr2 86942672 N DEL 39
A00404:155:HV27LDSXX:2:1654:29387:2315 chr4 189898160 N chr4 189898213 N DEL 14
A00404:155:HV27LDSXX:3:2603:29848:12602 chr7 140763364 N chr7 140763464 N DEL 5
A00297:158:HT275DSXX:3:1158:22968:2566 chr7 140763364 N chr7 140763464 N DEL 11
A00404:156:HV37TDSXX:2:1518:12825:15562 chr7 140763282 N chr7 140763508 N DEL 17
A00297:158:HT275DSXX:2:1614:19506:23030 chr7 140763338 N chr7 140763565 N DEL 5
A00404:155:HV27LDSXX:2:2468:2763:10285 chr1 194303748 N chr1 194303817 N DUP 9
A00404:156:HV37TDSXX:2:2204:4996:15530 chr1 194303724 N chr1 194303797 N DUP 10
A00404:156:HV37TDSXX:3:2316:27425:13949 chr1 194303724 N chr1 194303797 N DUP 10
A00404:155:HV27LDSXX:2:1619:32479:9706 chr1 194303792 N chr1 194303983 N DEL 10
A00404:155:HV27LDSXX:2:1619:32570:8829 chr1 194303792 N chr1 194303983 N DEL 10
A00297:158:HT275DSXX:2:2114:8250:31469 chr1 194303724 N chr1 194303797 N DUP 10
A00404:156:HV37TDSXX:1:1258:11921:21010 chr1 194303724 N chr1 194303797 N DUP 10
A00404:155:HV27LDSXX:1:1658:1380:26303 chr1 194303792 N chr1 194303983 N DEL 10
A00404:155:HV27LDSXX:1:1658:1651:23140 chr1 194303792 N chr1 194303983 N DEL 10
A00404:156:HV37TDSXX:3:1526:11876:34773 chr1 194303724 N chr1 194303797 N DUP 10
A00297:158:HT275DSXX:3:1561:17418:27398 chr1 194303724 N chr1 194303797 N DUP 10
A00404:156:HV37TDSXX:2:2515:22652:14074 chr1 194303724 N chr1 194303797 N DUP 10
A00404:156:HV37TDSXX:3:2161:2374:5102 chr1 194303724 N chr1 194303834 N DUP 8
A00404:155:HV27LDSXX:2:2524:31946:28980 chr1 194303724 N chr1 194303797 N DUP 10
A00297:158:HT275DSXX:1:2331:3803:6355 chr1 194303783 N chr1 194303974 N DEL 15
A00297:158:HT275DSXX:2:1630:19714:18098 chr1 194303792 N chr1 194303983 N DEL 10
A00404:155:HV27LDSXX:4:2305:13449:13354 chr1 194303793 N chr1 194303863 N DUP 8
A00404:156:HV37TDSXX:3:2239:23755:35744 chr1 194303724 N chr1 194303797 N DUP 10
A00404:155:HV27LDSXX:2:2430:31114:25974 chr1 194303724 N chr1 194303834 N DUP 8
A00297:158:HT275DSXX:1:1654:4996:23610 chr1 194303829 N chr1 194303983 N DEL 9
A00297:158:HT275DSXX:3:1152:7509:30373 chr1 194303724 N chr1 194303834 N DUP 9
A00297:158:HT275DSXX:1:1221:22236:23719 chr1 194303821 N chr1 194303979 N DEL 19
A00297:158:HT275DSXX:2:1646:24108:21355 chr1 194303793 N chr1 194303863 N DUP 8
A00404:156:HV37TDSXX:2:1539:3432:18427 chr1 194303724 N chr1 194303797 N DUP 10
A00404:155:HV27LDSXX:1:2160:21287:15875 chr1 194303979 N chr1 194304052 N DUP 16
A00404:155:HV27LDSXX:1:2372:10755:27132 chr1 194303979 N chr1 194304085 N DUP 26
A00404:156:HV37TDSXX:3:2445:3179:21746 chr1 194303793 N chr1 194303863 N DUP 8
A00404:155:HV27LDSXX:1:2214:12391:25050 chr1 194303724 N chr1 194303797 N DUP 10
A00404:155:HV27LDSXX:4:2442:29595:12477 chr1 194303979 N chr1 194304085 N DUP 27
A00404:155:HV27LDSXX:2:2430:31114:25974 chr1 194303793 N chr1 194303863 N DUP 8
A00404:155:HV27LDSXX:4:1538:3423:14716 chr1 194303793 N chr1 194303863 N DUP 8
A00404:156:HV37TDSXX:2:1539:3432:18427 chr1 194303793 N chr1 194303863 N DUP 8
A00404:155:HV27LDSXX:3:1541:32117:17848 chr1 194303793 N chr1 194303863 N DUP 8
A00297:158:HT275DSXX:4:1123:15628:1251 chr1 194303793 N chr1 194303863 N DUP 8
A00404:155:HV27LDSXX:3:2275:32606:16438 chr1 194303793 N chr1 194303863 N DUP 8
A00404:155:HV27LDSXX:1:1420:28384:35305 chr1 194303724 N chr1 194303871 N DUP 6
A00404:156:HV37TDSXX:2:2427:3721:36808 chr1 194303724 N chr1 194303908 N DUP 6
A00404:155:HV27LDSXX:4:1337:7898:34679 chr1 194303724 N chr1 194303871 N DUP 8
A00404:156:HV37TDSXX:1:2509:28420:31485 chr1 194303748 N chr1 194303854 N DUP 14
A00297:158:HT275DSXX:1:2331:3803:6355 chr1 194303748 N chr1 194303854 N DUP 14
A00404:156:HV37TDSXX:4:1265:28194:8766 chr1 194303793 N chr1 194303863 N DUP 8
A00404:155:HV27LDSXX:4:1626:29044:34006 chr1 194303724 N chr1 194303871 N DUP 10
A00404:155:HV27LDSXX:1:1469:26431:3458 chr1 194303724 N chr1 194303871 N DUP 10
A00297:158:HT275DSXX:3:1517:26250:24972 chr1 194303724 N chr1 194303834 N DUP 10
A00297:158:HT275DSXX:3:2328:11143:29904 chr1 194303724 N chr1 194303871 N DUP 10
A00404:155:HV27LDSXX:1:2526:18891:37027 chr1 194303793 N chr1 194303863 N DUP 8
A00404:156:HV37TDSXX:3:2463:4372:5838 chr1 194303748 N chr1 194303891 N DUP 14
A00297:158:HT275DSXX:2:1538:7220:25958 chr1 194303748 N chr1 194303854 N DUP 14
A00404:155:HV27LDSXX:1:1665:26973:26256 chr1 194303793 N chr1 194303900 N DUP 8
A00404:156:HV37TDSXX:2:2261:27778:33880 chr1 194303748 N chr1 194303891 N DUP 14
A00404:156:HV37TDSXX:2:1525:23348:10050 chr1 194303724 N chr1 194303871 N DUP 10
A00297:158:HT275DSXX:4:2176:3703:13291 chr1 194303748 N chr1 194303891 N DUP 14
A00297:158:HT275DSXX:3:2152:13955:8719 chr1 194303724 N chr1 194303871 N DUP 10
A00404:156:HV37TDSXX:2:1321:7093:2378 chr1 194303793 N chr1 194303900 N DUP 8
A00297:158:HT275DSXX:4:2637:5484:21136 chr1 194303748 N chr1 194303928 N DUP 9
A00404:155:HV27LDSXX:1:1658:1380:26303 chr1 194303735 N chr1 194303882 N DUP 5
A00404:155:HV27LDSXX:1:1658:1651:23140 chr1 194303735 N chr1 194303882 N DUP 5
A00404:156:HV37TDSXX:1:1560:11695:26318 chr1 194303748 N chr1 194303928 N DUP 9
A00404:156:HV37TDSXX:4:1261:5122:8140 chr1 194303748 N chr1 194303928 N DUP 9
A00297:158:HT275DSXX:1:1338:24894:13291 chr1 194303735 N chr1 194303882 N DUP 5
A00404:156:HV37TDSXX:1:2138:15148:2143 chr1 194303748 N chr1 194303928 N DUP 12
A00404:156:HV37TDSXX:2:2472:21350:33583 chr1 194303735 N chr1 194303919 N DUP 2
A00297:158:HT275DSXX:2:2263:27154:18051 chr1 194303735 N chr1 194303882 N DUP 5
A00404:155:HV27LDSXX:3:2560:28185:6840 chr1 194303735 N chr1 194303882 N DUP 5
A00297:158:HT275DSXX:3:1220:13657:23202 chr1 194303724 N chr1 194303908 N DUP 9
A00297:158:HT275DSXX:4:2449:6940:33207 chr1 194303748 N chr1 194303928 N DUP 13
A00404:156:HV37TDSXX:3:1247:29460:12336 chr1 194303793 N chr1 194303863 N DUP 8
A00404:155:HV27LDSXX:3:1331:3839:23860 chr1 194303735 N chr1 194303919 N DUP 4
A00297:158:HT275DSXX:2:1646:24108:21355 chr1 194303724 N chr1 194303908 N DUP 7
A00297:158:HT275DSXX:3:2436:13530:30311 chr1 194303735 N chr1 194303919 N DUP 5
A00404:156:HV37TDSXX:4:2148:28085:21919 chr1 194303793 N chr1 194303900 N DUP 8
A00404:155:HV27LDSXX:3:2430:21558:17096 chr1 194303793 N chr1 194303900 N DUP 8
A00297:158:HT275DSXX:3:1431:25997:3928 chr1 194303783 N chr1 194303974 N DEL 16
A00404:155:HV27LDSXX:1:2526:18891:37027 chr1 194303820 N chr1 194303974 N DEL 15
A00404:156:HV37TDSXX:3:2333:19316:1877 chr1 194303820 N chr1 194303974 N DEL 15
A00297:158:HT275DSXX:2:2573:21133:36495 chr1 194303820 N chr1 194303974 N DEL 15
A00404:156:HV37TDSXX:1:1103:27507:35227 chr1 194303820 N chr1 194303974 N DEL 15
A00404:155:HV27LDSXX:2:1352:6994:3458 chr1 194303820 N chr1 194303974 N DEL 15
A00404:155:HV27LDSXX:1:1122:10664:1423 chr1 194303784 N chr1 194303933 N DEL 5
A00404:155:HV27LDSXX:3:2208:16803:34757 chr1 194303785 N chr1 194303980 N DEL 19
A00404:155:HV27LDSXX:4:2305:13449:13354 chr1 194303792 N chr1 194303983 N DEL 10
A00297:158:HT275DSXX:2:2114:8250:31469 chr1 194303954 N chr1 194304032 N DUP 15
A00404:156:HV37TDSXX:2:2120:24297:17174 chr1 194303954 N chr1 194304032 N DUP 15
A00404:156:HV37TDSXX:1:1622:30147:7326 chr1 194303954 N chr1 194304032 N DUP 15
A00297:158:HT275DSXX:2:1538:7220:25958 chr1 194303954 N chr1 194304032 N DUP 15
A00404:156:HV37TDSXX:2:2204:4996:15530 chr1 194303954 N chr1 194304032 N DUP 12
A00297:158:HT275DSXX:3:1164:21233:25676 chr1 194303784 N chr1 194303979 N DEL 24
A00297:158:HT275DSXX:2:1630:19714:18098 chr1 194303781 N chr1 194303974 N DEL 22
A00297:158:HT275DSXX:2:1501:19705:29669 chr1 194303784 N chr1 194303979 N DEL 22
A00404:156:HV37TDSXX:4:2106:19587:9424 chr1 194303784 N chr1 194303979 N DEL 21
A00297:158:HT275DSXX:3:2442:15971:1532 chr1 194303784 N chr1 194303979 N DEL 19
A00404:155:HV27LDSXX:1:1469:26431:3458 chr1 194303784 N chr1 194303979 N DEL 19
A00404:155:HV27LDSXX:1:1252:6325:13197 chr1 194303784 N chr1 194303979 N DEL 19
A00404:155:HV27LDSXX:1:1252:7509:26459 chr1 194303784 N chr1 194303979 N DEL 19
A00404:156:HV37TDSXX:2:2472:21350:33583 chr1 194303822 N chr1 194303980 N DEL 19
A00404:156:HV37TDSXX:3:1637:30517:26569 chr1 194303784 N chr1 194303979 N DEL 19
A00404:155:HV27LDSXX:4:1469:15591:1814 chr1 194303783 N chr1 194303974 N DEL 15
A00404:155:HV27LDSXX:4:1469:17698:11569 chr1 194303783 N chr1 194303974 N DEL 15
A00404:155:HV27LDSXX:2:2675:4842:1297 chr1 194303786 N chr1 194303981 N DEL 19
A00297:158:HT275DSXX:2:1647:15492:25003 chr1 194303783 N chr1 194303974 N DEL 15
A00297:158:HT275DSXX:3:2263:11270:29872 chr1 194303786 N chr1 194303981 N DEL 19
A00404:156:HV37TDSXX:1:2377:6632:14669 chr1 194303783 N chr1 194303974 N DEL 15
A00404:156:HV37TDSXX:1:1602:8621:6809 chr1 194303711 N chr1 194303980 N DEL 14
A00297:158:HT275DSXX:4:2637:5484:21136 chr1 194303754 N chr1 194303982 N DEL 7
A00297:158:HT275DSXX:2:2359:1289:5729 chrY 10683266 N chrY 10683402 N DEL 8
A00404:156:HV37TDSXX:3:2642:6705:10410 chrY 10683266 N chrY 10683402 N DEL 8
A00404:156:HV37TDSXX:3:2642:7184:10238 chrY 10683266 N chrY 10683402 N DEL 8
A00404:156:HV37TDSXX:1:2359:22128:14262 chrY 10683262 N chrY 10683403 N DEL 12
A00404:155:HV27LDSXX:2:2235:13774:31767 chrY 10683282 N chrY 10683418 N DEL 4
A00404:155:HV27LDSXX:4:1573:1723:28432 chrY 10683282 N chrY 10683418 N DEL 4
A00404:155:HV27LDSXX:1:1521:14443:15045 chrY 10683265 N chrY 10683406 N DEL 9
A00297:158:HT275DSXX:2:2631:20844:20744 chrY 10683251 N chrY 10683432 N DEL 2
A00297:158:HT275DSXX:3:1471:32859:30185 chrY 10683251 N chrY 10683432 N DEL 2
A00404:156:HV37TDSXX:1:1473:19587:1720 chr9 8892663 N chr9 8892838 N DUP 5
A00297:158:HT275DSXX:1:1116:23366:10614 chr1 22678742 N chr1 22679086 N DUP 5
A00404:155:HV27LDSXX:4:2166:11686:7294 chr1 22679317 N chr1 22679481 N DEL 2
A00404:156:HV37TDSXX:2:1442:19759:11663 chr1 22679317 N chr1 22679481 N DEL 2
A00404:156:HV37TDSXX:2:2633:21567:5181 chr1 22679317 N chr1 22679481 N DEL 9
A00404:156:HV37TDSXX:4:2656:29957:30201 chr1 22679316 N chr1 22679480 N DEL 14
A00404:155:HV27LDSXX:3:2530:24659:3521 chr1 22679317 N chr1 22679481 N DEL 9
A00297:158:HT275DSXX:4:1314:15383:26600 chr1 22679376 N chr1 22679538 N DUP 18
A00404:155:HV27LDSXX:1:1404:14398:7983 chr1 22679376 N chr1 22679538 N DUP 17
A00404:155:HV27LDSXX:3:2467:21016:2597 chr1 22679379 N chr1 22679541 N DUP 12
A00404:156:HV37TDSXX:3:1358:15076:16454 chr1 22679379 N chr1 22679541 N DUP 12
A00404:156:HV37TDSXX:3:2450:30337:7373 chr1 22679444 N chr1 22679614 N DEL 27
A00404:155:HV27LDSXX:1:2617:4119:34303 chr8 3651801 N chr8 3651871 N DEL 5
A00404:155:HV27LDSXX:3:1527:14443:20964 chr8 3651801 N chr8 3651871 N DEL 5
A00297:158:HT275DSXX:1:2631:27208:21151 chr17 41149643 N chr17 41149809 N DEL 5
A00404:155:HV27LDSXX:4:1209:22046:8735 chr17 41149643 N chr17 41149809 N DEL 5
A00404:156:HV37TDSXX:2:1565:12075:11725 chr17 41149643 N chr17 41149809 N DEL 5
A00404:155:HV27LDSXX:4:1361:3794:19053 chr17 41149673 N chr17 41149852 N DUP 30
A00404:156:HV37TDSXX:3:2169:23945:5603 chr17 41149673 N chr17 41149852 N DUP 30
A00404:156:HV37TDSXX:4:2247:10339:8625 chr17 41149673 N chr17 41149852 N DUP 29
A00404:155:HV27LDSXX:3:1543:23140:27195 chr17 41149673 N chr17 41149852 N DUP 27
A00404:155:HV27LDSXX:1:2361:18231:4194 chr17 41149678 N chr17 41149812 N DUP 10
A00404:155:HV27LDSXX:1:2362:18258:8625 chr17 41149678 N chr17 41149812 N DUP 10
A00404:156:HV37TDSXX:4:1543:5873:14481 chr17 41149676 N chr17 41149810 N DUP 12
A00404:156:HV37TDSXX:4:1140:31846:13651 chr17 41149675 N chr17 41149809 N DUP 13
A00404:156:HV37TDSXX:4:2533:9968:9706 chr17 41149615 N chr17 41149839 N DUP 2
A00404:155:HV27LDSXX:2:1150:17155:16329 chr17 41149615 N chr17 41149839 N DUP 5
A00404:155:HV27LDSXX:3:2333:15293:7216 chr17 41149635 N chr17 41149861 N DEL 5
A00297:158:HT275DSXX:1:2310:5041:23249 chr3 48056242 N chr3 48056618 N DEL 2
A00404:155:HV27LDSXX:3:1244:15709:28260 chr3 48056265 N chr3 48056362 N DEL 19
A00297:158:HT275DSXX:1:2358:2130:21339 chr3 48056281 N chr3 48056557 N DEL 5
A00404:156:HV37TDSXX:4:1644:18954:36605 chr3 48056258 N chr3 48056359 N DEL 1
A00404:156:HV37TDSXX:1:1640:19804:5228 chr3 48056432 N chr3 48056660 N DEL 5
A00404:156:HV37TDSXX:2:2110:27814:5040 chr3 48056290 N chr3 48056389 N DEL 5
A00404:155:HV27LDSXX:4:2469:16170:23422 chr3 48056506 N chr3 48056557 N DEL 6
A00404:155:HV27LDSXX:2:2152:4246:32268 chr3 48056446 N chr3 48056523 N DUP 5
A00404:155:HV27LDSXX:3:2450:31241:12540 chr3 48056556 N chr3 48056656 N DEL 8
A00404:155:HV27LDSXX:2:2358:11605:26224 chr3 48056587 N chr3 48056638 N DEL 15
A00297:158:HT275DSXX:2:2606:15935:33004 chr3 48056397 N chr3 48056573 N DUP 5
A00404:156:HV37TDSXX:2:1221:15673:21057 chr3 48056519 N chr3 48056617 N DUP 9
A00404:156:HV37TDSXX:2:1636:10059:4100 chr3 48056415 N chr3 48056641 N DUP 8
A00404:156:HV37TDSXX:3:2575:11776:22576 chr3 48056369 N chr3 48056646 N DEL 6
A00404:156:HV37TDSXX:1:2261:9634:9345 chr2 161836634 N chr2 161836773 N DEL 2
A00404:156:HV37TDSXX:3:2347:16007:31313 chr2 161836634 N chr2 161836773 N DEL 2
A00404:155:HV27LDSXX:3:2256:8431:19445 chr2 161836637 N chr2 161836767 N DEL 5
A00404:156:HV37TDSXX:1:2131:3540:34147 chr2 47502684 N chr2 47502791 N DUP 11
A00404:155:HV27LDSXX:3:1515:13467:23907 chr2 47502689 N chr2 47502780 N DUP 8
A00297:158:HT275DSXX:4:2472:22489:31673 chr2 47502587 N chr2 47502816 N DEL 3
A00404:156:HV37TDSXX:3:2157:11433:8672 chr8 2475319 N chr8 2475389 N DEL 13
A00404:155:HV27LDSXX:3:1524:16658:36072 chr8 3385047 N chr8 3385187 N DEL 3
A00404:156:HV37TDSXX:3:2554:30346:16376 chr2 57455606 N chr2 57455665 N DUP 10
A00404:156:HV37TDSXX:3:2554:30517:16642 chr2 57455606 N chr2 57455665 N DUP 10
A00297:158:HT275DSXX:3:1533:8522:18067 chr2 57455606 N chr2 57455665 N DUP 10
A00297:158:HT275DSXX:1:1623:31232:27085 chr2 57455606 N chr2 57455695 N DUP 9
A00404:156:HV37TDSXX:3:1273:18638:24001 chr2 57455606 N chr2 57455665 N DUP 6
A00404:155:HV27LDSXX:4:1236:17897:5932 chr2 57455606 N chr2 57455665 N DUP 11
A00404:155:HV27LDSXX:2:1134:6054:13730 chr2 57455632 N chr2 57455723 N DEL 5
A00404:156:HV37TDSXX:4:2542:7301:6402 chr2 57455643 N chr2 57455734 N DEL 4
A00404:155:HV27LDSXX:4:1673:5773:18881 chr5 176837902 N chr5 176837960 N DUP 3
A00404:156:HV37TDSXX:4:2504:3839:9956 chr7 122645382 N chr7 122645585 N DEL 2
A00404:155:HV27LDSXX:3:2368:19515:27085 chr7 122645382 N chr7 122645585 N DEL 7
A00404:155:HV27LDSXX:2:2659:6379:24471 chr7 122645382 N chr7 122645585 N DEL 8
A00297:158:HT275DSXX:2:1118:11406:13949 chr7 122645393 N chr7 122645446 N DEL 13
A00297:158:HT275DSXX:1:1259:5014:35853 chr7 122645393 N chr7 122645446 N DEL 13
A00404:155:HV27LDSXX:3:2548:6370:25582 chr7 122645393 N chr7 122645446 N DEL 13
A00404:155:HV27LDSXX:2:1662:1271:2628 chr7 122645393 N chr7 122645446 N DEL 13
A00404:156:HV37TDSXX:2:1641:13702:24251 chr7 122645469 N chr7 122645548 N DEL 5
A00404:155:HV27LDSXX:1:2370:19551:32628 chr7 122645403 N chr7 122645496 N DUP 5
A00297:158:HT275DSXX:3:2402:5855:9251 chr7 122645406 N chr7 122645461 N DUP 5
A00404:155:HV27LDSXX:2:1623:28980:29168 chr7 122645422 N chr7 122645553 N DUP 3
A00404:155:HV27LDSXX:2:1351:30942:7482 chr1 37896988 N chr1 37897066 N DEL 5
A00297:158:HT275DSXX:1:2302:18141:23171 chr1 37896815 N chr1 37896994 N DUP 5
A00404:155:HV27LDSXX:2:1549:25717:36980 chr1 37896810 N chr1 37896989 N DUP 6
A00297:158:HT275DSXX:1:2459:9471:12320 chr1 37896810 N chr1 37896989 N DUP 10
A00404:155:HV27LDSXX:1:1612:12563:28447 chr1 37896818 N chr1 37896997 N DUP 10
A00404:155:HV27LDSXX:2:1142:20283:34616 chr1 37896859 N chr1 37897040 N DEL 10
A00404:155:HV27LDSXX:4:1436:17607:4210 chr1 37896859 N chr1 37897040 N DEL 5
A00404:156:HV37TDSXX:3:1347:11397:15749 chr16 88015144 N chr16 88015239 N DEL 5
A00404:155:HV27LDSXX:4:1210:27064:15358 chr16 88015144 N chr16 88015239 N DEL 5
A00404:156:HV37TDSXX:2:2629:23014:28604 chr16 88015144 N chr16 88015239 N DEL 5
A00404:156:HV37TDSXX:4:2231:27353:5055 chr16 88015172 N chr16 88015448 N DEL 4
A00404:155:HV27LDSXX:4:1205:32714:4476 chr11 16907376 N chr11 16907553 N DEL 5
A00404:155:HV27LDSXX:2:1632:26467:35587 chr11 16907263 N chr11 16907360 N DUP 15
A00297:158:HT275DSXX:1:2128:30065:35744 chr11 16907261 N chr11 16907407 N DUP 5
A00404:156:HV37TDSXX:3:2653:23014:32800 chr11 16907492 N chr11 16907620 N DEL 2
A00404:155:HV27LDSXX:3:1474:29731:18787 chr11 16907295 N chr11 16907394 N DEL 1
A00297:158:HT275DSXX:2:1406:13069:7717 chr11 16907507 N chr11 16907684 N DEL 5
A00297:158:HT275DSXX:2:1644:13196:16548 chr11 16907521 N chr11 16907647 N DUP 5
A00297:158:HT275DSXX:4:1215:7572:24064 chr11 16907534 N chr11 16907711 N DEL 5
A00404:155:HV27LDSXX:1:1138:23095:1846 chr11 16907358 N chr11 16907711 N DEL 5
A00297:158:HT275DSXX:4:1520:18295:20118 chr11 16907575 N chr11 16907654 N DEL 2
A00404:156:HV37TDSXX:4:2377:26006:33567 chr11 16907286 N chr11 16907688 N DEL 5
A00297:158:HT275DSXX:2:2120:20112:31939 chr11 16907442 N chr11 16907746 N DEL 20
A00404:156:HV37TDSXX:2:1523:23149:20509 chr11 16907489 N chr11 16907871 N DEL 10
A00297:158:HT275DSXX:2:1623:32217:5431 chr11 16907392 N chr11 16907823 N DEL 2
A00404:156:HV37TDSXX:2:1523:23149:20509 chr11 16907489 N chr11 16907871 N DEL 10
A00404:156:HV37TDSXX:4:2103:28194:36793 chr11 16907650 N chr11 16907904 N DEL 27
A00404:155:HV27LDSXX:3:1241:28745:15327 chr11 16907489 N chr11 16907871 N DEL 5
A00404:155:HV27LDSXX:2:2306:6406:23265 chr16 34769747 N chr16 34769913 N DUP 5
A00297:158:HT275DSXX:1:1358:23095:13620 chr10 24767771 N chr10 24767845 N DUP 3
A00404:155:HV27LDSXX:3:1357:27100:19335 chr1 150823850 N chr1 150824143 N DEL 6
A00297:158:HT275DSXX:3:2109:14669:35070 chr1 150823867 N chr1 150824159 N DEL 5
A00404:156:HV37TDSXX:4:2258:26594:19492 chr1 150823885 N chr1 150824177 N DEL 30
A00297:158:HT275DSXX:3:1331:9136:22764 chr1 150823936 N chr1 150824228 N DEL 5
A00404:156:HV37TDSXX:4:2678:6867:15139 chr1 150823838 N chr1 150824129 N DUP 5
A00297:158:HT275DSXX:3:1331:9136:22764 chr1 150823936 N chr1 150824228 N DEL 37
A00297:158:HT275DSXX:3:2109:14073:32471 chr1 150823892 N chr1 150824184 N DEL 5
A00404:155:HV27LDSXX:1:1319:4616:9549 chr1 150823952 N chr1 150824244 N DEL 5
A00404:156:HV37TDSXX:1:2404:28754:2503 chr19 50456207 N chr19 50456468 N DEL 6
A00404:155:HV27LDSXX:4:2641:10276:25332 chr19 50456443 N chr19 50456526 N DUP 2
A00297:158:HT275DSXX:4:2143:22824:8672 chr19 50456443 N chr19 50456526 N DUP 3
A00404:155:HV27LDSXX:2:2610:19208:21825 chr19 50456443 N chr19 50456526 N DUP 4
A00297:158:HT275DSXX:3:1138:30879:9001 chr19 50456233 N chr19 50456538 N DEL 25
A00297:158:HT275DSXX:4:1615:7826:3771 chr19 50456166 N chr19 50456531 N DEL 9
A00297:158:HT275DSXX:1:1434:12057:10128 chr19 50456166 N chr19 50456531 N DEL 9
A00297:158:HT275DSXX:2:2526:21016:16344 chr19 50456341 N chr19 50456553 N DEL 1
A00404:155:HV27LDSXX:3:2376:16984:29528 chr4 8211355 N chr4 8211544 N DUP 5
A00404:156:HV37TDSXX:4:2218:12617:21339 chr4 8211552 N chr4 8211625 N DUP 20
A00404:156:HV37TDSXX:3:2148:15799:21183 chr4 8211395 N chr4 8211553 N DEL 10
A00404:155:HV27LDSXX:3:2656:15646:26209 chr4 8211398 N chr4 8211556 N DEL 10
A00404:156:HV37TDSXX:1:1135:9670:16548 chr8 10852168 N chr8 10852330 N DUP 3
A00404:156:HV37TDSXX:1:2247:1787:33614 chr16 21524909 N chr16 21525146 N DEL 9
A00297:158:HT275DSXX:4:1112:15320:17096 chr16 21524987 N chr16 21525396 N DEL 8
A00404:155:HV27LDSXX:4:1646:12093:7247 chr16 21525010 N chr16 21525268 N DEL 1
A00404:155:HV27LDSXX:2:1249:11876:20556 chr16 21525031 N chr16 21525417 N DUP 3
A00404:155:HV27LDSXX:1:2220:6343:23938 chr16 21524848 N chr16 21525105 N DUP 11
A00404:155:HV27LDSXX:1:2220:6361:23938 chr16 21524848 N chr16 21525105 N DUP 11
A00404:155:HV27LDSXX:3:1324:25961:34397 chr16 21525294 N chr16 21525425 N DEL 16
A00404:155:HV27LDSXX:1:1208:15031:5134 chr16 21525054 N chr16 21525377 N DEL 24
A00404:155:HV27LDSXX:3:1324:25961:34397 chr16 21525294 N chr16 21525425 N DEL 22
A00297:158:HT275DSXX:4:2323:22480:16376 chr21 42140468 N chr21 42140559 N DEL 5
A00297:158:HT275DSXX:1:1654:3170:3223 chr21 42140496 N chr21 42140587 N DEL 1
A00297:158:HT275DSXX:3:1656:5394:18349 chr21 42140451 N chr21 42140586 N DUP 5
A00404:155:HV27LDSXX:1:1652:6578:8500 chr21 42140451 N chr21 42140586 N DUP 5
A00297:158:HT275DSXX:1:1514:20943:2628 chr22 46644367 N chr22 46644476 N DUP 5
A00297:158:HT275DSXX:2:1110:3061:26303 chr22 46644377 N chr22 46644642 N DEL 3
A00404:156:HV37TDSXX:3:2635:17246:18865 chr22 46644386 N chr22 46644717 N DEL 1
A00404:156:HV37TDSXX:2:1478:32389:31782 chr22 46644617 N chr22 46644772 N DEL 10
A00297:158:HT275DSXX:1:1626:20943:30592 chr16 52340348 N chr16 52340429 N DEL 3
A00404:155:HV27LDSXX:3:2533:11767:30201 chr16 52340348 N chr16 52340429 N DEL 5
A00404:156:HV37TDSXX:2:2466:5755:27680 chr16 52340306 N chr16 52340600 N DUP 5
A00404:156:HV37TDSXX:2:1334:13304:13479 chr17 860402 N chr17 860808 N DEL 6
A00404:156:HV37TDSXX:2:2320:23565:15624 chr17 860402 N chr17 860538 N DEL 10
A00404:156:HV37TDSXX:2:2455:17074:28087 chr17 860430 N chr17 860701 N DEL 5
A00404:155:HV27LDSXX:1:2563:24334:1799 chr17 860560 N chr17 860831 N DEL 5
A00404:155:HV27LDSXX:3:2667:7229:20964 chr17 860560 N chr17 860831 N DEL 5
A00404:155:HV27LDSXX:2:2345:4101:36996 chr19 291580 N chr19 291785 N DEL 28
A00404:155:HV27LDSXX:2:2347:17255:10394 chr3 181150146 N chr3 181150310 N DEL 9
A00297:158:HT275DSXX:4:1472:5656:34554 chr3 181150146 N chr3 181150310 N DEL 9
A00404:155:HV27LDSXX:3:1220:11975:30373 chr17 72473680 N chr17 72473747 N DUP 23
A00404:156:HV37TDSXX:4:1564:26060:19664 chr17 72473641 N chr17 72473718 N DEL 16
A00297:158:HT275DSXX:1:1643:18096:5431 chr17 72473641 N chr17 72473718 N DEL 16
A00404:155:HV27LDSXX:3:1610:28167:19617 chr17 72473568 N chr17 72473723 N DEL 7
A00297:158:HT275DSXX:2:2666:26802:4539 chr17 72473574 N chr17 72473729 N DEL 4
A00404:156:HV37TDSXX:2:2266:14751:35524 chr17 72473865 N chr17 72473916 N DUP 19
A00297:158:HT275DSXX:4:1363:19831:14168 chr17 72473865 N chr17 72473916 N DUP 20
A00404:155:HV27LDSXX:3:1524:2257:23469 chr4 32345482 N chr4 32345694 N DEL 6
A00404:156:HV37TDSXX:2:2468:15826:15655 chr2 122452858 N chr2 122452935 N DEL 5
A00404:155:HV27LDSXX:3:2303:2627:31313 chr2 122452858 N chr2 122452935 N DEL 5
A00404:155:HV27LDSXX:3:1110:25409:3286 chr2 122452878 N chr2 122452953 N DUP 5
A00404:156:HV37TDSXX:1:1105:19018:29230 chr2 122452885 N chr2 122452960 N DUP 5
A00404:155:HV27LDSXX:3:1370:3983:16595 chr6 170453167 N chr6 170453303 N DEL 4
A00404:155:HV27LDSXX:4:1675:29803:21699 chr6 170453217 N chr6 170453343 N DUP 5
A00404:155:HV27LDSXX:2:1150:4571:17926 chr16 52618628 N chr16 52618930 N DEL 2
A00297:158:HT275DSXX:4:2606:13910:31876 chr4 162153834 N chr4 162153909 N DEL 27
A00404:155:HV27LDSXX:1:1353:3794:35618 chr4 162153834 N chr4 162153909 N DEL 27
A00404:156:HV37TDSXX:3:2269:3143:2863 chr4 162153792 N chr4 162153871 N DEL 16
A00404:156:HV37TDSXX:4:1224:5936:4852 chr2 35638050 N chr2 35638194 N DEL 5
A00297:158:HT275DSXX:2:2302:14968:10441 chr19 433127 N chr19 433244 N DEL 5
A00404:155:HV27LDSXX:4:1477:9164:18176 chr19 433128 N chr19 433187 N DEL 5
A00297:158:HT275DSXX:1:2147:10429:4930 chr9 2450499 N chr9 2450552 N DEL 18
A00404:156:HV37TDSXX:4:2566:2220:25535 chr9 2450591 N chr9 2450650 N DUP 10
A00297:158:HT275DSXX:2:2303:26413:2613 chr9 2450591 N chr9 2450650 N DUP 8
A00404:156:HV37TDSXX:2:1261:28917:32753 chr22 47814791 N chr22 47814952 N DUP 3
A00404:156:HV37TDSXX:4:1352:31910:12790 chr22 47814787 N chr22 47814964 N DUP 10
A00404:155:HV27LDSXX:3:1361:23918:31078 chr22 47814803 N chr22 47814998 N DUP 4
A00297:158:HT275DSXX:3:1505:3233:3959 chr22 47814808 N chr22 47814967 N DEL 13
A00297:158:HT275DSXX:3:2460:14055:16720 chr19 57990212 N chr19 57990531 N DEL 8
A00404:156:HV37TDSXX:2:2566:22146:28510 chr11 530558 N chr11 530727 N DEL 15
A00297:158:HT275DSXX:4:1632:28022:12508 chr11 530596 N chr11 530653 N DEL 3
A00297:158:HT275DSXX:1:1578:23665:29575 chr11 530596 N chr11 530653 N DEL 5
A00297:158:HT275DSXX:4:1222:19877:35759 chr11 530596 N chr11 530653 N DEL 6
A00297:158:HT275DSXX:2:2602:10203:1814 chr11 530596 N chr11 530653 N DEL 10
A00404:156:HV37TDSXX:4:1420:25889:33176 chr11 530596 N chr11 530653 N DEL 10
A00404:155:HV27LDSXX:4:2178:21269:6699 chr11 530596 N chr11 530653 N DEL 10
A00404:155:HV27LDSXX:1:1502:19036:30326 chr11 530596 N chr11 530653 N DEL 10
A00404:155:HV27LDSXX:1:1502:20645:28855 chr11 530596 N chr11 530653 N DEL 10
A00297:158:HT275DSXX:1:2157:10239:27649 chr11 530596 N chr11 531129 N DEL 10
A00404:155:HV27LDSXX:3:2566:26259:11929 chr11 530596 N chr11 531129 N DEL 10
A00297:158:HT275DSXX:4:1511:16441:4100 chr11 530596 N chr11 531129 N DEL 10
A00297:158:HT275DSXX:4:2122:3143:3114 chr11 530596 N chr11 531129 N DEL 10
A00404:155:HV27LDSXX:1:2574:26259:7012 chr11 530648 N chr11 530761 N DEL 5
A00297:158:HT275DSXX:4:2634:5900:15436 chr11 530648 N chr11 530761 N DEL 5
A00297:158:HT275DSXX:2:1457:8947:18834 chr11 530596 N chr11 530709 N DEL 10
A00297:158:HT275DSXX:1:2207:32687:23156 chr11 530656 N chr11 531217 N DEL 5
A00404:156:HV37TDSXX:1:1251:5837:7968 chr11 530623 N chr11 530736 N DEL 5
A00404:156:HV37TDSXX:4:2224:28348:19742 chr11 530623 N chr11 530736 N DEL 5
A00404:156:HV37TDSXX:4:2224:29640:20008 chr11 530623 N chr11 530736 N DEL 5
A00404:155:HV27LDSXX:3:1231:11849:12900 chr11 530623 N chr11 530736 N DEL 5
A00404:155:HV27LDSXX:3:2409:2573:10269 chr11 530623 N chr11 530736 N DEL 5
A00404:155:HV27LDSXX:4:1450:27868:31031 chr11 530623 N chr11 530736 N DEL 5
A00404:156:HV37TDSXX:4:2461:10565:7670 chr11 530623 N chr11 530736 N DEL 5
A00404:155:HV27LDSXX:1:1613:9661:26772 chr11 530623 N chr11 530876 N DEL 10
A00404:155:HV27LDSXX:3:2525:2293:25191 chr11 530623 N chr11 530736 N DEL 5
A00404:155:HV27LDSXX:1:2254:17671:15875 chr11 530680 N chr11 531267 N DUP 5
A00404:155:HV27LDSXX:4:2267:32217:29669 chr11 530631 N chr11 531022 N DUP 5
A00404:155:HV27LDSXX:4:2267:32217:29669 chr11 530636 N chr11 531027 N DUP 4
A00404:155:HV27LDSXX:4:2658:13829:15421 chr11 530699 N chr11 531064 N DEL 15
A00297:158:HT275DSXX:3:1376:7428:19429 chr11 530606 N chr11 530663 N DEL 5
A00297:158:HT275DSXX:4:2649:10610:7560 chr11 531036 N chr11 531287 N DUP 15
A00404:155:HV27LDSXX:3:2566:26259:11929 chr11 530820 N chr11 531155 N DUP 3
A00297:158:HT275DSXX:2:2510:28230:14058 chr11 530708 N chr11 531129 N DEL 10
A00297:158:HT275DSXX:2:1516:9146:13886 chr11 530708 N chr11 531129 N DEL 10
A00297:158:HT275DSXX:3:2118:9995:21089 chr11 530708 N chr11 531129 N DEL 10
A00404:155:HV27LDSXX:2:1562:18484:3881 chr11 530623 N chr11 530820 N DEL 5
A00404:155:HV27LDSXX:4:2403:1868:12649 chr11 530687 N chr11 530742 N DUP 5
A00297:158:HT275DSXX:1:1378:4616:7357 chr11 530708 N chr11 531129 N DEL 10
A00404:156:HV37TDSXX:4:1417:30499:6245 chr11 530643 N chr11 530700 N DEL 5
A00297:158:HT275DSXX:2:2171:32606:22733 chr11 530681 N chr11 530736 N DUP 5
A00404:155:HV27LDSXX:1:2421:14597:22451 chr11 530740 N chr11 531019 N DUP 10
A00297:158:HT275DSXX:2:1142:26350:20259 chr11 530811 N chr11 531232 N DEL 5
A00404:155:HV27LDSXX:1:1551:30951:30013 chr11 530616 N chr11 530811 N DUP 10
A00404:155:HV27LDSXX:4:1407:9986:23109 chr11 530735 N chr11 530792 N DEL 5
A00404:155:HV27LDSXX:2:2526:26413:35023 chr11 530714 N chr11 530797 N DUP 5
A00404:155:HV27LDSXX:2:1208:23728:27367 chr11 530708 N chr11 531129 N DEL 10
A00404:155:HV27LDSXX:1:1156:16288:9283 chr11 530811 N chr11 531232 N DEL 10
A00404:156:HV37TDSXX:2:2315:15727:15170 chr11 530708 N chr11 531129 N DEL 15
A00297:158:HT275DSXX:3:1431:9923:31735 chr11 530811 N chr11 531232 N DEL 10
A00404:155:HV27LDSXX:2:2467:6479:14497 chr11 530811 N chr11 531204 N DEL 10
A00404:155:HV27LDSXX:3:1655:13557:7999 chr11 530831 N chr11 530988 N DEL 31
A00297:158:HT275DSXX:2:1142:26350:20259 chr11 530708 N chr11 531129 N DEL 15
A00404:155:HV27LDSXX:2:2421:27724:6167 chr11 530831 N chr11 530988 N DEL 31
A00404:156:HV37TDSXX:2:2302:24243:35806 chr11 530737 N chr11 530990 N DEL 5
A00404:155:HV27LDSXX:3:2101:21395:10300 chr11 530811 N chr11 531204 N DEL 15
A00404:156:HV37TDSXX:4:2421:16975:23062 chr11 530623 N chr11 530830 N DUP 20
A00297:158:HT275DSXX:2:2171:32606:22733 chr11 531017 N chr11 531156 N DUP 10
A00404:155:HV27LDSXX:1:1613:9661:26772 chr11 531064 N chr11 531287 N DUP 10
A00297:158:HT275DSXX:2:2622:10059:13557 chr11 530643 N chr11 530812 N DEL 5
A00404:155:HV27LDSXX:4:2159:15600:12947 chr11 530812 N chr11 531035 N DUP 10
A00297:158:HT275DSXX:4:1348:3631:1986 chr11 530735 N chr11 530792 N DEL 5
A00404:155:HV27LDSXX:1:2229:29053:20055 chr11 530812 N chr11 531035 N DUP 10
A00404:155:HV27LDSXX:1:2421:14597:22451 chr11 530708 N chr11 530793 N DEL 10
A00297:158:HT275DSXX:3:1247:23321:13792 chr11 530821 N chr11 531044 N DUP 9
A00297:158:HT275DSXX:3:1676:28863:19319 chr11 530708 N chr11 531129 N DEL 15
A00404:156:HV37TDSXX:1:2119:12780:21120 chr11 530708 N chr11 531129 N DEL 15
A00404:155:HV27LDSXX:2:2455:17336:10473 chr11 530923 N chr11 530980 N DEL 10
A00404:155:HV27LDSXX:4:2368:31774:17315 chr11 530658 N chr11 530855 N DEL 9
A00404:155:HV27LDSXX:2:2455:17336:10473 chr11 531156 N chr11 531295 N DUP 13
A00404:155:HV27LDSXX:1:1502:20645:28855 chr11 530621 N chr11 530706 N DEL 2
A00297:158:HT275DSXX:2:1457:8947:18834 chr11 530700 N chr11 530755 N DUP 5
A00404:155:HV27LDSXX:2:2313:32145:13197 chr11 530644 N chr11 530811 N DUP 10
A00297:158:HT275DSXX:1:1455:12518:30906 chr11 530783 N chr11 531176 N DEL 5
A00297:158:HT275DSXX:2:1150:23493:20008 chr11 530951 N chr11 531288 N DEL 15
A00404:155:HV27LDSXX:3:2622:32136:12430 chr11 530755 N chr11 531176 N DEL 2
A00297:158:HT275DSXX:4:2649:10610:7560 chr11 530932 N chr11 531099 N DUP 10
A00404:156:HV37TDSXX:4:1148:20591:20243 chr11 530775 N chr11 530988 N DEL 26
A00404:155:HV27LDSXX:3:1327:17400:18004 chr11 530945 N chr11 531058 N DEL 1
A00404:155:HV27LDSXX:4:2368:31774:17315 chr11 530597 N chr11 530792 N DUP 10
A00297:158:HT275DSXX:3:1468:10294:34695 chr11 530811 N chr11 531204 N DEL 10
A00404:155:HV27LDSXX:4:1532:2935:12524 chr11 530811 N chr11 531204 N DEL 10
A00297:158:HT275DSXX:4:1511:16441:4100 chr11 530831 N chr11 530988 N DEL 31
A00404:156:HV37TDSXX:2:1173:6325:11631 chr11 530713 N chr11 530966 N DEL 10
A00404:155:HV27LDSXX:3:2622:25391:29904 chr11 530735 N chr11 530960 N DEL 13
A00404:156:HV37TDSXX:1:1567:21395:25300 chr11 530792 N chr11 531017 N DEL 10
A00297:158:HT275DSXX:3:2217:18665:10895 chr11 530980 N chr11 531035 N DUP 10
A00297:158:HT275DSXX:3:1409:31756:16125 chr11 530719 N chr11 530988 N DEL 24
A00404:155:HV27LDSXX:4:2477:22797:7153 chr11 531010 N chr11 531093 N DUP 10
A00297:158:HT275DSXX:3:2549:20980:30373 chr11 531008 N chr11 531091 N DUP 10
A00297:158:HT275DSXX:3:1431:9923:31735 chr11 530811 N chr11 531232 N DEL 9
A00404:155:HV27LDSXX:4:1564:6858:33317 chr11 530988 N chr11 531111 N DUP 29
A00297:158:HT275DSXX:3:1271:20781:20603 chr11 530980 N chr11 531315 N DUP 18
A00404:155:HV27LDSXX:1:2156:17074:22357 chr11 530680 N chr11 531099 N DUP 10
A00404:155:HV27LDSXX:3:2622:26142:29042 chr11 530711 N chr11 531048 N DEL 3
A00404:155:HV27LDSXX:2:2103:24876:31266 chr11 530742 N chr11 531105 N DUP 10
A00404:156:HV37TDSXX:1:2349:19343:35305 chr11 531129 N chr11 531212 N DUP 5
A00404:155:HV27LDSXX:2:2273:4517:33520 chr11 530760 N chr11 530983 N DUP 3
A00404:155:HV27LDSXX:2:1433:14931:22592 chr11 530616 N chr11 530811 N DUP 10
A00404:155:HV27LDSXX:1:1218:25635:23844 chr11 530792 N chr11 531129 N DEL 5
A00404:156:HV37TDSXX:4:2678:29903:35869 chr11 531156 N chr11 531267 N DUP 10
A00404:156:HV37TDSXX:2:1665:15320:26240 chr11 530682 N chr11 531017 N DUP 5
A00297:158:HT275DSXX:3:2413:10637:36824 chr11 530848 N chr11 531155 N DUP 10
A00404:155:HV27LDSXX:1:1566:26286:25034 chr11 530651 N chr11 530820 N DEL 5
A00404:155:HV27LDSXX:4:2365:18295:31140 chr11 531156 N chr11 531267 N DUP 10
A00404:155:HV27LDSXX:1:1535:16315:11553 chr11 531212 N chr11 531267 N DUP 10
A00404:155:HV27LDSXX:4:1309:22950:11428 chr11 530811 N chr11 531204 N DEL 14
A00297:158:HT275DSXX:4:2133:29649:18333 chr11 530811 N chr11 531204 N DEL 15
A00297:158:HT275DSXX:3:2168:27109:2722 chr11 530811 N chr11 531204 N DEL 15
A00297:158:HT275DSXX:3:2168:28293:2769 chr11 530811 N chr11 531204 N DEL 15
A00404:155:HV27LDSXX:2:2273:4517:33520 chr11 530708 N chr11 531239 N DUP 5
A00297:158:HT275DSXX:2:2402:11324:3756 chr11 530699 N chr11 531204 N DEL 15
A00297:158:HT275DSXX:3:2217:18665:10895 chr11 530615 N chr11 530980 N DEL 10
A00404:155:HV27LDSXX:1:1509:18801:15859 chr11 530817 N chr11 531238 N DEL 6
A00404:155:HV27LDSXX:3:2622:32136:12430 chr11 531017 N chr11 531186 N DEL 14
A00404:155:HV27LDSXX:3:2543:8368:33238 chr11 530625 N chr11 531016 N DUP 5
A00404:155:HV27LDSXX:4:1625:4110:8923 chr11 530699 N chr11 531204 N DEL 6
A00297:158:HT275DSXX:3:1413:12924:30420 chr11 531021 N chr11 531190 N DEL 10
A00404:155:HV27LDSXX:1:2359:14986:9408 chr11 530699 N chr11 531204 N DEL 5
A00297:158:HT275DSXX:4:2256:18005:11256 chr11 530951 N chr11 531288 N DEL 10
A00404:156:HV37TDSXX:2:1154:7202:6042 chr11 531155 N chr11 531268 N DEL 11
A00404:156:HV37TDSXX:1:2126:4318:35336 chr11 530690 N chr11 531361 N DUP 9
A00404:156:HV37TDSXX:1:2126:4327:35196 chr11 530690 N chr11 531361 N DUP 9
A00404:156:HV37TDSXX:3:2573:30020:14559 chr11 530690 N chr11 531361 N DUP 10
A00404:156:HV37TDSXX:1:2335:21730:25880 chr11 530755 N chr11 531288 N DEL 12
A00404:156:HV37TDSXX:1:1403:28411:7357 chr11 530690 N chr11 531361 N DUP 10
A00404:155:HV27LDSXX:2:2222:15944:7905 chr11 530690 N chr11 531361 N DUP 10
A00404:156:HV37TDSXX:4:2163:31955:29872 chr11 530755 N chr11 531288 N DEL 5
A00404:155:HV27LDSXX:4:1478:18322:32283 chr11 530643 N chr11 531288 N DEL 10
A00404:155:HV27LDSXX:2:2402:19271:26443 chr11 530643 N chr11 531288 N DEL 10
A00404:155:HV27LDSXX:2:2313:32533:13526 chr11 530643 N chr11 531288 N DEL 10
A00404:155:HV27LDSXX:3:1103:28565:15483 chr11 530643 N chr11 531288 N DEL 10
A00404:155:HV27LDSXX:3:1467:28004:15922 chr11 530643 N chr11 531288 N DEL 10
A00404:156:HV37TDSXX:4:2269:22779:3364 chr11 530727 N chr11 531288 N DEL 5
A00404:156:HV37TDSXX:4:1560:21730:12164 chr11 530791 N chr11 531352 N DEL 15
A00404:156:HV37TDSXX:4:2617:25156:32221 chr11 530643 N chr11 531288 N DEL 5
A00404:156:HV37TDSXX:2:2227:30337:3646 chr11 530615 N chr11 531288 N DEL 5
A00404:156:HV37TDSXX:3:2666:9263:6856 chr11 530619 N chr11 531292 N DEL 5
A00404:155:HV27LDSXX:4:1526:25789:18505 chr11 531261 N chr11 531374 N DEL 40
A00404:155:HV27LDSXX:4:2227:20184:35634 chr11 530791 N chr11 531380 N DEL 55
A00404:156:HV37TDSXX:3:1354:4788:19366 chr11 531093 N chr11 531374 N DEL 23
A00404:155:HV27LDSXX:4:2227:20184:35634 chr11 530623 N chr11 531380 N DEL 15
A00404:155:HV27LDSXX:1:1178:26060:26490 chr5 165345537 N chr5 165345626 N DUP 7
A00404:155:HV27LDSXX:4:1450:14859:20682 chr5 165345541 N chr5 165345656 N DUP 8
A00404:155:HV27LDSXX:4:1450:15736:19820 chr5 165345541 N chr5 165345656 N DUP 8
A00297:158:HT275DSXX:3:2665:30246:26349 chr14 103616107 N chr14 103616586 N DEL 8
A00297:158:HT275DSXX:2:1622:29279:36354 chr14 103616107 N chr14 103616586 N DEL 10
A00404:155:HV27LDSXX:3:1664:31159:13651 chr14 103616155 N chr14 103616310 N DEL 5
A00404:156:HV37TDSXX:2:2556:22290:2988 chr14 103616155 N chr14 103616310 N DEL 5
A00404:155:HV27LDSXX:3:1163:30689:32315 chr14 103616134 N chr14 103616611 N DUP 6
A00404:156:HV37TDSXX:4:1246:13612:19366 chr14 103616175 N chr14 103616328 N DUP 5
A00404:156:HV37TDSXX:4:1246:13666:19617 chr14 103616175 N chr14 103616328 N DUP 5
A00404:156:HV37TDSXX:3:2365:8458:11506 chr14 103616176 N chr14 103616329 N DUP 4
A00404:156:HV37TDSXX:3:1334:27905:3818 chr11 2472196 N chr11 2472342 N DUP 2
A00404:156:HV37TDSXX:3:1477:8359:12336 chr11 2472196 N chr11 2472342 N DUP 5
A00404:156:HV37TDSXX:3:1477:8531:12696 chr11 2472196 N chr11 2472342 N DUP 5
A00297:158:HT275DSXX:2:1518:24478:17769 chr11 2472196 N chr11 2472342 N DUP 5
A00404:155:HV27LDSXX:4:2553:15971:2722 chr11 2472196 N chr11 2472342 N DUP 5
A00404:155:HV27LDSXX:1:2448:23583:15029 chr11 2472254 N chr11 2472402 N DEL 5
A00404:155:HV27LDSXX:4:2307:9733:19695 chr11 2472132 N chr11 2472402 N DEL 5
A00297:158:HT275DSXX:2:2651:26883:36025 chr11 2472132 N chr11 2472402 N DEL 5
A00297:158:HT275DSXX:3:1302:20021:13338 chr11 2472144 N chr11 2472414 N DEL 3
A00404:156:HV37TDSXX:4:1650:18710:6652 chr11 2472145 N chr11 2472415 N DEL 2
A00297:158:HT275DSXX:3:2227:32515:20635 chr2 236594072 N chr2 236594374 N DEL 5
A00297:158:HT275DSXX:3:2227:32515:20635 chr2 236594072 N chr2 236594374 N DEL 7
A00404:156:HV37TDSXX:1:1169:31964:13823 chr2 236594114 N chr2 236594220 N DEL 36
A00404:155:HV27LDSXX:1:2269:23701:27132 chr3 40212259 N chr3 40212338 N DEL 4
A00404:155:HV27LDSXX:1:1412:17472:11146 chr3 40212267 N chr3 40212346 N DEL 9
A00404:155:HV27LDSXX:4:1535:22562:14700 chr3 40212250 N chr3 40212303 N DEL 5
A00297:158:HT275DSXX:3:1371:5927:33739 chr3 40212279 N chr3 40212334 N DEL 15
A00404:156:HV37TDSXX:1:2651:22589:17159 chr3 40212279 N chr3 40212334 N DEL 17
A00404:155:HV27LDSXX:4:2553:22390:33191 chr3 40212279 N chr3 40212334 N DEL 17
A00297:158:HT275DSXX:4:2552:5141:21981 chr3 40212279 N chr3 40212334 N DEL 17
A00404:155:HV27LDSXX:2:1233:26648:23750 chr3 40212279 N chr3 40212334 N DEL 17
A00404:155:HV27LDSXX:2:1233:27064:23218 chr3 40212279 N chr3 40212334 N DEL 17
A00404:155:HV27LDSXX:2:1233:27633:23516 chr3 40212279 N chr3 40212334 N DEL 17
A00404:155:HV27LDSXX:4:1120:14868:36793 chr3 40212279 N chr3 40212334 N DEL 26
A00404:155:HV27LDSXX:4:1120:15474:36151 chr3 40212279 N chr3 40212334 N DEL 26
A00404:156:HV37TDSXX:4:1410:13449:32142 chr3 40212279 N chr3 40212334 N DEL 31
A00297:158:HT275DSXX:2:1424:25192:7232 chr3 40212279 N chr3 40212334 N DEL 34
A00404:156:HV37TDSXX:2:1658:32063:20384 chr3 40212279 N chr3 40212334 N DEL 40
A00297:158:HT275DSXX:3:2253:27245:15577 chr3 40212279 N chr3 40212334 N DEL 21
A00404:155:HV27LDSXX:4:2213:32090:12414 chr3 40212279 N chr3 40212334 N DEL 15
A00404:156:HV37TDSXX:4:2255:10755:25222 chr1 161243725 N chr1 161244009 N DUP 5
A00297:158:HT275DSXX:2:2311:28754:17660 chr1 161243725 N chr1 161244009 N DUP 5
A00404:156:HV37TDSXX:1:2646:14751:36182 chr1 161243725 N chr1 161244009 N DUP 5
A00404:155:HV27LDSXX:1:1323:10357:36871 chr1 161243725 N chr1 161244009 N DUP 5
A00404:155:HV27LDSXX:2:1139:19714:3192 chr1 161243725 N chr1 161244009 N DUP 5
A00404:155:HV27LDSXX:4:1647:26196:16986 chr1 161243725 N chr1 161244009 N DUP 5
A00297:158:HT275DSXX:3:1547:5177:26584 chr1 161243725 N chr1 161244009 N DUP 5
A00404:156:HV37TDSXX:2:2360:1895:9846 chr1 161243725 N chr1 161244009 N DUP 5
A00297:158:HT275DSXX:1:2626:13548:10676 chr1 161243742 N chr1 161244028 N DEL 5
A00404:156:HV37TDSXX:3:1616:25654:3521 chrX 153891705 N chrX 153892000 N DEL 5
A00404:155:HV27LDSXX:2:1343:24614:4507 chrX 153891685 N chrX 153891978 N DUP 5
A00404:156:HV37TDSXX:3:1322:3287:22654 chrX 153891582 N chrX 153891877 N DEL 4
A00297:158:HT275DSXX:4:2520:20889:26584 chr12 93226062 N chr12 93226112 N DUP 8
A00404:156:HV37TDSXX:1:2128:23836:32878 chr12 93226062 N chr12 93226112 N DUP 8
A00404:156:HV37TDSXX:4:2332:8721:19100 chr12 93226062 N chr12 93226112 N DUP 8
A00297:158:HT275DSXX:4:2506:22797:14575 chr12 93226062 N chr12 93226112 N DUP 8
A00404:156:HV37TDSXX:3:1529:8250:5541 chr12 93226113 N chr12 93226171 N DEL 10
A00404:155:HV27LDSXX:3:1457:32678:27211 chr12 93226113 N chr12 93226171 N DEL 26
A00404:156:HV37TDSXX:3:1107:5113:15984 chr12 93226113 N chr12 93226171 N DEL 26
A00404:155:HV27LDSXX:3:2512:30427:7748 chr12 93226113 N chr12 93226171 N DEL 26
A00404:156:HV37TDSXX:3:2309:19461:30812 chr12 93226113 N chr12 93226171 N DEL 26
A00297:158:HT275DSXX:1:2178:19452:16297 chr12 93226113 N chr12 93226171 N DEL 20
A00297:158:HT275DSXX:2:2111:2013:30342 chr12 93226113 N chr12 93226171 N DEL 12
A00297:158:HT275DSXX:1:2675:8594:33129 chr12 93226113 N chr12 93226171 N DEL 17
A00404:155:HV27LDSXX:4:1142:31087:28056 chr12 93226113 N chr12 93226171 N DEL 8
A00404:155:HV27LDSXX:4:2119:8666:21825 chr12 93226045 N chr12 93226171 N DEL 8
A00297:158:HT275DSXX:4:1153:27010:17300 chr10 739761 N chr10 739888 N DUP 4
A00297:158:HT275DSXX:1:1237:4390:7185 chr10 739739 N chr10 739894 N DUP 11
A00297:158:HT275DSXX:2:2124:11324:6887 chr10 739746 N chr10 739901 N DEL 11
A00404:156:HV37TDSXX:4:1303:26377:5525 chr10 739746 N chr10 739901 N DEL 11
A00297:158:HT275DSXX:3:1172:2211:1971 chr10 739778 N chr10 739913 N DEL 3
A00404:155:HV27LDSXX:2:1222:29405:17534 chr8 26929328 N chr8 26929387 N DEL 6
A00404:156:HV37TDSXX:1:1363:18936:26960 chr12 52935547 N chr12 52935692 N DUP 1
A00404:156:HV37TDSXX:2:1571:8992:11240 chr12 52935544 N chr12 52935678 N DUP 2
A00404:156:HV37TDSXX:1:2239:28266:16814 chr2 201260035 N chr2 201260114 N DUP 1
A00297:158:HT275DSXX:2:2522:8829:32471 chr17 82579585 N chr17 82580145 N DEL 5
A00404:156:HV37TDSXX:3:1277:5475:29951 chr17 82579689 N chr17 82580739 N DEL 4
A00297:158:HT275DSXX:3:1340:12888:14857 chr17 82579784 N chr17 82579992 N DUP 5
A00404:156:HV37TDSXX:1:1138:15600:9314 chr17 82579994 N chr17 82580135 N DEL 5
A00297:158:HT275DSXX:4:2626:19090:35963 chr17 82580106 N chr17 82580247 N DEL 5
A00404:156:HV37TDSXX:3:1508:12400:34835 chr17 82580016 N chr17 82580085 N DUP 5
A00297:158:HT275DSXX:2:2140:20943:27837 chr17 82580104 N chr17 82580245 N DEL 5
A00404:156:HV37TDSXX:1:2224:2474:35556 chr17 82580174 N chr17 82580245 N DEL 5
A00404:156:HV37TDSXX:1:2503:17047:29230 chr17 82579856 N chr17 82580067 N DEL 6
A00404:156:HV37TDSXX:1:1323:27091:23140 chr17 82580177 N chr17 82580248 N DEL 5
A00404:156:HV37TDSXX:2:2502:21305:16344 chr17 82579670 N chr17 82580158 N DUP 4
A00404:156:HV37TDSXX:1:1430:26368:28651 chr17 82579672 N chr17 82580162 N DEL 5
A00297:158:HT275DSXX:4:2626:19090:35963 chr17 82579666 N chr17 82580576 N DEL 5
A00297:158:HT275DSXX:3:2347:31575:17879 chr17 82579990 N chr17 82580271 N DEL 5
A00297:158:HT275DSXX:1:2232:17074:3630 chr17 82580179 N chr17 82580248 N DUP 5
A00404:156:HV37TDSXX:1:2224:2474:35556 chr17 82579727 N chr17 82580427 N DEL 5
A00404:156:HV37TDSXX:2:2332:24523:29841 chr17 82579672 N chr17 82580372 N DEL 10
A00297:158:HT275DSXX:3:2239:17381:18537 chr17 82579695 N chr17 82580535 N DEL 5
A00404:156:HV37TDSXX:3:1274:20518:30201 chr17 82580400 N chr17 82580472 N DEL 5
A00404:156:HV37TDSXX:4:2550:17815:30436 chr17 82580034 N chr17 82580455 N DEL 10
A00404:156:HV37TDSXX:3:1508:12400:34835 chr17 82579596 N chr17 82580506 N DEL 5
A00404:155:HV27LDSXX:4:2155:10176:9815 chr17 82580575 N chr17 82580786 N DEL 5
A00404:155:HV27LDSXX:4:1360:23719:10942 chr17 82580226 N chr17 82580575 N DUP 3
A00297:158:HT275DSXX:4:2114:30635:17002 chr17 82580227 N chr17 82580716 N DUP 5
A00297:158:HT275DSXX:4:2443:20681:18552 chr17 82580506 N chr17 82580785 N DUP 5
A00404:155:HV27LDSXX:2:2403:24162:2628 chr17 82579899 N chr17 82580738 N DUP 5
A00404:156:HV37TDSXX:2:1458:19027:33786 chr17 82579667 N chr17 82580085 N DUP 5
A00404:155:HV27LDSXX:3:1275:7392:18803 chr17 82580506 N chr17 82580785 N DUP 5
A00404:155:HV27LDSXX:3:1612:28031:11741 chr17 82580088 N chr17 82580789 N DEL 5
A00404:156:HV37TDSXX:2:2310:3007:6073 chr17 82580642 N chr17 82580711 N DUP 5
A00404:156:HV37TDSXX:2:1474:12943:1986 chr17 82580477 N chr17 82580756 N DUP 5
A00404:155:HV27LDSXX:3:2656:8757:8891 chr17 82580506 N chr17 82580785 N DUP 5
A00404:155:HV27LDSXX:3:1417:19081:29496 chr17 82580109 N chr17 82580738 N DUP 5
A00404:155:HV27LDSXX:4:1360:23719:10942 chr17 82579684 N chr17 82580032 N DUP 4
A00297:158:HT275DSXX:1:1636:23728:26960 chr17 82580253 N chr17 82581024 N DEL 5
A00404:156:HV37TDSXX:2:1655:21513:21809 chr17 82580087 N chr17 82581068 N DEL 5
A00404:156:HV37TDSXX:2:1655:21513:21809 chr17 82580087 N chr17 82581068 N DEL 5
A00404:155:HV27LDSXX:3:1117:13268:31735 chr17 82580088 N chr17 82581069 N DEL 5
A00297:158:HT275DSXX:1:1174:13801:4163 chr22 48956663 N chr22 48957028 N DEL 7
A00404:155:HV27LDSXX:4:2511:20790:24815 chr22 48956601 N chr22 48957034 N DEL 2
A00404:156:HV37TDSXX:1:2242:11559:33661 chr22 48956510 N chr22 48957092 N DEL 1
A00404:156:HV37TDSXX:1:2406:30011:3615 chr22 48956510 N chr22 48957092 N DEL 1
A00297:158:HT275DSXX:1:1432:2474:28228 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:1:1633:12680:11522 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:1:2364:30273:21699 chr6 154481281 N chr6 154481553 N DUP 7
A00404:155:HV27LDSXX:3:2609:31177:13933 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:2:1449:4083:18521 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:4:2329:11767:10473 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:3:2260:31250:18192 chr6 154481281 N chr6 154481553 N DUP 7
A00404:156:HV37TDSXX:3:2264:32009:16720 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:2:1429:31340:17628 chr6 154481281 N chr6 154481553 N DUP 7
A00404:155:HV27LDSXX:3:1133:26096:15217 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:4:1360:20193:1360 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:4:1618:5104:17848 chr6 154481281 N chr6 154481553 N DUP 7
A00297:158:HT275DSXX:1:1321:14606:19304 chr6 154481281 N chr6 154481553 N DEL 7
A00404:156:HV37TDSXX:3:1435:26196:6527 chr6 154481281 N chr6 154481553 N DEL 7
A00404:155:HV27LDSXX:3:2163:11686:5635 chr2 141324073 N chr2 141324146 N DEL 11
A00404:156:HV37TDSXX:3:1305:27190:24095 chr2 141324072 N chr2 141324145 N DEL 10
A00404:155:HV27LDSXX:1:2647:2013:13777 chr2 141324039 N chr2 141324180 N DEL 7
A00404:155:HV27LDSXX:2:1626:4417:20635 chr2 141324040 N chr2 141324181 N DEL 7
A00297:158:HT275DSXX:3:1259:18945:26130 chr2 141324181 N chr2 141324330 N DUP 8
A00297:158:HT275DSXX:2:1123:1362:36730 chr2 141324043 N chr2 141324184 N DEL 7
A00297:158:HT275DSXX:2:1123:1515:36902 chr2 141324043 N chr2 141324184 N DEL 7
A00404:155:HV27LDSXX:3:2612:27163:16783 chr2 141324044 N chr2 141324187 N DEL 9
A00404:155:HV27LDSXX:4:2662:16893:35133 chr2 141324052 N chr2 141324193 N DEL 2
A00404:156:HV37TDSXX:1:1309:19985:18161 chr8 23040423 N chr8 23040476 N DEL 5
A00297:158:HT275DSXX:3:2502:19343:13166 chr8 23040423 N chr8 23040476 N DEL 5
A00404:156:HV37TDSXX:3:1306:4010:22404 chr8 23040423 N chr8 23040558 N DEL 8
A00404:155:HV27LDSXX:1:2430:1163:3630 chr8 23040423 N chr8 23040558 N DEL 16
A00404:156:HV37TDSXX:4:1629:2718:17754 chr8 23040423 N chr8 23040558 N DEL 20
A00404:156:HV37TDSXX:3:2263:30535:28980 chr8 23040423 N chr8 23040558 N DEL 22
A00404:156:HV37TDSXX:3:2227:19253:21527 chr8 23040443 N chr8 23040520 N DEL 28
A00404:155:HV27LDSXX:1:2628:18466:1219 chr8 23040443 N chr8 23040520 N DEL 28
A00404:155:HV27LDSXX:3:2354:27489:2910 chr8 23040443 N chr8 23040520 N DEL 28
A00404:156:HV37TDSXX:2:1477:13829:14700 chr8 23040443 N chr8 23040520 N DEL 28
A00404:155:HV27LDSXX:4:2562:1461:7529 chr8 23040443 N chr8 23040520 N DEL 14
A00404:156:HV37TDSXX:3:1651:30599:31469 chr8 23040548 N chr8 23040603 N DUP 21
A00404:156:HV37TDSXX:3:2140:19759:6151 chr8 23040548 N chr8 23040603 N DUP 21
A00297:158:HT275DSXX:2:2327:15393:12618 chr8 23040548 N chr8 23040603 N DUP 20
A00404:156:HV37TDSXX:2:1162:17146:29559 chr8 23040548 N chr8 23040603 N DUP 19
A00404:155:HV27LDSXX:3:2318:29188:34381 chr8 23040548 N chr8 23040603 N DUP 13
A00404:155:HV27LDSXX:3:2319:32063:1344 chr8 23040548 N chr8 23040603 N DUP 13
A00404:156:HV37TDSXX:2:2578:5909:30295 chr8 23040514 N chr8 23040574 N DEL 10
A00404:155:HV27LDSXX:4:2450:19678:5509 chr8 23040514 N chr8 23040574 N DEL 10
A00404:155:HV27LDSXX:2:2472:23357:5024 chr8 23040514 N chr8 23040574 N DEL 10
A00404:156:HV37TDSXX:2:1318:1606:5588 chr8 23040514 N chr8 23040574 N DEL 10
A00297:158:HT275DSXX:2:2160:29857:23390 chr8 23040514 N chr8 23040574 N DEL 10
A00404:156:HV37TDSXX:4:2115:3622:4038 chr8 23040488 N chr8 23040574 N DEL 8
A00404:155:HV27LDSXX:1:1638:18991:9737 chr8 23040516 N chr8 23040576 N DEL 6
A00404:155:HV27LDSXX:1:2253:10212:28635 chr8 23040423 N chr8 23040616 N DEL 7
A00297:158:HT275DSXX:4:2252:23565:16250 chr8 23040424 N chr8 23040617 N DEL 7
A00297:158:HT275DSXX:4:2252:23701:19617 chr8 23040424 N chr8 23040617 N DEL 7
A00404:156:HV37TDSXX:3:1306:4010:22404 chr8 23040477 N chr8 23040620 N DEL 7
A00297:158:HT275DSXX:1:2371:19045:23484 chr8 23040478 N chr8 23040621 N DEL 7
A00404:156:HV37TDSXX:1:1509:28194:33411 chr13 76480616 N chr13 76480665 N DUP 10
A00404:155:HV27LDSXX:1:1512:9064:9236 chr10 80357054 N chr10 80357130 N DEL 14
A00404:155:HV27LDSXX:2:2545:2121:27492 chr6 47418043 N chr6 47418120 N DUP 6
A00404:156:HV37TDSXX:4:2629:2492:35399 chr14 84099656 N chr14 84099749 N DEL 5
A00404:156:HV37TDSXX:2:2477:9598:21746 chr14 84099656 N chr14 84099749 N DEL 5
A00404:155:HV27LDSXX:4:1133:9173:23140 chr14 84099907 N chr14 84100140 N DEL 5
A00297:158:HT275DSXX:3:1348:2257:22529 chr14 84099853 N chr14 84099934 N DEL 21
A00297:158:HT275DSXX:3:1348:2257:22529 chr14 84099934 N chr14 84100162 N DUP 13
A00404:156:HV37TDSXX:2:1359:21043:21120 chr1 4964478 N chr1 4964538 N DUP 5
A00297:158:HT275DSXX:1:1318:21974:34068 chr17 77809939 N chr17 77810190 N DEL 1
A00404:155:HV27LDSXX:2:2110:30418:28275 chr17 77809976 N chr17 77810239 N DEL 5
A00404:156:HV37TDSXX:3:1644:7184:25551 chr17 77810018 N chr17 77810254 N DEL 5
A00404:155:HV27LDSXX:3:1564:24804:36746 chr17 77810044 N chr17 77810258 N DEL 1
A00404:155:HV27LDSXX:2:2514:2193:19914 chr11 1429384 N chr11 1429480 N DEL 7
A00297:158:HT275DSXX:2:1429:15374:6793 chr11 1429384 N chr11 1429480 N DEL 9
A00297:158:HT275DSXX:3:1265:6533:15154 chr11 1429384 N chr11 1429480 N DEL 19
A00297:158:HT275DSXX:4:1259:13955:11036 chr11 1429305 N chr11 1429556 N DUP 4
A00404:155:HV27LDSXX:2:2368:15845:10488 chr11 1429392 N chr11 1429488 N DEL 7
A00404:156:HV37TDSXX:1:2134:25229:4726 chr11 1429392 N chr11 1429488 N DEL 7
A00404:155:HV27LDSXX:4:1335:21124:34882 chr11 1429395 N chr11 1429491 N DEL 4
A00404:155:HV27LDSXX:4:1335:22236:29293 chr11 1429395 N chr11 1429491 N DEL 4
A00404:156:HV37TDSXX:4:1572:32750:9236 chr11 1429394 N chr11 1429490 N DEL 5
A00404:155:HV27LDSXX:1:2235:2727:31673 chr5 157849014 N chr5 157849151 N DEL 31
A00297:158:HT275DSXX:4:1501:19940:6621 chr5 157895076 N chr5 157895260 N DEL 6
A00404:156:HV37TDSXX:1:1144:31684:19633 chr5 157895150 N chr5 157895334 N DEL 14
A00297:158:HT275DSXX:1:2160:2862:10300 chr5 157895060 N chr5 157895244 N DEL 7
A00404:156:HV37TDSXX:1:1144:31684:19633 chr5 157895150 N chr5 157895334 N DEL 28
A00404:156:HV37TDSXX:3:1659:11586:1705 chr11 3217035 N chr11 3217105 N DUP 6
A00404:156:HV37TDSXX:4:2307:1597:25958 chr8 100723910 N chr8 100724042 N DUP 4
A00297:158:HT275DSXX:3:2315:23023:16595 chr8 100723851 N chr8 100723987 N DEL 16
A00297:158:HT275DSXX:1:2449:3613:35305 chrX 3434773 N chrX 3435141 N DEL 14
A00404:156:HV37TDSXX:1:1114:1199:9111 chr13 60601172 N chr13 60601227 N DEL 34
A00404:155:HV27LDSXX:2:2404:27163:31657 chr7 57444620 N chr7 57444922 N DUP 1
A00404:155:HV27LDSXX:4:1604:2148:13416 chr7 57444929 N chr7 57445069 N DEL 10
A00404:155:HV27LDSXX:1:2607:4146:29496 chr7 57444535 N chr7 57444965 N DUP 2
A00404:156:HV37TDSXX:1:2376:4218:8516 chr7 57444669 N chr7 57444965 N DUP 6
A00404:155:HV27LDSXX:2:1161:20030:12320 chr7 57444869 N chr7 57444971 N DUP 4
A00297:158:HT275DSXX:3:1443:13648:22122 chr7 57444691 N chr7 57444909 N DEL 7
A00404:155:HV27LDSXX:3:2345:18756:34601 chr7 57444946 N chr7 57445084 N DUP 7
A00297:158:HT275DSXX:3:2238:14904:22388 chr7 57444646 N chr7 57444952 N DEL 4
A00404:156:HV37TDSXX:4:1374:23041:25864 chr10 128129464 N chr10 128129519 N DEL 12
A00404:155:HV27LDSXX:2:1675:16016:13792 chr10 128129464 N chr10 128129519 N DEL 14
A00404:155:HV27LDSXX:1:1451:21612:25739 chr10 128129464 N chr10 128129519 N DEL 15
A00404:156:HV37TDSXX:3:2326:29839:14434 chr10 128129464 N chr10 128129519 N DEL 26
A00404:155:HV27LDSXX:2:1205:17137:33739 chr10 128129464 N chr10 128129519 N DEL 26
A00404:156:HV37TDSXX:2:2227:25247:27618 chr10 128129464 N chr10 128129519 N DEL 26
A00404:156:HV37TDSXX:1:2351:32768:2033 chr10 128129489 N chr10 128129542 N DUP 5
A00404:156:HV37TDSXX:2:2411:3558:9220 chr10 128129464 N chr10 128129519 N DEL 19
A00404:155:HV27LDSXX:4:1102:10773:9095 chr10 128129471 N chr10 128129526 N DEL 4
A00297:158:HT275DSXX:4:1223:4571:23093 chr7 73648713 N chr7 73649085 N DEL 6
A00297:158:HT275DSXX:4:1269:28284:30655 chr7 73648790 N chr7 73649156 N DUP 4
A00404:155:HV27LDSXX:1:2237:16830:23657 chr7 73648934 N chr7 73649099 N DEL 8
A00297:158:HT275DSXX:3:2356:19099:30686 chr7 73648616 N chr7 73649331 N DUP 5
A00404:156:HV37TDSXX:1:1424:19199:30107 chr1 194028671 N chr1 194028745 N DUP 15
A00297:158:HT275DSXX:3:1414:13856:20415 chr1 194028622 N chr1 194028684 N DEL 2
A00404:156:HV37TDSXX:3:1304:14814:17566 chr1 194028691 N chr1 194028765 N DUP 4
A00404:156:HV37TDSXX:3:1304:15013:18317 chr1 194028682 N chr1 194028756 N DUP 4
A00297:158:HT275DSXX:2:1613:32597:28917 chr1 194028632 N chr1 194028824 N DUP 4
A00404:155:HV27LDSXX:3:1138:4752:6151 chr1 194028626 N chr1 194028757 N DEL 6
A00404:155:HV27LDSXX:3:1138:5755:6950 chr1 194028626 N chr1 194028757 N DEL 6
A00297:158:HT275DSXX:2:1565:10013:12352 chr1 194028706 N chr1 194028850 N DEL 12
A00404:155:HV27LDSXX:4:1514:12427:18474 chr1 194028709 N chr1 194028853 N DEL 12
A00297:158:HT275DSXX:2:2545:32000:21402 chr1 194028713 N chr1 194028857 N DEL 8
A00297:158:HT275DSXX:2:2545:32344:21308 chr1 194028713 N chr1 194028857 N DEL 8
A00297:158:HT275DSXX:2:2643:7030:33739 chr1 194028713 N chr1 194028857 N DEL 8
A00297:158:HT275DSXX:2:1253:32452:21402 chr15 80400864 N chr15 80401193 N DEL 17
A00404:155:HV27LDSXX:2:1339:29387:13714 chr12 129538960 N chr12 129539081 N DEL 5
A00297:158:HT275DSXX:3:2463:5077:34804 chr12 129538960 N chr12 129539081 N DEL 5
A00404:155:HV27LDSXX:2:2678:21929:32925 chr12 129538960 N chr12 129539081 N DEL 5
A00404:156:HV37TDSXX:1:2233:32768:18443 chr12 129538960 N chr12 129539081 N DEL 5
A00404:156:HV37TDSXX:3:1664:24469:9204 chr12 129538960 N chr12 129539081 N DEL 5
A00404:155:HV27LDSXX:2:1333:26521:29199 chr12 129538960 N chr12 129539081 N DEL 5
A00404:156:HV37TDSXX:2:2273:19759:18239 chr12 129538960 N chr12 129539081 N DEL 5
A00404:155:HV27LDSXX:1:1127:7591:23469 chr12 129538960 N chr12 129539081 N DEL 5
A00404:156:HV37TDSXX:1:1355:3766:30185 chr12 129538960 N chr12 129539081 N DEL 5
A00404:156:HV37TDSXX:2:2139:20961:29309 chr12 129538969 N chr12 129539050 N DEL 5
A00404:155:HV27LDSXX:3:1464:30065:14105 chr12 129538961 N chr12 129539080 N DUP 2
A00404:155:HV27LDSXX:1:1541:2483:12649 chr12 129538961 N chr12 129539080 N DUP 5
A00297:158:HT275DSXX:2:1309:5990:3161 chr12 129538961 N chr12 129539080 N DUP 5
A00297:158:HT275DSXX:2:1309:7274:28964 chr12 129538961 N chr12 129539080 N DUP 5
A00297:158:HT275DSXX:2:1309:7283:28948 chr12 129538961 N chr12 129539080 N DUP 5
A00297:158:HT275DSXX:1:1527:14425:13260 chr12 129539024 N chr12 129539144 N DUP 16
A00297:158:HT275DSXX:3:1365:7726:32597 chr12 129539036 N chr12 129539115 N DUP 18
A00297:158:HT275DSXX:3:2563:8739:31908 chr12 129539036 N chr12 129539155 N DUP 14
A00404:156:HV37TDSXX:4:2511:20618:17942 chr12 129539036 N chr12 129539155 N DUP 10
A00297:158:HT275DSXX:2:1576:8829:19319 chr12 129539024 N chr12 129539144 N DUP 12
A00404:155:HV27LDSXX:1:1634:24460:23124 chr12 129539036 N chr12 129539115 N DUP 14
A00404:156:HV37TDSXX:3:2613:11062:24064 chr12 129539036 N chr12 129539155 N DUP 10
A00404:156:HV37TDSXX:3:2613:11505:23860 chr12 129539036 N chr12 129539155 N DUP 10
A00297:158:HT275DSXX:3:1528:12418:14982 chr12 129539036 N chr12 129539115 N DUP 15
A00404:155:HV27LDSXX:4:2203:29541:21026 chr12 129538961 N chr12 129539080 N DUP 20
A00404:155:HV27LDSXX:2:2469:16776:36245 chr12 129539064 N chr12 129539144 N DUP 20
A00404:156:HV37TDSXX:3:1443:22164:14888 chr12 129539036 N chr12 129539115 N DUP 8
A00297:158:HT275DSXX:1:1311:27552:26318 chr12 129539036 N chr12 129539115 N DUP 2
A00297:158:HT275DSXX:1:2674:2166:6057 chr12 129539036 N chr12 129539115 N DUP 5
A00297:158:HT275DSXX:3:2563:8739:31908 chr12 129539036 N chr12 129539115 N DUP 2
A00404:156:HV37TDSXX:3:1664:24469:9204 chr12 129539050 N chr12 129539129 N DUP 10
A00297:158:HT275DSXX:3:1150:20690:33254 chr12 129539024 N chr12 129539144 N DUP 17
A00297:158:HT275DSXX:4:2476:6090:9251 chr12 129539036 N chr12 129539115 N DUP 5
A00404:155:HV27LDSXX:4:1531:19813:21590 chr12 129539024 N chr12 129539144 N DUP 17
A00404:155:HV27LDSXX:2:1106:16333:26678 chr12 129539050 N chr12 129539129 N DUP 10
A00404:156:HV37TDSXX:1:1108:3613:27759 chr12 129539036 N chr12 129539115 N DUP 4
A00297:158:HT275DSXX:2:2109:9824:13150 chr12 129539036 N chr12 129539115 N DUP 5
A00404:156:HV37TDSXX:2:1639:26268:17080 chr12 129539050 N chr12 129539129 N DUP 10
A00404:156:HV37TDSXX:3:1618:17029:35399 chr12 129538961 N chr12 129539080 N DUP 5
A00297:158:HT275DSXX:1:2672:27905:2503 chr12 129539050 N chr12 129539129 N DUP 10
A00297:158:HT275DSXX:1:2354:22327:23469 chr12 129539036 N chr12 129539115 N DUP 5
A00297:158:HT275DSXX:2:1659:3224:33129 chr12 129539036 N chr12 129539155 N DUP 15
A00297:158:HT275DSXX:4:2630:7256:5760 chr12 129538984 N chr12 129539144 N DUP 12
A00404:155:HV27LDSXX:1:2446:25997:17989 chr12 129539050 N chr12 129539129 N DUP 10
A00297:158:HT275DSXX:2:1341:32280:25645 chr12 129539064 N chr12 129539144 N DUP 17
A00404:155:HV27LDSXX:3:1655:22661:17691 chr12 129538961 N chr12 129539080 N DUP 5
A00297:158:HT275DSXX:4:1637:12156:24361 chr12 129539036 N chr12 129539115 N DUP 5
A00404:155:HV27LDSXX:3:2638:26377:18771 chr12 129539050 N chr12 129539129 N DUP 10
A00404:156:HV37TDSXX:4:2563:7717:20870 chr12 129539036 N chr12 129539115 N DUP 5
A00404:155:HV27LDSXX:4:2102:32298:18599 chr12 129539050 N chr12 129539129 N DUP 10
A00404:156:HV37TDSXX:2:1264:17607:34961 chr12 129539036 N chr12 129539155 N DUP 18
A00404:155:HV27LDSXX:3:1664:23204:11929 chr12 129539050 N chr12 129539129 N DUP 10
A00297:158:HT275DSXX:1:1623:16486:2519 chr12 129539036 N chr12 129539155 N DUP 16
A00404:156:HV37TDSXX:1:2565:6560:31798 chr12 129539050 N chr12 129539129 N DUP 11
A00404:156:HV37TDSXX:1:1557:24822:21872 chr12 129538961 N chr12 129539080 N DUP 20
A00404:155:HV27LDSXX:2:2541:22968:26209 chr12 129538984 N chr12 129539144 N DUP 13
A00297:158:HT275DSXX:3:2432:3839:31438 chr12 129538984 N chr12 129539144 N DUP 18
A00404:155:HV27LDSXX:1:2105:19397:34679 chr12 129539059 N chr12 129539140 N DEL 5
A00404:156:HV37TDSXX:4:1449:2410:23484 chr7 2459244 N chr7 2459570 N DUP 2
A00297:158:HT275DSXX:2:2333:29704:23187 chr7 2459244 N chr7 2459570 N DUP 2
A00404:155:HV27LDSXX:2:1335:26955:36401 chr7 2459261 N chr7 2459579 N DEL 3
A00297:158:HT275DSXX:3:2636:17861:5588 chr10 62369951 N chr10 62370716 N DEL 4
A00404:155:HV27LDSXX:4:1654:24044:18302 chr10 62369951 N chr10 62370716 N DEL 5
A00404:156:HV37TDSXX:2:2155:31774:8923 chr10 62369940 N chr10 62370339 N DEL 5
A00297:158:HT275DSXX:1:1625:20627:31328 chr10 62370009 N chr10 62370322 N DEL 1
A00297:158:HT275DSXX:3:1565:4996:28119 chr10 62370009 N chr10 62370322 N DEL 4
A00404:155:HV27LDSXX:3:1361:11225:36088 chr10 62370009 N chr10 62370322 N DEL 9
A00297:158:HT275DSXX:4:1169:3296:33285 chr10 62370009 N chr10 62370322 N DEL 9
A00297:158:HT275DSXX:4:1150:15962:26193 chr10 62369956 N chr10 62370037 N DUP 9
A00297:158:HT275DSXX:1:2356:11397:17065 chr10 62369956 N chr10 62370037 N DUP 9
A00404:156:HV37TDSXX:4:1638:1497:32612 chr10 62369940 N chr10 62370057 N DEL 4
A00404:156:HV37TDSXX:3:1453:10484:30671 chr10 62370058 N chr10 62370711 N DUP 1
A00404:155:HV27LDSXX:3:2603:1298:2581 chr10 62369981 N chr10 62370042 N DEL 7
A00404:155:HV27LDSXX:3:1413:25409:1658 chr10 62369956 N chr10 62370037 N DUP 7
A00404:155:HV27LDSXX:3:1350:6316:12430 chr10 62370049 N chr10 62370384 N DUP 7
A00297:158:HT275DSXX:4:2302:28619:26162 chr10 62370049 N chr10 62370384 N DUP 7
A00404:156:HV37TDSXX:3:2266:4191:35556 chr10 62370054 N chr10 62370361 N DUP 7
A00404:155:HV27LDSXX:1:2450:24225:9752 chr10 62369981 N chr10 62370042 N DEL 7
A00404:155:HV27LDSXX:2:1361:22589:34538 chr10 62369956 N chr10 62370009 N DUP 7
A00404:156:HV37TDSXX:2:2115:27335:21872 chr10 62369956 N chr10 62370009 N DUP 7
A00404:155:HV27LDSXX:3:1572:12545:36746 chr10 62369981 N chr10 62370042 N DEL 7
A00404:155:HV27LDSXX:4:2557:32660:2190 chr10 62369981 N chr10 62370042 N DEL 7
A00404:156:HV37TDSXX:2:2317:6967:35509 chr10 62369956 N chr10 62370037 N DUP 7
A00404:156:HV37TDSXX:2:2407:18783:8249 chr10 62369981 N chr10 62370042 N DEL 7
A00404:155:HV27LDSXX:3:2645:18150:10254 chr10 62370054 N chr10 62370361 N DUP 7
A00404:156:HV37TDSXX:1:2223:7283:36777 chr10 62370151 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:1:1639:18078:6120 chr10 62370037 N chr10 62370322 N DEL 7
A00404:156:HV37TDSXX:2:2374:7193:8625 chr10 62370057 N chr10 62370730 N DUP 2
A00404:155:HV27LDSXX:4:2259:11785:32706 chr10 62370151 N chr10 62370322 N DEL 7
A00404:156:HV37TDSXX:2:2268:30526:12023 chr10 62370037 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:3:1522:5186:30984 chr10 62370037 N chr10 62370322 N DEL 7
A00404:155:HV27LDSXX:1:2606:26756:4178 chr10 62370009 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:1:1556:7346:13870 chr10 62370009 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:3:1157:23556:19961 chr10 62370009 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:1:2447:3739:13260 chr10 62370037 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:1:2447:3748:13244 chr10 62370037 N chr10 62370322 N DEL 7
A00404:155:HV27LDSXX:2:2102:5403:27195 chr10 62370037 N chr10 62370322 N DEL 7
A00404:155:HV27LDSXX:2:2102:5755:27211 chr10 62370037 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:2:1247:27046:35430 chr10 62370037 N chr10 62370322 N DEL 7
A00404:156:HV37TDSXX:2:1632:23086:24126 chr10 62370037 N chr10 62370322 N DEL 7
A00404:156:HV37TDSXX:4:1320:21965:8500 chr10 62370047 N chr10 62370332 N DEL 7
A00404:155:HV27LDSXX:2:2149:26720:36025 chr10 62370037 N chr10 62370322 N DEL 7
A00404:155:HV27LDSXX:4:2411:5502:5572 chr10 62370037 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:2:1632:4806:35243 chr10 62370037 N chr10 62370322 N DEL 7
A00404:155:HV27LDSXX:1:1408:2510:23187 chr10 62370009 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:3:1266:7654:35728 chr10 62370009 N chr10 62370322 N DEL 7
A00404:156:HV37TDSXX:1:1438:30065:34491 chr10 62369981 N chr10 62370322 N DEL 7
A00404:156:HV37TDSXX:2:1632:23086:24126 chr10 62369981 N chr10 62370322 N DEL 7
A00297:158:HT275DSXX:4:1304:29740:24752 chr10 62369981 N chr10 62370322 N DEL 7
A00404:156:HV37TDSXX:4:2438:4580:3223 chr10 62370442 N chr10 62371227 N DEL 19
A00404:156:HV37TDSXX:4:1378:5593:9706 chr10 62370456 N chr10 62370520 N DEL 14
A00297:158:HT275DSXX:4:2619:29044:14246 chr10 62370442 N chr10 62370816 N DEL 14
A00404:155:HV27LDSXX:4:2259:11785:32706 chr10 62370419 N chr10 62370548 N DUP 3
A00404:155:HV27LDSXX:3:1577:25409:1470 chr10 62371177 N chr10 62371344 N DEL 19
A00404:155:HV27LDSXX:3:2650:24370:9565 chr10 62370470 N chr10 62370525 N DUP 6
A00404:155:HV27LDSXX:2:2278:27905:1438 chr10 62370667 N chr10 62371215 N DEL 4
A00404:155:HV27LDSXX:1:2265:5656:15076 chr10 62370773 N chr10 62370824 N DEL 1
A00404:155:HV27LDSXX:3:1668:19524:16767 chr10 62370707 N chr10 62370801 N DUP 13
A00404:155:HV27LDSXX:3:2668:16920:11569 chr10 62370707 N chr10 62370801 N DUP 13
A00404:155:HV27LDSXX:4:1566:18367:33990 chr10 62370707 N chr10 62370801 N DUP 13
A00297:158:HT275DSXX:2:2459:10203:3975 chr10 62370750 N chr10 62370828 N DUP 21
A00297:158:HT275DSXX:4:2209:24252:2159 chr10 62371037 N chr10 62371190 N DUP 27
A00404:155:HV27LDSXX:2:2163:18276:31704 chr10 62371032 N chr10 62371246 N DUP 19
A00404:155:HV27LDSXX:3:2539:30129:17848 chr10 62371128 N chr10 62371264 N DUP 34
A00404:155:HV27LDSXX:2:2602:1768:3897 chr10 62371212 N chr10 62371307 N DUP 13
A00297:158:HT275DSXX:4:2462:8693:11256 chr10 62371212 N chr10 62371307 N DUP 13
A00297:158:HT275DSXX:4:1469:23520:10535 chr10 62371209 N chr10 62371293 N DUP 36
A00404:155:HV27LDSXX:3:2162:9236:3051 chr10 62370823 N chr10 62371280 N DUP 1
A00404:156:HV37TDSXX:2:2313:1904:29841 chr10 62370440 N chr10 62371324 N DUP 7
A00404:156:HV37TDSXX:4:1261:21856:5932 chr10 62371160 N chr10 62371240 N DEL 1
A00404:155:HV27LDSXX:4:2553:14335:3051 chr10 62370440 N chr10 62371324 N DUP 7
A00297:158:HT275DSXX:4:2647:27751:31798 chr10 62370440 N chr10 62371324 N DUP 8
A00297:158:HT275DSXX:4:2462:8693:11256 chr10 62370436 N chr10 62371329 N DUP 17
A00404:155:HV27LDSXX:1:1239:27109:15843 chr10 62371227 N chr10 62371449 N DUP 23
A00404:156:HV37TDSXX:2:2313:1904:29841 chr10 62371350 N chr10 62371447 N DUP 29
A00297:158:HT275DSXX:1:2212:14796:35258 chr10 62371362 N chr10 62371499 N DEL 10
A00297:158:HT275DSXX:1:1454:19316:20071 chr10 62371362 N chr10 62371499 N DEL 9
A00404:156:HV37TDSXX:1:2147:5132:9815 chr10 62371362 N chr10 62371499 N DEL 9
A00297:158:HT275DSXX:3:2433:1389:13041 chr10 62370483 N chr10 62371471 N DEL 9
A00297:158:HT275DSXX:4:2351:14931:4366 chr10 62370792 N chr10 62371475 N DEL 8
A00404:156:HV37TDSXX:3:2101:5385:34397 chr10 62371347 N chr10 62371486 N DEL 5
A00404:155:HV27LDSXX:2:2450:17237:5666 chr10 62371362 N chr10 62371499 N DEL 19
A00297:158:HT275DSXX:4:1257:1895:34648 chr10 62371362 N chr10 62371499 N DEL 19
A00297:158:HT275DSXX:1:2447:30517:4492 chr10 62371367 N chr10 62371522 N DEL 21
A00404:155:HV27LDSXX:1:1542:14190:8030 chr10 62371368 N chr10 62371523 N DEL 21
A00297:158:HT275DSXX:2:2109:23357:25598 chr20 64287327 N chr20 64287529 N DUP 9
A00297:158:HT275DSXX:2:2256:24316:32205 chr20 64286944 N chr20 64287521 N DUP 14
A00404:156:HV37TDSXX:2:2516:5864:32941 chr20 64286943 N chr20 64287511 N DUP 16
A00404:155:HV27LDSXX:3:2609:12581:28573 chr20 64286943 N chr20 64287511 N DUP 13
A00404:155:HV27LDSXX:2:1367:8142:25207 chr20 64287074 N chr20 64287236 N DEL 5
A00404:156:HV37TDSXX:4:1139:21676:6684 chr20 64286960 N chr20 64287043 N DUP 14
A00297:158:HT275DSXX:1:2654:22833:36025 chr20 64287173 N chr20 64287284 N DEL 18
A00404:155:HV27LDSXX:1:2355:16414:25567 chr20 64287167 N chr20 64287327 N DEL 1
A00404:155:HV27LDSXX:2:2322:14425:17300 chr20 64286966 N chr20 64287354 N DEL 6
A00404:156:HV37TDSXX:4:2547:29713:9580 chr20 64286894 N chr20 64287457 N DUP 2
A00297:158:HT275DSXX:4:1664:25003:4805 chr20 64286867 N chr20 64287360 N DEL 6
A00404:155:HV27LDSXX:3:2331:23909:19225 chr20 64286931 N chr20 64287422 N DUP 6
A00404:155:HV27LDSXX:1:1465:22001:6339 chr20 64286858 N chr20 64287584 N DUP 6
A00404:155:HV27LDSXX:2:2136:6632:4773 chr20 64287290 N chr20 64287473 N DEL 12
A00404:155:HV27LDSXX:3:1573:15899:2785 chr20 64287488 N chr20 64287686 N DUP 6
A00404:155:HV27LDSXX:3:2529:24813:17378 chr20 64287291 N chr20 64287474 N DEL 7
A00404:156:HV37TDSXX:4:2513:25211:1564 chr20 64287457 N chr20 64287630 N DUP 32
A00297:158:HT275DSXX:1:1424:9769:29716 chr20 64287363 N chr20 64287580 N DEL 5
A00297:158:HT275DSXX:3:1510:8567:36025 chr20 64286940 N chr20 64287606 N DEL 3
A00404:156:HV37TDSXX:2:1233:6940:23563 chr20 64286927 N chr20 64287680 N DEL 15
A00297:158:HT275DSXX:3:2548:32696:8954 chr20 64287156 N chr20 64287660 N DEL 4
A00404:155:HV27LDSXX:2:2555:28248:31939 chr20 64286865 N chr20 64287673 N DEL 11
A00297:158:HT275DSXX:4:2315:8910:19304 chr20 64286866 N chr20 64287674 N DEL 10
A00297:158:HT275DSXX:3:1174:30825:33677 chr20 64287556 N chr20 64287726 N DEL 28
A00404:155:HV27LDSXX:1:1159:21766:35963 chr20 64286863 N chr20 64287683 N DEL 1
A00404:156:HV37TDSXX:2:1136:29460:9612 chr20 64286865 N chr20 64287679 N DEL 5
A00404:156:HV37TDSXX:2:1330:30273:4413 chr20 64287314 N chr20 64287748 N DEL 33
A00404:156:HV37TDSXX:1:1167:8052:9956 chr1 57290829 N chr1 57290984 N DEL 2
A00297:158:HT275DSXX:3:1676:14968:17519 chr1 57290829 N chr1 57290984 N DEL 5
A00404:155:HV27LDSXX:3:1518:2456:13823 chr1 57290829 N chr1 57290984 N DEL 5
A00297:158:HT275DSXX:1:2127:7527:25113 chr1 57290829 N chr1 57290984 N DEL 5
A00404:156:HV37TDSXX:2:2333:10185:14403 chr1 57290829 N chr1 57290984 N DEL 5
A00404:156:HV37TDSXX:2:2333:10402:13119 chr1 57290829 N chr1 57290984 N DEL 5
A00404:156:HV37TDSXX:4:2139:21432:33098 chr1 57290847 N chr1 57291000 N DUP 5
A00404:156:HV37TDSXX:2:2545:19171:22357 chr1 57290849 N chr1 57291002 N DUP 5
A00404:155:HV27LDSXX:4:1422:32922:30921 chr19 14362683 N chr19 14362810 N DEL 4
A00404:155:HV27LDSXX:3:2441:25518:10551 chr7 29263641 N chr7 29263758 N DEL 5
A00404:156:HV37TDSXX:1:2263:1488:27837 chr7 29263668 N chr7 29263785 N DEL 24
A00404:155:HV27LDSXX:2:2211:29577:16673 chr7 29263717 N chr7 29263834 N DEL 40
A00404:156:HV37TDSXX:2:1233:20618:30279 chr7 29263944 N chr7 29264368 N DEL 45
A00404:156:HV37TDSXX:3:1451:19723:16892 chr7 29264100 N chr7 29264210 N DEL 5
A00404:155:HV27LDSXX:2:2424:3206:26991 chr7 29264100 N chr7 29264210 N DEL 5
A00404:156:HV37TDSXX:1:1404:24858:8093 chr7 29264118 N chr7 29264226 N DUP 5
A00404:155:HV27LDSXX:3:2654:2826:7639 chr7 29264120 N chr7 29264228 N DUP 5
A00404:156:HV37TDSXX:1:2624:5990:26240 chr7 29264120 N chr7 29264228 N DUP 5
A00404:156:HV37TDSXX:1:1159:25120:9298 chr7 29264122 N chr7 29264230 N DUP 5
A00297:158:HT275DSXX:2:2643:18502:15781 chr7 29264123 N chr7 29264231 N DUP 5
A00404:155:HV27LDSXX:4:1162:21522:33254 chr7 29264221 N chr7 29264377 N DEL 31
A00404:155:HV27LDSXX:3:1611:15058:32925 chr7 29263602 N chr7 29264219 N DEL 1
A00404:155:HV27LDSXX:1:1654:26485:16078 chr7 29263789 N chr7 29264366 N DEL 6
A00404:155:HV27LDSXX:4:2507:13440:7200 chr7 29264288 N chr7 29264444 N DEL 5
A00297:158:HT275DSXX:4:1469:23005:30123 chr7 29264288 N chr7 29264444 N DEL 5
A00404:155:HV27LDSXX:2:2336:22218:8061 chr7 29264288 N chr7 29264444 N DEL 5
A00404:155:HV27LDSXX:3:1111:4345:28275 chr7 29264288 N chr7 29264444 N DEL 5
A00404:156:HV37TDSXX:4:1239:25699:18881 chr7 29264288 N chr7 29264444 N DEL 5
A00404:155:HV27LDSXX:2:1574:7563:7795 chr7 29263790 N chr7 29264444 N DEL 5
A00404:155:HV27LDSXX:1:2134:20537:4272 chr7 29263790 N chr7 29264444 N DEL 5
A00404:156:HV37TDSXX:1:1274:14271:26334 chr7 29263790 N chr7 29264444 N DEL 5
A00404:156:HV37TDSXX:1:1274:14470:26772 chr7 29263790 N chr7 29264444 N DEL 5
A00404:156:HV37TDSXX:1:1274:14470:26804 chr7 29263790 N chr7 29264444 N DEL 5
A00404:155:HV27LDSXX:3:1140:10682:36276 chr1 13038079 N chr1 13038201 N DEL 13
A00404:156:HV37TDSXX:1:2657:32542:34491 chr1 13038075 N chr1 13038201 N DEL 12
A00404:156:HV37TDSXX:3:2669:29324:29857 chr21 46069103 N chr21 46069438 N DEL 8
A00404:155:HV27LDSXX:3:1550:29342:36432 chr21 46069507 N chr21 46069588 N DUP 4
A00404:155:HV27LDSXX:3:1320:27624:6339 chr21 46069510 N chr21 46069591 N DUP 1
A00404:156:HV37TDSXX:4:2423:26015:27258 chr7 113712956 N chr7 113713035 N DEL 9
A00297:158:HT275DSXX:4:2138:8630:12023 chr7 113712956 N chr7 113713035 N DEL 9
A00297:158:HT275DSXX:1:1309:23565:17347 chr7 113712956 N chr7 113713035 N DEL 9
A00404:155:HV27LDSXX:3:1235:4237:5666 chr7 113712956 N chr7 113713035 N DEL 9
A00404:156:HV37TDSXX:4:1166:15194:13307 chr7 113712956 N chr7 113713035 N DEL 9
A00404:155:HV27LDSXX:2:2414:2446:34413 chr7 113712956 N chr7 113713035 N DEL 9
A00297:158:HT275DSXX:2:2560:14615:29434 chr7 113712872 N chr7 113713043 N DEL 7
A00297:158:HT275DSXX:2:2560:14687:29496 chr7 113712872 N chr7 113713043 N DEL 7
A00404:155:HV27LDSXX:4:2447:1669:16752 chr7 101113451 N chr7 101113518 N DEL 5
A00404:155:HV27LDSXX:1:2219:3414:20055 chr17 78893544 N chr17 78893603 N DEL 5
A00404:155:HV27LDSXX:3:1334:25861:3505 chr17 78893292 N chr17 78893563 N DEL 5
A00404:156:HV37TDSXX:2:1263:27552:28604 chr17 78893292 N chr17 78893563 N DEL 5
A00404:156:HV37TDSXX:2:2468:7717:10723 chr17 78893292 N chr17 78893563 N DEL 5
A00404:156:HV37TDSXX:1:1473:32976:20744 chr21 32507940 N chr21 32508076 N DUP 1
A00404:155:HV27LDSXX:2:1376:7374:33238 chr4 14836515 N chr4 14836594 N DEL 5
A00297:158:HT275DSXX:4:2164:4155:25504 chr4 14836524 N chr4 14837396 N DEL 1
A00404:156:HV37TDSXX:4:1455:9155:4476 chr4 14836524 N chr4 14837396 N DEL 1
A00404:156:HV37TDSXX:1:1547:4517:34992 chr4 14836524 N chr4 14837396 N DEL 2
A00297:158:HT275DSXX:1:1260:18114:37027 chr4 14836535 N chr4 14837389 N DEL 3
A00404:156:HV37TDSXX:4:2603:24053:25739 chr4 14836691 N chr4 14836771 N DUP 23
A00404:155:HV27LDSXX:3:1112:7726:36448 chr4 14836584 N chr4 14836818 N DUP 14
A00404:155:HV27LDSXX:3:1112:7925:36573 chr4 14836584 N chr4 14836818 N DUP 14
A00404:155:HV27LDSXX:3:1112:9019:36620 chr4 14836584 N chr4 14836818 N DUP 14
A00404:156:HV37TDSXX:2:2140:19271:23563 chr4 14836655 N chr4 14836762 N DUP 10
A00404:156:HV37TDSXX:4:1370:6741:15233 chr4 14836597 N chr4 14836772 N DUP 18
A00404:156:HV37TDSXX:2:2316:28872:6997 chr4 14836691 N chr4 14836771 N DUP 23
A00404:156:HV37TDSXX:3:2135:27299:30702 chr4 14836691 N chr4 14836771 N DUP 23
A00297:158:HT275DSXX:2:1640:5104:28526 chr4 14836691 N chr4 14836771 N DUP 22
A00297:158:HT275DSXX:4:2631:5077:26694 chr4 14836691 N chr4 14836771 N DUP 22
A00404:155:HV27LDSXX:3:1373:3369:6918 chr4 14836691 N chr4 14836771 N DUP 22
A00404:156:HV37TDSXX:1:1473:20302:13448 chr4 14836691 N chr4 14836771 N DUP 22
A00404:156:HV37TDSXX:1:1246:27489:14810 chr4 14836691 N chr4 14836771 N DUP 21
A00297:158:HT275DSXX:2:1609:16803:7921 chr4 14836631 N chr4 14836700 N DEL 19
A00404:155:HV27LDSXX:4:2629:20329:7420 chr4 14836691 N chr4 14836771 N DUP 24
A00404:156:HV37TDSXX:1:2317:22507:35336 chr4 14836691 N chr4 14836771 N DUP 24
A00404:155:HV27LDSXX:4:2608:7482:20306 chr4 14836691 N chr4 14836771 N DUP 24
A00297:158:HT275DSXX:2:1157:7527:13777 chr4 14836703 N chr4 14836754 N DUP 26
A00297:158:HT275DSXX:2:2531:15817:6214 chr4 14836715 N chr4 14836812 N DUP 17
A00404:155:HV27LDSXX:4:2423:23511:15311 chr4 14837251 N chr4 14837556 N DEL 10
A00404:155:HV27LDSXX:4:2423:24198:12931 chr4 14837251 N chr4 14837556 N DEL 10
A00297:158:HT275DSXX:1:1238:26142:15201 chr4 14837185 N chr4 14837578 N DUP 11
A00404:156:HV37TDSXX:2:1350:20772:28792 chr4 14837127 N chr4 14837559 N DUP 31
A00297:158:HT275DSXX:3:1543:22607:6511 chr4 14837022 N chr4 14837351 N DUP 2
A00404:156:HV37TDSXX:3:1413:27877:27602 chr4 14837169 N chr4 14837296 N DUP 9
A00297:158:HT275DSXX:3:1523:18050:10050 chr4 14837308 N chr4 14837437 N DUP 10
A00297:158:HT275DSXX:3:1523:20446:12164 chr4 14837308 N chr4 14837437 N DUP 10
A00297:158:HT275DSXX:2:1538:17716:2049 chr4 14837556 N chr4 14837636 N DUP 17
A00404:156:HV37TDSXX:3:1526:10330:20322 chr4 14837131 N chr4 14837415 N DUP 11
A00404:156:HV37TDSXX:3:1526:10330:20322 chr4 14836569 N chr4 14837584 N DEL 17
A00404:156:HV37TDSXX:3:1560:2935:20603 chr4 14837535 N chr4 14837623 N DEL 21
A00297:158:HT275DSXX:2:2422:14877:14763 chr4 14836765 N chr4 14837627 N DEL 11
A00404:156:HV37TDSXX:3:1236:28492:22654 chr4 14836766 N chr4 14837628 N DEL 10
A00297:158:HT275DSXX:3:1533:3152:15718 chr10 119360139 N chr10 119360237 N DEL 9
A00297:158:HT275DSXX:1:1367:6370:14779 chr19 52907096 N chr19 52907433 N DEL 1
A00297:158:HT275DSXX:1:1131:2591:3474 chr19 52906885 N chr19 52907220 N DUP 1
A00297:158:HT275DSXX:1:1210:23276:22044 chr19 52906933 N chr19 52907270 N DEL 10
A00297:158:HT275DSXX:2:1420:26178:26944 chr19 52906933 N chr19 52907270 N DEL 10
A00404:155:HV27LDSXX:2:2422:28709:12759 chr19 52906667 N chr19 52907256 N DEL 5
A00404:156:HV37TDSXX:2:2461:11840:15859 chr19 52907130 N chr19 52907467 N DEL 10
A00297:158:HT275DSXX:1:2268:8684:22576 chr19 52907109 N chr19 52907446 N DEL 2
A00404:155:HV27LDSXX:4:2311:18295:19085 chr1 212749563 N chr1 212749641 N DEL 4
A00404:155:HV27LDSXX:1:1648:30355:9909 chr9 43346512 N chr9 43346632 N DUP 5
A00404:156:HV37TDSXX:1:1349:6596:31266 chr7 67385838 N chr7 67386004 N DEL 20
A00404:156:HV37TDSXX:4:1340:25220:1830 chr11 88359181 N chr11 88359351 N DUP 10
A00404:156:HV37TDSXX:4:2247:26395:32299 chr11 88359183 N chr11 88359353 N DUP 8
A00404:155:HV27LDSXX:4:2251:2347:8218 chr5 930828 N chr5 931053 N DEL 6
A00404:156:HV37TDSXX:1:2211:17336:6590 chr10 45870076 N chr10 45870294 N DEL 17
A00297:158:HT275DSXX:2:1317:26775:29982 chr18 79339392 N chr18 79339591 N DEL 10
A00404:155:HV27LDSXX:3:2635:3034:5525 chr18 79339392 N chr18 79339591 N DEL 12
A00297:158:HT275DSXX:1:2448:21169:5368 chr18 79339392 N chr18 79339591 N DEL 12
A00404:155:HV27LDSXX:1:1428:31458:26694 chr18 79339315 N chr18 79339408 N DEL 5
A00404:156:HV37TDSXX:3:1151:2971:15342 chr18 79339317 N chr18 79339410 N DEL 5
A00404:156:HV37TDSXX:3:1151:3477:13056 chr18 79339317 N chr18 79339410 N DEL 5
A00404:155:HV27LDSXX:3:1461:16333:12461 chr18 79339417 N chr18 79339637 N DUP 2
A00404:155:HV27LDSXX:3:2460:17508:27336 chr18 79339417 N chr18 79339637 N DUP 2
A00297:158:HT275DSXX:2:2376:24840:11694 chr16 50755268 N chr16 50755351 N DEL 5
A00404:156:HV37TDSXX:3:1323:9471:19805 chr16 80243533 N chr16 80244138 N DEL 5
A00404:156:HV37TDSXX:3:1323:9471:19805 chr16 80243527 N chr16 80244132 N DEL 15
A00297:158:HT275DSXX:4:1638:22507:22404 chr16 80243546 N chr16 80244151 N DEL 14
A00404:156:HV37TDSXX:2:2359:5565:1705 chr16 80243591 N chr16 80244325 N DEL 5
A00404:155:HV27LDSXX:2:1349:26612:6997 chr16 80243659 N chr16 80244340 N DEL 5
A00404:155:HV27LDSXX:1:1342:12454:6778 chr16 80243555 N chr16 80243653 N DEL 1
A00404:155:HV27LDSXX:2:1435:9733:15248 chr16 80243720 N chr16 80244048 N DEL 20
A00404:156:HV37TDSXX:3:1358:16405:30655 chr16 80243797 N chr16 80243896 N DEL 5
A00297:158:HT275DSXX:1:1323:27263:14982 chr16 80243758 N chr16 80244211 N DUP 1
A00297:158:HT275DSXX:2:2550:21766:2143 chr16 80243816 N chr16 80244269 N DUP 10
A00404:155:HV27LDSXX:2:1349:26612:6997 chr16 80243811 N chr16 80244363 N DUP 8
A00297:158:HT275DSXX:2:2160:29125:20995 chr16 80243550 N chr16 80243828 N DEL 9
A00404:156:HV37TDSXX:1:2219:4698:26506 chr16 80244028 N chr16 80244284 N DEL 5
A00404:156:HV37TDSXX:2:1577:3531:28369 chr16 80243704 N chr16 80244030 N DUP 5
A00404:156:HV37TDSXX:2:1577:3531:28369 chr16 80243831 N chr16 80244030 N DUP 5
A00297:158:HT275DSXX:4:2223:12807:14967 chr16 80244030 N chr16 80244159 N DEL 11
A00404:155:HV27LDSXX:2:1619:3586:17002 chr16 80243704 N chr16 80244030 N DUP 5
A00404:155:HV27LDSXX:2:1631:7672:35759 chr16 80243558 N chr16 80243983 N DEL 1
A00297:158:HT275DSXX:3:1222:31015:15029 chr16 80244072 N chr16 80244377 N DEL 5
A00404:155:HV27LDSXX:1:2101:1624:6809 chr16 80243534 N chr16 80244137 N DUP 5
A00404:156:HV37TDSXX:4:2350:30662:10848 chr16 80244150 N chr16 80244328 N DEL 10
A00404:156:HV37TDSXX:2:2520:9607:9674 chr16 80243823 N chr16 80244151 N DEL 5
A00297:158:HT275DSXX:2:2160:29125:20995 chr16 80244278 N chr16 80244329 N DEL 18
A00404:156:HV37TDSXX:2:2210:28700:22388 chr16 80244157 N chr16 80244335 N DEL 5
A00404:155:HV27LDSXX:1:2321:29270:3427 chr16 80243629 N chr16 80244363 N DEL 5
A00404:156:HV37TDSXX:1:1127:19678:5447 chr16 80244081 N chr16 80244386 N DEL 19
A00297:158:HT275DSXX:3:1611:10285:22717 chr16 80244083 N chr16 80244388 N DEL 9
A00404:156:HV37TDSXX:2:2306:3721:5212 chr1 58518379 N chr1 58518437 N DEL 20
A00404:155:HV27LDSXX:2:1323:10926:4319 chr1 58518453 N chr1 58518504 N DEL 5
A00297:158:HT275DSXX:1:2462:16188:32628 chr1 58518453 N chr1 58518504 N DEL 5
A00404:155:HV27LDSXX:4:2433:4535:34554 chr1 58518453 N chr1 58518504 N DEL 5
A00404:155:HV27LDSXX:3:1129:7717:32925 chr1 58518448 N chr1 58518504 N DEL 5
A00404:155:HV27LDSXX:4:2232:4472:11647 chr1 58518441 N chr1 58518507 N DEL 5
A00404:155:HV27LDSXX:4:2232:4490:12054 chr1 58518441 N chr1 58518507 N DEL 5
A00404:156:HV37TDSXX:1:1341:6958:13166 chr2 91498248 N chr2 91498333 N DEL 5
A00297:158:HT275DSXX:2:2273:24650:14058 chr2 91498242 N chr2 91498353 N DUP 5
A00404:156:HV37TDSXX:4:1575:4155:31454 chr2 91498419 N chr2 91498529 N DEL 6
A00297:158:HT275DSXX:2:2233:32633:17989 chr2 91498419 N chr2 91498529 N DEL 6
A00404:155:HV27LDSXX:4:1360:10257:13902 chr2 91498597 N chr2 91498651 N DEL 9
A00297:158:HT275DSXX:4:2524:3803:34319 chr2 91498442 N chr2 91498544 N DEL 4
A00404:155:HV27LDSXX:4:1309:17571:9126 chr6 5035696 N chr6 5035936 N DEL 6
A00404:156:HV37TDSXX:1:1262:16179:11318 chr19 7419201 N chr19 7419409 N DEL 5
A00404:155:HV27LDSXX:4:1412:20130:32659 chr10 1375997 N chr10 1376121 N DUP 5
A00297:158:HT275DSXX:4:2153:19379:28541 chr10 1375957 N chr10 1376122 N DUP 5
A00297:158:HT275DSXX:4:2153:20772:29418 chr10 1375957 N chr10 1376122 N DUP 5
A00404:156:HV37TDSXX:3:2475:15176:34381 chr10 1376010 N chr10 1376136 N DEL 5
A00404:155:HV27LDSXX:3:2636:22444:13056 chr10 1375975 N chr10 1376142 N DEL 5
A00404:156:HV37TDSXX:2:2322:19651:3803 chr21 23807802 N chr21 23807853 N DEL 5
A00404:155:HV27LDSXX:2:1428:13838:27618 chr21 23807802 N chr21 23807853 N DEL 5
A00404:156:HV37TDSXX:4:1607:3676:21981 chr21 23807802 N chr21 23807853 N DEL 6
A00404:155:HV27LDSXX:2:1213:6063:27336 chr21 23807802 N chr21 23807853 N DEL 10
A00297:158:HT275DSXX:2:1305:25834:13949 chr21 23807802 N chr21 23807853 N DEL 17
A00404:155:HV27LDSXX:1:2277:11749:25254 chr21 23807802 N chr21 23807853 N DEL 18
A00404:155:HV27LDSXX:1:2277:7075:14372 chr21 23807802 N chr21 23807853 N DEL 18
A00297:158:HT275DSXX:4:1630:11794:14309 chr21 23807802 N chr21 23807853 N DEL 19
A00404:156:HV37TDSXX:1:2602:5737:32753 chr21 23807802 N chr21 23807853 N DEL 23
A00404:156:HV37TDSXX:2:1464:12237:2018 chr21 23807802 N chr21 23807853 N DEL 30
A00404:155:HV27LDSXX:4:1227:7753:10942 chr21 23807802 N chr21 23807853 N DEL 33
A00404:155:HV27LDSXX:2:2130:27028:23469 chr21 23807802 N chr21 23807853 N DEL 39
A00404:156:HV37TDSXX:1:1375:17824:21496 chr21 23807802 N chr21 23807853 N DEL 40
A00297:158:HT275DSXX:4:1106:18457:25191 chr14 106531010 N chr14 106531068 N DEL 5
A00404:155:HV27LDSXX:4:2667:22408:11146 chr14 106531010 N chr14 106531145 N DEL 5
A00404:155:HV27LDSXX:1:1440:5448:25989 chr17 2268769 N chr17 2268902 N DUP 4
A00297:158:HT275DSXX:2:1506:4598:4351 chr20 33701351 N chr20 33701507 N DEL 45
A00297:158:HT275DSXX:4:2543:4029:15452 chr1 12274514 N chr1 12274651 N DEL 14
A00404:155:HV27LDSXX:3:1616:11360:4758 chr6 52825449 N chr6 52825902 N DEL 5
A00404:155:HV27LDSXX:2:1660:15772:31344 chr6 52825417 N chr6 52825684 N DEL 32
A00404:155:HV27LDSXX:2:1660:15790:31344 chr6 52825417 N chr6 52825684 N DEL 32
A00404:155:HV27LDSXX:2:1544:17915:27539 chr6 52825556 N chr6 52825785 N DEL 17
A00404:155:HV27LDSXX:1:2307:16712:34851 chr6 52825805 N chr6 52825880 N DEL 5
A00297:158:HT275DSXX:1:2223:29423:7451 chr6 52825693 N chr6 52825843 N DUP 5
A00404:156:HV37TDSXX:1:2239:29071:17989 chr6 52825693 N chr6 52825843 N DUP 5
A00297:158:HT275DSXX:1:2163:19669:31641 chr6 52825620 N chr6 52825809 N DEL 5
A00297:158:HT275DSXX:1:2166:22209:3724 chr6 52825620 N chr6 52825809 N DEL 5
A00404:156:HV37TDSXX:2:2102:32542:23030 chr6 52825622 N chr6 52825811 N DEL 5
A00297:158:HT275DSXX:4:1603:29821:37012 chr6 52825619 N chr6 52825845 N DEL 5
A00297:158:HT275DSXX:4:1426:24813:4069 chr6 52825643 N chr6 52825869 N DEL 2
A00404:155:HV27LDSXX:2:1544:17915:27539 chr6 52825643 N chr6 52825869 N DEL 2
A00404:156:HV37TDSXX:3:2158:25048:26334 chr6 52825683 N chr6 52825909 N DEL 35
A00404:155:HV27LDSXX:1:1578:10086:11882 chr6 52825494 N chr6 52825947 N DEL 5
A00404:155:HV27LDSXX:4:1459:24560:25989 chr1 186307104 N chr1 186307813 N DEL 19
A00404:155:HV27LDSXX:1:2448:20853:19476 chr1 186307070 N chr1 186307188 N DEL 5
A00297:158:HT275DSXX:2:2321:31168:35681 chr1 186307258 N chr1 186307536 N DUP 10
A00404:155:HV27LDSXX:4:2202:19244:6825 chr1 186307387 N chr1 186307526 N DEL 7
A00404:155:HV27LDSXX:1:1364:22625:20697 chr1 186307540 N chr1 186307805 N DEL 11
A00404:156:HV37TDSXX:2:2102:29948:4946 chr1 186307024 N chr1 186307491 N DUP 5
A00404:156:HV37TDSXX:1:1268:14977:9079 chr1 186307584 N chr1 186308041 N DEL 1
A00404:155:HV27LDSXX:1:2159:27905:26647 chr1 186307060 N chr1 186307532 N DEL 13
A00297:158:HT275DSXX:4:2372:1344:35102 chr1 186307932 N chr1 186308116 N DEL 9
A00297:158:HT275DSXX:2:2428:1696:9345 chr1 186307696 N chr1 186307983 N DUP 8
A00404:155:HV27LDSXX:1:1363:17644:10254 chr1 186307201 N chr1 186308142 N DUP 7
A00404:156:HV37TDSXX:4:1369:29812:17863 chr17 62123119 N chr17 62123218 N DEL 9
A00404:156:HV37TDSXX:3:1554:7274:33129 chr17 62123092 N chr17 62123218 N DEL 9
A00404:155:HV27LDSXX:4:2641:10402:13182 chr17 62123194 N chr17 62123300 N DEL 6
A00404:155:HV27LDSXX:4:2641:10411:13166 chr17 62123194 N chr17 62123300 N DEL 6
A00404:155:HV27LDSXX:3:2263:25753:27837 chr6 132384364 N chr6 132384433 N DUP 6
A00297:158:HT275DSXX:4:2420:24994:26021 chr6 132384364 N chr6 132384433 N DUP 6
A00404:156:HV37TDSXX:3:1347:12201:12164 chr10 131890568 N chr10 131890755 N DEL 5
A00404:156:HV37TDSXX:4:1443:26702:12978 chr10 131890702 N chr10 131890785 N DEL 1
A00404:155:HV27LDSXX:3:1525:5439:31610 chr10 131890724 N chr10 131890927 N DUP 5
A00404:156:HV37TDSXX:4:1621:19162:28823 chr4 174405113 N chr4 174405279 N DEL 3
A00404:155:HV27LDSXX:2:2237:7636:33473 chr12 66068995 N chr12 66069481 N DEL 4
A00404:156:HV37TDSXX:4:2362:2293:21402 chr12 66069072 N chr12 66069237 N DEL 11
A00404:155:HV27LDSXX:3:2122:13720:35055 chr12 66068986 N chr12 66069062 N DEL 13
A00404:155:HV27LDSXX:4:2215:22399:22247 chr12 66068986 N chr12 66069062 N DEL 16
A00297:158:HT275DSXX:2:1166:13295:14027 chr12 66068943 N chr12 66069006 N DEL 5
A00404:155:HV27LDSXX:3:1375:15121:33004 chr12 66068948 N chr12 66069011 N DEL 3
A00297:158:HT275DSXX:4:2646:23647:34741 chr12 66068947 N chr12 66069010 N DEL 4
A00297:158:HT275DSXX:4:2646:24731:35086 chr12 66068947 N chr12 66069010 N DEL 4
A00404:156:HV37TDSXX:4:2560:19931:26459 chr12 66068875 N chr12 66069110 N DEL 1
A00404:155:HV27LDSXX:4:1470:24487:1313 chr12 66069268 N chr12 66069361 N DEL 2
A00404:155:HV27LDSXX:1:1551:19099:13964 chr12 66068980 N chr12 66069276 N DUP 9
A00404:156:HV37TDSXX:1:1462:2031:8328 chr12 66069170 N chr12 66069256 N DUP 5
A00404:155:HV27LDSXX:3:1426:27516:34773 chr12 66068852 N chr12 66069543 N DUP 9
A00404:155:HV27LDSXX:3:2249:6180:13542 chr12 66068852 N chr12 66069616 N DUP 5
A00404:155:HV27LDSXX:4:2159:17318:11256 chr12 66068852 N chr12 66069591 N DUP 8
A00404:156:HV37TDSXX:4:2107:25256:7341 chr12 66069603 N chr12 66069677 N DUP 21
A00404:155:HV27LDSXX:4:2321:14651:26929 chr12 66069603 N chr12 66069677 N DUP 22
A00404:156:HV37TDSXX:3:1172:20889:9173 chr12 66069603 N chr12 66069677 N DUP 15
A00297:158:HT275DSXX:2:1526:10710:4288 chr12 66068876 N chr12 66069569 N DEL 10
A00404:155:HV27LDSXX:1:1604:23393:2863 chr12 66069603 N chr12 66069677 N DUP 19
A00297:158:HT275DSXX:1:2316:25256:12571 chr12 66068876 N chr12 66069569 N DEL 9
A00404:156:HV37TDSXX:4:2665:20971:30044 chr12 66069603 N chr12 66069652 N DUP 11
A00404:155:HV27LDSXX:4:2353:7844:16861 chr12 66069603 N chr12 66069677 N DUP 12
A00297:158:HT275DSXX:3:1544:18738:9925 chr12 66069603 N chr12 66069677 N DUP 12
A00404:156:HV37TDSXX:1:1544:21197:27680 chr12 66068877 N chr12 66069693 N DEL 5
A00404:155:HV27LDSXX:1:2159:29613:6527 chr12 66068905 N chr12 66069694 N DEL 5
A00404:155:HV27LDSXX:1:2159:30481:15013 chr12 66068905 N chr12 66069694 N DEL 5
A00404:156:HV37TDSXX:1:2429:18692:6746 chr14 42650141 N chr14 42650190 N DUP 10
A00404:155:HV27LDSXX:3:1421:26223:5603 chr14 42650141 N chr14 42650190 N DUP 10
A00297:158:HT275DSXX:4:1631:8721:24799 chr17 80160265 N chr17 80160358 N DEL 10
A00404:156:HV37TDSXX:2:2367:27073:10802 chr19 47991828 N chr19 47992043 N DEL 56
A00297:158:HT275DSXX:1:2615:10628:36464 chr16 2857146 N chr16 2857499 N DEL 10
A00297:158:HT275DSXX:1:2658:20799:19319 chr16 2857157 N chr16 2857556 N DEL 5
A00297:158:HT275DSXX:1:2369:30843:34366 chr16 2857339 N chr16 2857531 N DEL 2
A00404:156:HV37TDSXX:1:2566:24252:36699 chr16 2857348 N chr16 2857421 N DEL 5
A00404:155:HV27LDSXX:1:1473:28330:33019 chr16 2857387 N chr16 2857530 N DUP 13
A00297:158:HT275DSXX:4:2623:19180:5337 chr16 2857355 N chr16 2857476 N DEL 5
A00297:158:HT275DSXX:2:2147:7292:28213 chr16 2857175 N chr16 2857481 N DEL 11
A00404:155:HV27LDSXX:2:2503:19099:8296 chr16 2857177 N chr16 2857482 N DEL 5
A00297:158:HT275DSXX:4:2101:17707:14559 chr16 2857179 N chr16 2857554 N DEL 17
A00297:158:HT275DSXX:4:1359:9317:6167 chr21 45376161 N chr21 45376320 N DEL 8
A00404:155:HV27LDSXX:4:1232:27172:22811 chr21 45376093 N chr21 45376225 N DUP 5
A00297:158:HT275DSXX:4:1359:9317:6167 chr21 45376114 N chr21 45376212 N DEL 5
A00404:156:HV37TDSXX:2:1210:19768:17409 chr16 56580929 N chr16 56581014 N DUP 5
A00404:156:HV37TDSXX:4:1232:9218:2018 chr16 56580929 N chr16 56581014 N DUP 11
A00404:155:HV27LDSXX:1:1219:5945:25629 chr16 56580929 N chr16 56581014 N DUP 14
A00297:158:HT275DSXX:2:1429:12183:29637 chr16 56580927 N chr16 56581019 N DEL 10
A00404:156:HV37TDSXX:3:2267:27335:35775 chr18 48180079 N chr18 48180274 N DEL 3
A00404:156:HV37TDSXX:2:1524:10764:10019 chr18 48180144 N chr18 48180319 N DEL 5
A00297:158:HT275DSXX:3:1217:9263:19727 chr18 48180030 N chr18 48180335 N DEL 13
A00297:158:HT275DSXX:2:2435:21251:34538 chr22 45981015 N chr22 45981269 N DUP 5
A00404:155:HV27LDSXX:3:2327:21296:18771 chr22 45981043 N chr22 45981265 N DEL 14
A00404:155:HV27LDSXX:3:2519:12020:27602 chr8 141488172 N chr8 141488267 N DEL 5
A00297:158:HT275DSXX:3:2634:30101:11381 chr8 141488198 N chr8 141488291 N DUP 5
A00297:158:HT275DSXX:2:2332:9408:35978 chr8 141488206 N chr8 141488299 N DUP 5
A00404:155:HV27LDSXX:1:1552:30906:12054 chr14 105186475 N chr14 105186612 N DEL 5
A00297:158:HT275DSXX:4:1331:12599:26162 chr14 105187025 N chr14 105187076 N DUP 10
A00297:158:HT275DSXX:4:2210:1913:28197 chr14 105187027 N chr14 105187078 N DUP 10
A00404:155:HV27LDSXX:2:2272:16215:28604 chr14 105187218 N chr14 105187344 N DEL 12
A00297:158:HT275DSXX:2:2340:20166:7263 chr4 24493415 N chr4 24493490 N DUP 3
A00404:155:HV27LDSXX:1:2132:11623:6214 chr7 84791764 N chr7 84791817 N DEL 3
A00404:155:HV27LDSXX:2:1555:6036:30577 chrY 11017322 N chrY 11017396 N DUP 5
A00404:155:HV27LDSXX:3:2261:21368:9815 chrY 11017322 N chrY 11017396 N DUP 5
A00404:155:HV27LDSXX:3:1640:32452:25567 chrY 11017322 N chrY 11017396 N DUP 69
A00404:155:HV27LDSXX:3:1640:32452:25567 chrY 11017322 N chrY 11017396 N DUP 71
A00404:156:HV37TDSXX:1:1476:17137:15515 chrY 11017389 N chrY 11017521 N DEL 5
A00404:155:HV27LDSXX:2:2248:1344:30624 chrY 11017379 N chrY 11017521 N DEL 5
A00404:156:HV37TDSXX:1:2442:28483:37012 chrY 11017322 N chrY 11017395 N DUP 15
A00404:155:HV27LDSXX:3:2220:25120:16532 chrY 11017339 N chrY 11017521 N DEL 5
A00404:156:HV37TDSXX:3:1676:31783:23156 chrY 11017336 N chrY 11017522 N DEL 5
A00404:156:HV37TDSXX:1:1627:12843:4351 chrY 11017336 N chrY 11017522 N DEL 5
A00404:156:HV37TDSXX:1:1627:13783:3035 chrY 11017336 N chrY 11017522 N DEL 5
A00297:158:HT275DSXX:3:1229:6171:29027 chrY 11017336 N chrY 11017524 N DEL 5
A00404:155:HV27LDSXX:3:2156:19072:26475 chrY 11017360 N chrY 11017581 N DEL 5
A00404:156:HV37TDSXX:3:1615:32497:29590 chrY 11017355 N chrY 11017644 N DEL 10
A00404:155:HV27LDSXX:3:2156:19072:26475 chrY 11017322 N chrY 11017396 N DUP 70
A00404:156:HV37TDSXX:2:1141:27715:31078 chrY 11017322 N chrY 11017396 N DUP 9
A00404:156:HV37TDSXX:2:1666:4598:23015 chrY 11017322 N chrY 11017396 N DUP 67
A00297:158:HT275DSXX:4:1334:2700:16188 chrY 11017322 N chrY 11017394 N DUP 71
A00404:155:HV27LDSXX:2:1427:30120:2362 chrY 11017322 N chrY 11017395 N DUP 71
A00404:156:HV37TDSXX:3:2373:14253:10238 chrY 11017322 N chrY 11017395 N DUP 71
A00404:156:HV37TDSXX:4:1515:25220:17300 chrY 11017322 N chrY 11017396 N DUP 71
A00404:155:HV27LDSXX:4:1575:18783:36777 chrY 11017322 N chrY 11017395 N DUP 68
A00404:155:HV27LDSXX:4:1343:20428:35618 chrY 11017322 N chrY 11017396 N DUP 71
A00404:156:HV37TDSXX:2:2574:13141:9189 chrY 11017322 N chrY 11017396 N DUP 71
A00404:155:HV27LDSXX:4:1424:32633:31454 chrY 11017322 N chrY 11017396 N DUP 71
A00297:158:HT275DSXX:2:1210:12292:8469 chrY 11017322 N chrY 11017396 N DUP 71
A00404:155:HV27LDSXX:3:1348:6298:20603 chrY 11017322 N chrY 11017396 N DUP 71
A00404:155:HV27LDSXX:2:1608:21974:9987 chrY 11017322 N chrY 11017396 N DUP 71
A00297:158:HT275DSXX:1:2373:23493:14309 chrY 11017336 N chrY 11017784 N DEL 3
A00404:156:HV37TDSXX:3:1676:31783:23156 chrY 11017322 N chrY 11017396 N DUP 45
A00404:156:HV37TDSXX:1:1614:7627:11130 chrY 11017322 N chrY 11017396 N DUP 25
A00297:158:HT275DSXX:3:2518:21856:4085 chr16 46382709 N chr16 46382855 N DUP 4
A00297:158:HT275DSXX:4:1156:4092:23547 chr16 46382709 N chr16 46382855 N DUP 4
A00404:155:HV27LDSXX:1:1270:8386:21590 chr16 46382709 N chr16 46382855 N DUP 4
A00404:155:HV27LDSXX:2:1146:4074:11303 chr16 46382709 N chr16 46382855 N DUP 4
A00404:155:HV27LDSXX:2:1331:11740:4069 chr16 46382711 N chr16 46382782 N DUP 2
A00404:155:HV27LDSXX:2:1627:28908:27320 chr16 46382709 N chr16 46382855 N DUP 4
A00404:155:HV27LDSXX:2:2313:29378:7435 chr16 46382711 N chr16 46382782 N DUP 2
A00404:155:HV27LDSXX:3:1615:3775:30608 chr16 46382709 N chr16 46382855 N DUP 4
A00404:155:HV27LDSXX:4:1432:23213:27226 chr16 46382711 N chr16 46382782 N DUP 2
A00404:156:HV37TDSXX:1:1447:16893:29528 chr16 46382711 N chr16 46382782 N DUP 2
A00404:156:HV37TDSXX:2:1137:31891:20995 chr16 46382709 N chr16 46382855 N DUP 4
A00404:156:HV37TDSXX:2:1624:30499:20932 chr16 46382709 N chr16 46382855 N DUP 4
A00404:156:HV37TDSXX:2:2110:9995:28134 chr16 46382709 N chr16 46382855 N DUP 4
A00404:156:HV37TDSXX:2:2202:30337:19335 chr16 46382711 N chr16 46382782 N DUP 2
A00404:156:HV37TDSXX:2:2218:30346:29528 chr16 46382711 N chr16 46382782 N DUP 2
A00404:156:HV37TDSXX:4:2572:2917:33692 chr16 46382709 N chr16 46382855 N DUP 4
A00404:156:HV37TDSXX:2:2312:16251:27884 chr12 25174502 N chr12 25174639 N DEL 21
A00404:155:HV27LDSXX:3:2261:7554:9408 chr12 25174539 N chr12 25174600 N DUP 13
A00404:155:HV27LDSXX:2:1559:21965:20055 chr12 25174539 N chr12 25174600 N DUP 15
A00404:155:HV27LDSXX:2:1539:2609:22670 chr12 25174546 N chr12 25174607 N DUP 17
A00404:155:HV27LDSXX:1:1458:10990:21903 chr12 25174547 N chr12 25174608 N DUP 18
A00297:158:HT275DSXX:3:2365:9489:14074 chr12 25174548 N chr12 25174609 N DUP 19
A00297:158:HT275DSXX:4:1456:4924:18255 chr12 25174550 N chr12 25174611 N DUP 21
A00297:158:HT275DSXX:4:2433:28438:17644 chr12 25174577 N chr12 25174662 N DUP 22
A00404:155:HV27LDSXX:2:1370:11659:8594 chr12 25174558 N chr12 25174681 N DUP 19
A00404:155:HV27LDSXX:2:1370:12057:7686 chr12 25174558 N chr12 25174681 N DUP 19
A00404:155:HV27LDSXX:2:1552:25870:25285 chr12 25174577 N chr12 25174662 N DUP 21
A00404:155:HV27LDSXX:3:2103:11731:30420 chr12 25174577 N chr12 25174631 N DUP 24
A00404:156:HV37TDSXX:1:1527:21404:2832 chr12 25174557 N chr12 25174618 N DUP 6
A00297:158:HT275DSXX:1:2428:13376:18740 chr12 25174577 N chr12 25174662 N DUP 24
A00297:158:HT275DSXX:3:1115:4128:24298 chr12 25174557 N chr12 25174713 N DUP 21
A00297:158:HT275DSXX:3:1115:5168:23187 chr12 25174557 N chr12 25174713 N DUP 21
A00297:158:HT275DSXX:4:2315:22950:31344 chr12 25174557 N chr12 25174713 N DUP 20
A00297:158:HT275DSXX:4:1116:27353:25285 chr12 25174577 N chr12 25174631 N DUP 19
A00404:155:HV27LDSXX:1:1521:19027:31532 chr12 25174577 N chr12 25174631 N DUP 19
A00404:156:HV37TDSXX:2:1620:4372:2769 chr12 25174565 N chr12 25174697 N DUP 8
A00404:155:HV27LDSXX:2:1645:20717:2080 chr12 25174584 N chr12 25174837 N DUP 8
A00297:158:HT275DSXX:4:1204:12011:13056 chr12 25174565 N chr12 25174697 N DUP 13
A00404:156:HV37TDSXX:1:1166:22562:31829 chr12 25174510 N chr12 25174607 N DEL 22
A00404:156:HV37TDSXX:3:1668:23556:5963 chr12 25174577 N chr12 25174693 N DUP 23
A00297:158:HT275DSXX:2:2454:28782:12007 chr12 25174580 N chr12 25174705 N DUP 3
A00404:156:HV37TDSXX:1:1519:32235:5901 chr12 25174577 N chr12 25174662 N DUP 24
A00297:158:HT275DSXX:3:1115:4128:24298 chr12 25174584 N chr12 25174647 N DEL 10
A00297:158:HT275DSXX:3:1115:5168:23187 chr12 25174584 N chr12 25174647 N DEL 10
A00404:155:HV27LDSXX:2:1552:25870:25285 chr12 25174584 N chr12 25174647 N DEL 10
A00404:155:HV27LDSXX:3:2230:22914:33818 chr12 25174553 N chr12 25174647 N DEL 10
A00297:158:HT275DSXX:2:1477:10276:24298 chr12 25174540 N chr12 25174661 N DEL 1
A00404:155:HV27LDSXX:3:1439:6596:16203 chr12 25174703 N chr12 25174775 N DUP 14
A00297:158:HT275DSXX:4:2235:2645:8516 chr12 25174577 N chr12 25174742 N DUP 12
A00297:158:HT275DSXX:4:1257:30671:26522 chr12 25174577 N chr12 25174742 N DUP 12
A00404:155:HV27LDSXX:3:2619:22010:20134 chr12 25174604 N chr12 25174658 N DEL 22
A00404:156:HV37TDSXX:2:2640:15537:28275 chr12 25174604 N chr12 25174658 N DEL 22
A00404:156:HV37TDSXX:3:1366:31684:20635 chr12 25174604 N chr12 25174658 N DEL 24
A00297:158:HT275DSXX:4:2630:29984:1595 chr12 25174771 N chr12 25174823 N DUP 10
A00404:156:HV37TDSXX:1:2106:20076:19914 chr12 25174771 N chr12 25174823 N DUP 10
A00297:158:HT275DSXX:2:2324:16550:2848 chr12 25174581 N chr12 25174812 N DEL 5
A00297:158:HT275DSXX:2:2258:29116:23265 chr15 88554625 N chr15 88554686 N DEL 10
A00404:155:HV27LDSXX:1:1525:28510:23437 chr15 88554625 N chr15 88554686 N DEL 8
A00404:156:HV37TDSXX:3:1436:21504:31970 chr15 88554625 N chr15 88554686 N DEL 8
A00297:158:HT275DSXX:2:1674:27344:23390 chr15 88554628 N chr15 88554689 N DEL 5
A00404:156:HV37TDSXX:4:1425:20202:35697 chr15 88554628 N chr15 88554689 N DEL 5
A00404:156:HV37TDSXX:4:1415:17192:20525 chr15 88554622 N chr15 88554695 N DEL 5
A00404:156:HV37TDSXX:4:2572:11876:9032 chr6 19470482 N chr6 19470624 N DUP 8
A00404:156:HV37TDSXX:2:2562:7292:13307 chr18 559045 N chr18 559116 N DEL 9
A00297:158:HT275DSXX:3:1409:19651:27352 chr4 19771026 N chr4 19771093 N DEL 16
A00297:158:HT275DSXX:1:1304:30427:28291 chr2 217342313 N chr2 217342388 N DEL 9
A00404:155:HV27LDSXX:1:1463:22146:6433 chr2 217342314 N chr2 217342385 N DEL 10
A00404:155:HV27LDSXX:4:2555:9127:27320 chr7 136135289 N chr7 136135347 N DUP 6
A00404:156:HV37TDSXX:4:2405:16938:9533 chrX 46275320 N chrX 46275477 N DEL 5
A00297:158:HT275DSXX:2:1378:16459:16470 chrX 46275321 N chrX 46275478 N DEL 4
A00297:158:HT275DSXX:3:1244:30038:6950 chrX 46275324 N chrX 46275481 N DEL 1
A00404:155:HV27LDSXX:1:1418:6768:2566 chrX 46275321 N chrX 46275478 N DEL 4
A00404:155:HV27LDSXX:3:1543:11415:35540 chr3 141805130 N chr3 141805251 N DUP 5
A00404:155:HV27LDSXX:1:1353:15456:21652 chr10 123950282 N chr10 123950443 N DEL 32
A00404:156:HV37TDSXX:4:1232:24921:29465 chr2 239708552 N chr2 239708647 N DEL 6
A00404:156:HV37TDSXX:1:2341:4670:17597 chr2 239708567 N chr2 239708661 N DUP 7
A00404:156:HV37TDSXX:1:2341:4679:17581 chr2 239708567 N chr2 239708661 N DUP 7
A00404:155:HV27LDSXX:4:1454:27037:8015 chr1 143227141 N chr1 143227290 N DUP 5
A00404:155:HV27LDSXX:3:2221:29559:20901 chr1 143227163 N chr1 143227332 N DUP 6
A00297:158:HT275DSXX:3:1148:26006:19570 chr1 143227163 N chr1 143227332 N DUP 5
A00297:158:HT275DSXX:3:2115:1425:23563 chr1 143227163 N chr1 143227332 N DUP 5
A00404:155:HV27LDSXX:2:1533:10420:26177 chr1 143227184 N chr1 143227447 N DUP 5
A00404:155:HV27LDSXX:4:1628:23737:1642 chr1 143227184 N chr1 143227258 N DUP 5
A00404:156:HV37TDSXX:4:1668:5466:32847 chr1 143227184 N chr1 143227258 N DUP 5
A00297:158:HT275DSXX:4:2623:27624:17425 chr1 143227184 N chr1 143227258 N DUP 5
A00297:158:HT275DSXX:4:2623:27859:15483 chr1 143227184 N chr1 143227258 N DUP 5
A00297:158:HT275DSXX:4:2672:31910:34303 chr5 180594999 N chr5 180595088 N DUP 5
A00404:156:HV37TDSXX:4:2334:27868:33818 chr5 180595048 N chr5 180595105 N DUP 5
A00404:156:HV37TDSXX:1:2275:2871:18490 chr19 40470623 N chr19 40470950 N DEL 10
A00404:155:HV27LDSXX:3:1473:6207:18067 chr16 77714600 N chr16 77715030 N DUP 5
A00297:158:HT275DSXX:1:2450:27615:26271 chr16 85716579 N chr16 85716677 N DEL 3
